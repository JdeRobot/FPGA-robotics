// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 13 2019 00:12:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2Drone" view "INTERFACE"

module Pc2Drone (
    debug_state_output,
    uart_input,
    uart_data_rdy,
    debug_sinkdatavalid_output,
    uart_input_debug,
    frame_decoder_dv,
    clk_system);

    output [4:0] debug_state_output;
    input uart_input;
    output uart_data_rdy;
    output debug_sinkdatavalid_output;
    output uart_input_debug;
    output frame_decoder_dv;
    input clk_system;

    wire N__5663;
    wire N__5662;
    wire N__5661;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5616;
    wire N__5615;
    wire N__5614;
    wire N__5607;
    wire N__5606;
    wire N__5605;
    wire N__5598;
    wire N__5597;
    wire N__5596;
    wire N__5589;
    wire N__5588;
    wire N__5587;
    wire N__5580;
    wire N__5579;
    wire N__5578;
    wire N__5571;
    wire N__5570;
    wire N__5569;
    wire N__5552;
    wire N__5551;
    wire N__5550;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5511;
    wire N__5504;
    wire N__5503;
    wire N__5502;
    wire N__5501;
    wire N__5498;
    wire N__5497;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5492;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5464;
    wire N__5461;
    wire N__5460;
    wire N__5459;
    wire N__5458;
    wire N__5457;
    wire N__5456;
    wire N__5455;
    wire N__5450;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5432;
    wire N__5427;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5411;
    wire N__5406;
    wire N__5401;
    wire N__5398;
    wire N__5393;
    wire N__5378;
    wire N__5377;
    wire N__5376;
    wire N__5373;
    wire N__5372;
    wire N__5369;
    wire N__5368;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5361;
    wire N__5360;
    wire N__5359;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5338;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5318;
    wire N__5309;
    wire N__5300;
    wire N__5297;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5279;
    wire N__5278;
    wire N__5275;
    wire N__5274;
    wire N__5271;
    wire N__5266;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5245;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5233;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5212;
    wire N__5211;
    wire N__5208;
    wire N__5207;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5192;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5172;
    wire N__5167;
    wire N__5162;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5153;
    wire N__5148;
    wire N__5143;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5110;
    wire N__5105;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5099;
    wire N__5094;
    wire N__5089;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5074;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5057;
    wire N__5056;
    wire N__5055;
    wire N__5052;
    wire N__5051;
    wire N__5046;
    wire N__5041;
    wire N__5036;
    wire N__5033;
    wire N__5032;
    wire N__5031;
    wire N__5030;
    wire N__5027;
    wire N__5026;
    wire N__5021;
    wire N__5018;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5010;
    wire N__5009;
    wire N__5008;
    wire N__5003;
    wire N__5000;
    wire N__4995;
    wire N__4990;
    wire N__4987;
    wire N__4982;
    wire N__4979;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4942;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4893;
    wire N__4888;
    wire N__4883;
    wire N__4882;
    wire N__4881;
    wire N__4880;
    wire N__4879;
    wire N__4878;
    wire N__4877;
    wire N__4876;
    wire N__4875;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4871;
    wire N__4870;
    wire N__4869;
    wire N__4868;
    wire N__4867;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4860;
    wire N__4859;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4784;
    wire N__4781;
    wire N__4780;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4757;
    wire N__4754;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4731;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4719;
    wire N__4716;
    wire N__4709;
    wire N__4706;
    wire N__4705;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4688;
    wire N__4685;
    wire N__4684;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4667;
    wire N__4664;
    wire N__4663;
    wire N__4662;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4648;
    wire N__4643;
    wire N__4640;
    wire N__4639;
    wire N__4634;
    wire N__4633;
    wire N__4632;
    wire N__4631;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4617;
    wire N__4614;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4499;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4438;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4426;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4357;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4324;
    wire N__4321;
    wire N__4320;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4295;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4270;
    wire N__4269;
    wire N__4264;
    wire N__4261;
    wire N__4256;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4244;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4183;
    wire N__4182;
    wire N__4179;
    wire N__4174;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4156;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4093;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4081;
    wire N__4080;
    wire N__4077;
    wire N__4076;
    wire N__4071;
    wire N__4066;
    wire N__4061;
    wire N__4060;
    wire N__4059;
    wire N__4056;
    wire N__4051;
    wire N__4046;
    wire N__4045;
    wire N__4040;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4031;
    wire N__4024;
    wire N__4019;
    wire N__4018;
    wire N__4015;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4003;
    wire N__4002;
    wire N__4001;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3987;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3967;
    wire N__3966;
    wire N__3965;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3941;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3925;
    wire N__3924;
    wire N__3921;
    wire N__3920;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3886;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3851;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3843;
    wire N__3842;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3828;
    wire N__3821;
    wire N__3818;
    wire N__3817;
    wire N__3814;
    wire N__3813;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3801;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3780;
    wire N__3779;
    wire N__3774;
    wire N__3773;
    wire N__3772;
    wire N__3771;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3754;
    wire N__3749;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3730;
    wire N__3725;
    wire N__3722;
    wire N__3721;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3709;
    wire N__3704;
    wire N__3701;
    wire N__3700;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3682;
    wire N__3681;
    wire N__3678;
    wire N__3677;
    wire N__3676;
    wire N__3673;
    wire N__3672;
    wire N__3671;
    wire N__3670;
    wire N__3669;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3652;
    wire N__3651;
    wire N__3650;
    wire N__3647;
    wire N__3638;
    wire N__3635;
    wire N__3626;
    wire N__3619;
    wire N__3616;
    wire N__3613;
    wire N__3608;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3571;
    wire N__3568;
    wire N__3567;
    wire N__3566;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3539;
    wire N__3536;
    wire N__3535;
    wire N__3534;
    wire N__3531;
    wire N__3526;
    wire N__3521;
    wire N__3520;
    wire N__3517;
    wire N__3514;
    wire N__3513;
    wire N__3512;
    wire N__3511;
    wire N__3506;
    wire N__3505;
    wire N__3502;
    wire N__3501;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3483;
    wire N__3480;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3454;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3417;
    wire N__3412;
    wire N__3407;
    wire N__3404;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3396;
    wire N__3393;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3371;
    wire N__3370;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3362;
    wire N__3361;
    wire N__3360;
    wire N__3357;
    wire N__3356;
    wire N__3353;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3338;
    wire N__3335;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3317;
    wire N__3314;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3287;
    wire N__3284;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3260;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3242;
    wire N__3239;
    wire N__3238;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3221;
    wire N__3218;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3206;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3173;
    wire N__3172;
    wire N__3171;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3133;
    wire N__3132;
    wire N__3131;
    wire N__3130;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3098;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3080;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3065;
    wire N__3062;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3050;
    wire N__3047;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3035;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3023;
    wire N__3020;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3005;
    wire N__3002;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2990;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2978;
    wire N__2975;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2960;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2948;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2936;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2921;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2876;
    wire N__2875;
    wire N__2872;
    wire N__2869;
    wire N__2868;
    wire N__2867;
    wire N__2866;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2842;
    wire N__2841;
    wire N__2840;
    wire N__2831;
    wire N__2828;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2807;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2795;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2783;
    wire N__2782;
    wire N__2781;
    wire N__2778;
    wire N__2777;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2771;
    wire N__2764;
    wire N__2757;
    wire N__2750;
    wire N__2747;
    wire N__2744;
    wire N__2741;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2722;
    wire N__2721;
    wire N__2714;
    wire N__2711;
    wire N__2710;
    wire N__2709;
    wire N__2708;
    wire N__2707;
    wire N__2706;
    wire N__2705;
    wire N__2704;
    wire N__2701;
    wire N__2698;
    wire N__2697;
    wire N__2696;
    wire N__2693;
    wire N__2682;
    wire N__2677;
    wire N__2672;
    wire N__2663;
    wire N__2662;
    wire N__2661;
    wire N__2658;
    wire N__2657;
    wire N__2656;
    wire N__2653;
    wire N__2652;
    wire N__2651;
    wire N__2650;
    wire N__2649;
    wire N__2648;
    wire N__2645;
    wire N__2644;
    wire N__2633;
    wire N__2628;
    wire N__2623;
    wire N__2618;
    wire N__2609;
    wire N__2608;
    wire N__2607;
    wire N__2606;
    wire N__2605;
    wire N__2604;
    wire N__2603;
    wire N__2602;
    wire N__2601;
    wire N__2600;
    wire N__2599;
    wire N__2598;
    wire N__2587;
    wire N__2582;
    wire N__2575;
    wire N__2570;
    wire N__2561;
    wire N__2558;
    wire N__2555;
    wire N__2552;
    wire N__2549;
    wire N__2546;
    wire N__2543;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2528;
    wire N__2525;
    wire N__2522;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2507;
    wire N__2504;
    wire N__2501;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2489;
    wire N__2486;
    wire N__2483;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2471;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2447;
    wire N__2444;
    wire N__2441;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2429;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2417;
    wire N__2416;
    wire N__2413;
    wire N__2410;
    wire N__2405;
    wire N__2402;
    wire N__2399;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2374;
    wire N__2371;
    wire N__2366;
    wire N__2365;
    wire N__2362;
    wire N__2359;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2347;
    wire N__2342;
    wire N__2339;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2324;
    wire N__2321;
    wire GNDG0;
    wire VCCG0;
    wire frame_decoder_dv_c;
    wire uart_input_c;
    wire \uart_sync.aux_0__0_Z0Z_0 ;
    wire \uart_sync.aux_1__0_Z0Z_0 ;
    wire \uart_sync.aux_2__0_Z0Z_0 ;
    wire \uart_sync.aux_3__0_Z0Z_0 ;
    wire \uart.N_133_0_cascade_ ;
    wire \uart.N_133_0 ;
    wire \uart.data_Auxce_0_6_cascade_ ;
    wire \uart.CO1_0 ;
    wire bfn_8_1_0_;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire bfn_8_2_0_;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire bfn_8_3_0_;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \uart.data_Auxce_0_5 ;
    wire \uart.timer_Count_RNI9M0NZ0Z_1 ;
    wire \uart.timer_Count_RNILKMA1Z0Z_0_cascade_ ;
    wire \uart.un1_state_2_0_cascade_ ;
    wire \uart.un1_state_2_0 ;
    wire \uart.data_Auxce_0_0_4 ;
    wire \uart.data_Auxce_0_0_0 ;
    wire \uart.data_Auxce_0_1 ;
    wire \uart.data_Auxce_0_0_2 ;
    wire \uart.un1_state_5_0 ;
    wire \uart.bit_CountZ0Z_2 ;
    wire \uart.bit_CountZ0Z_1 ;
    wire \uart.bit_CountZ0Z_0 ;
    wire \uart.data_Auxce_0_3 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.reset6_14_cascade_ ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.count_1_1 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire \reset_module_System.reset6_3_cascade_ ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_11 ;
    wire \reset_module_System.reset6_19 ;
    wire \uart.N_169_cascade_ ;
    wire \uart.state_srsts_i_1_3_cascade_ ;
    wire \uart.data_AuxZ0Z_0 ;
    wire \uart.data_AuxZ0Z_2 ;
    wire \uart.data_AuxZ0Z_3 ;
    wire \uart.data_AuxZ0Z_5 ;
    wire \uart.data_AuxZ0Z_7 ;
    wire \uart.timer_Count10lto5_0_0_cascade_ ;
    wire \uart.N_177 ;
    wire \uart.N_168_cascade_ ;
    wire \uart.state_RNIAFHLZ0Z_4 ;
    wire \uart.stateZ0Z_1 ;
    wire \uart.N_151_cascade_ ;
    wire \uart.stateZ0Z_2 ;
    wire \uart.stateZ0Z_3 ;
    wire \uart.state_srsts_i_1_1_3 ;
    wire \uart.N_166_cascade_ ;
    wire \uart.state_srsts_0_1_0_cascade_ ;
    wire \uart.stateZ0Z_0 ;
    wire \uart_frame_decoder.N_43 ;
    wire \uart_frame_decoder.N_43_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_ ;
    wire \uart_frame_decoder.N_81_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ;
    wire uart_data_3;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_ ;
    wire uart_data_2;
    wire uart_data_5;
    wire uart_data_7;
    wire uart_data_0;
    wire \uart_frame_decoder.N_79_4 ;
    wire \uart_frame_decoder.N_79_4_cascade_ ;
    wire uart_input_sync;
    wire \uart.data_8_0_cascade_ ;
    wire \uart.state_srsts_0_a3_1_4 ;
    wire \uart.N_152_0_cascade_ ;
    wire \uart.N_167 ;
    wire \uart.N_159 ;
    wire \uart.N_167_cascade_ ;
    wire \uart.N_180 ;
    wire \uart.N_152_0 ;
    wire \uart.stateZ0Z_4 ;
    wire \uart.N_145_0 ;
    wire \uart.state_1_sqmuxa ;
    wire \uart.state_1_sqmuxa_cascade_ ;
    wire bfn_10_5_0_;
    wire \uart.timer_CountZ0Z_2 ;
    wire \uart.un4_timer_Count_1_cry_1 ;
    wire \uart.timer_CountZ0Z_3 ;
    wire \uart.un4_timer_Count_1_cry_2 ;
    wire \uart.timer_CountZ0Z_4 ;
    wire \uart.un4_timer_Count_1_cry_3 ;
    wire \uart.timer_CountZ0Z_5 ;
    wire \uart.un4_timer_Count_1_cry_4 ;
    wire \uart.timer_CountZ0Z_6 ;
    wire \uart.un4_timer_Count_1_cry_5 ;
    wire \uart.un4_timer_Count_1_cry_6 ;
    wire \uart.timer_CountZ0Z_7 ;
    wire bfn_11_1_0_;
    wire \uart_frame_decoder.count8_axb_1 ;
    wire \uart_frame_decoder.count8_cry_0 ;
    wire \uart_frame_decoder.count_i_2 ;
    wire \uart_frame_decoder.count8_cry_1 ;
    wire \uart_frame_decoder.count8 ;
    wire \uart_frame_decoder.count8_THRU_CO ;
    wire \uart_frame_decoder.count8_THRU_CO_cascade_ ;
    wire \uart_frame_decoder.N_37 ;
    wire \uart_frame_decoder.N_37_cascade_ ;
    wire \uart_frame_decoder.countZ0Z_1 ;
    wire \uart_frame_decoder.countZ0Z_2 ;
    wire CONSTANT_ONE_NET;
    wire \uart_frame_decoder.count8_0 ;
    wire \uart_frame_decoder.count8_0_i ;
    wire \uart_frame_decoder.N_4_0_cascade_ ;
    wire \uart_frame_decoder.g0_1_0_1 ;
    wire \uart_frame_decoder.g0_1_a3_3 ;
    wire \uart_frame_decoder.WDT8lto15_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10 ;
    wire \uart_frame_decoder.state_1_ns_i_i_a2_1_1_0 ;
    wire \uart_frame_decoder.state_1Z0Z_0 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_ ;
    wire \uart_frame_decoder.N_35_i_1 ;
    wire \uart.timer_CountZ0Z_1 ;
    wire \uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ;
    wire \uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_ ;
    wire \uart_frame_decoder.WDT8lt13_cascade_ ;
    wire \uart_frame_decoder.state_1_ns_i_i_a2_0_0 ;
    wire \uart_frame_decoder.WDT8lt13 ;
    wire \uart_frame_decoder.WDT8lto15 ;
    wire \uart_frame_decoder.N_80 ;
    wire \uart.timer_CountZ0Z_0 ;
    wire \uart.timer_Count_1_sqmuxa_i ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ;
    wire \uart_frame_decoder.N_99 ;
    wire \uart_frame_decoder.N_92 ;
    wire \uart.data_AuxZ0Z_1 ;
    wire uart_data_1;
    wire \uart.data_AuxZ0Z_4 ;
    wire uart_data_4;
    wire \uart.data_AuxZ0Z_6 ;
    wire uart_data_6;
    wire \uart.state_1_sqmuxa_0 ;
    wire \uart.timer_Count_RNIS4183Z0Z_7 ;
    wire \uart_frame_decoder.WDT8_0_i ;
    wire \uart_frame_decoder.WDTZ0Z_0 ;
    wire bfn_12_2_0_;
    wire \uart_frame_decoder.WDTZ0Z_1 ;
    wire \uart_frame_decoder.un1_WDT_cry_0 ;
    wire \uart_frame_decoder.WDTZ0Z_2 ;
    wire \uart_frame_decoder.un1_WDT_cry_1 ;
    wire \uart_frame_decoder.WDTZ0Z_3 ;
    wire \uart_frame_decoder.un1_WDT_cry_2 ;
    wire \uart_frame_decoder.WDTZ0Z_4 ;
    wire \uart_frame_decoder.un1_WDT_cry_3 ;
    wire \uart_frame_decoder.WDTZ0Z_5 ;
    wire \uart_frame_decoder.un1_WDT_cry_4 ;
    wire \uart_frame_decoder.WDTZ0Z_6 ;
    wire \uart_frame_decoder.un1_WDT_cry_5 ;
    wire \uart_frame_decoder.WDTZ0Z_7 ;
    wire \uart_frame_decoder.un1_WDT_cry_6 ;
    wire \uart_frame_decoder.un1_WDT_cry_7 ;
    wire \uart_frame_decoder.WDTZ0Z_8 ;
    wire bfn_12_3_0_;
    wire \uart_frame_decoder.WDTZ0Z_9 ;
    wire \uart_frame_decoder.un1_WDT_cry_8 ;
    wire \uart_frame_decoder.WDTZ0Z_10 ;
    wire \uart_frame_decoder.un1_WDT_cry_9 ;
    wire \uart_frame_decoder.WDTZ0Z_11 ;
    wire \uart_frame_decoder.un1_WDT_cry_10 ;
    wire \uart_frame_decoder.WDTZ0Z_12 ;
    wire \uart_frame_decoder.un1_WDT_cry_11 ;
    wire \uart_frame_decoder.WDTZ0Z_13 ;
    wire \uart_frame_decoder.un1_WDT_cry_12 ;
    wire \uart_frame_decoder.WDTZ0Z_14 ;
    wire \uart_frame_decoder.un1_WDT_cry_13 ;
    wire \uart_frame_decoder.un1_WDT_cry_14 ;
    wire \uart_frame_decoder.WDTZ0Z_15 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10 ;
    wire \uart_frame_decoder.state_1_ns_0_i_a2_0_d_10 ;
    wire \uart_frame_decoder.N_85 ;
    wire clk_system_c_g;
    wire reset_module_System_reset_iso;
    wire uart_data_rdy_c;
    wire reset_system;
    wire \uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ;
    wire \uart_frame_decoder.state_1Z0Z_4 ;
    wire uart_frame_decoder_N_307_i;
    wire \uart_frame_decoder.state_1Z0Z_8 ;
    wire uart_frame_decoder_N_308_i;
    wire \uart_frame_decoder.state_1Z0Z_1 ;
    wire \uart_frame_decoder.state_1Z0Z_9 ;
    wire \uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_ ;
    wire \uart_frame_decoder.state_1Z0Z_5 ;
    wire uart_frame_decoder_N_305_i;
    wire \uart_frame_decoder.state_1Z0Z_6 ;
    wire \uart_frame_decoder.state_1Z0Z_7 ;
    wire \uart_frame_decoder.N_306_1 ;
    wire \uart_frame_decoder.state_1Z0Z_2 ;
    wire \uart_frame_decoder.state_1Z0Z_3 ;
    wire \uart_frame_decoder.N_306_1_cascade_ ;
    wire \uart_frame_decoder.state_1Z0Z_10 ;
    wire uart_frame_decoder_N_306_i;
    wire _gnd_net_;

    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5661),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__5663),
            .DIN(N__5662),
            .DOUT(N__5661),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__5663),
            .PADOUT(N__5662),
            .PADIN(N__5661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD debug_state_output_obuf_4_iopad (
            .OE(N__5652),
            .DIN(N__5651),
            .DOUT(N__5650),
            .PACKAGEPIN(debug_state_output[4]));
    defparam debug_state_output_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_4_preio (
            .PADOEN(N__5652),
            .PADOUT(N__5651),
            .PADIN(N__5650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_1_iopad (
            .OE(N__5643),
            .DIN(N__5642),
            .DOUT(N__5641),
            .PACKAGEPIN(debug_state_output[1]));
    defparam debug_state_output_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_1_preio (
            .PADOEN(N__5643),
            .PADOUT(N__5642),
            .PADIN(N__5641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4970),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_data_rdy_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_data_rdy_obuf_iopad (
            .OE(N__5634),
            .DIN(N__5633),
            .DOUT(N__5632),
            .PACKAGEPIN(uart_data_rdy));
    defparam uart_data_rdy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_data_rdy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_data_rdy_obuf_preio (
            .PADOEN(N__5634),
            .PADOUT(N__5633),
            .PADIN(N__5632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5503),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_3_iopad (
            .OE(N__5625),
            .DIN(N__5624),
            .DOUT(N__5623),
            .PACKAGEPIN(debug_state_output[3]));
    defparam debug_state_output_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_3_preio (
            .PADOEN(N__5625),
            .PADOUT(N__5624),
            .PADIN(N__5623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_sinkdatavalid_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_sinkdatavalid_output_obuf_iopad (
            .OE(N__5616),
            .DIN(N__5615),
            .DOUT(N__5614),
            .PACKAGEPIN(debug_sinkdatavalid_output));
    defparam debug_sinkdatavalid_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_sinkdatavalid_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_sinkdatavalid_output_obuf_preio (
            .PADOEN(N__5616),
            .PADOUT(N__5615),
            .PADIN(N__5614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam frame_decoder_dv_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD frame_decoder_dv_obuf_iopad (
            .OE(N__5607),
            .DIN(N__5606),
            .DOUT(N__5605),
            .PACKAGEPIN(frame_decoder_dv));
    defparam frame_decoder_dv_obuf_preio.NEG_TRIGGER=1'b0;
    defparam frame_decoder_dv_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO frame_decoder_dv_obuf_preio (
            .PADOEN(N__5607),
            .PADOUT(N__5606),
            .PADIN(N__5605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2393),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_ibuf_iopad (
            .OE(N__5598),
            .DIN(N__5597),
            .DOUT(N__5596),
            .PACKAGEPIN(uart_input));
    defparam uart_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_ibuf_preio (
            .PADOEN(N__5598),
            .PADOUT(N__5597),
            .PADIN(N__5596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_0_iopad (
            .OE(N__5589),
            .DIN(N__5588),
            .DOUT(N__5587),
            .PACKAGEPIN(debug_state_output[0]));
    defparam debug_state_output_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_0_preio (
            .PADOEN(N__5589),
            .PADOUT(N__5588),
            .PADIN(N__5587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5138),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_state_output_obuf_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_state_output_obuf_2_iopad (
            .OE(N__5580),
            .DIN(N__5579),
            .DOUT(N__5578),
            .PACKAGEPIN(debug_state_output[2]));
    defparam debug_state_output_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam debug_state_output_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_state_output_obuf_2_preio (
            .PADOEN(N__5580),
            .PADOUT(N__5579),
            .PADIN(N__5578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5261),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_debug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_debug_obuf_iopad (
            .OE(N__5571),
            .DIN(N__5570),
            .DOUT(N__5569),
            .PACKAGEPIN(uart_input_debug));
    defparam uart_input_debug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_debug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO uart_input_debug_obuf_preio (
            .PADOEN(N__5571),
            .PADOUT(N__5570),
            .PADIN(N__5569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    SRMux I__1274 (
            .O(N__5552),
            .I(N__5546));
    SRMux I__1273 (
            .O(N__5551),
            .I(N__5543));
    SRMux I__1272 (
            .O(N__5550),
            .I(N__5540));
    SRMux I__1271 (
            .O(N__5549),
            .I(N__5537));
    LocalMux I__1270 (
            .O(N__5546),
            .I(N__5533));
    LocalMux I__1269 (
            .O(N__5543),
            .I(N__5530));
    LocalMux I__1268 (
            .O(N__5540),
            .I(N__5527));
    LocalMux I__1267 (
            .O(N__5537),
            .I(N__5524));
    SRMux I__1266 (
            .O(N__5536),
            .I(N__5521));
    Span4Mux_v I__1265 (
            .O(N__5533),
            .I(N__5518));
    Span4Mux_s0_v I__1264 (
            .O(N__5530),
            .I(N__5511));
    Span4Mux_v I__1263 (
            .O(N__5527),
            .I(N__5511));
    Span4Mux_v I__1262 (
            .O(N__5524),
            .I(N__5511));
    LocalMux I__1261 (
            .O(N__5521),
            .I(reset_module_System_reset_iso));
    Odrv4 I__1260 (
            .O(N__5518),
            .I(reset_module_System_reset_iso));
    Odrv4 I__1259 (
            .O(N__5511),
            .I(reset_module_System_reset_iso));
    CascadeMux I__1258 (
            .O(N__5504),
            .I(N__5498));
    IoInMux I__1257 (
            .O(N__5503),
            .I(N__5488));
    IoInMux I__1256 (
            .O(N__5502),
            .I(N__5485));
    InMux I__1255 (
            .O(N__5501),
            .I(N__5482));
    InMux I__1254 (
            .O(N__5498),
            .I(N__5479));
    InMux I__1253 (
            .O(N__5497),
            .I(N__5464));
    InMux I__1252 (
            .O(N__5496),
            .I(N__5464));
    InMux I__1251 (
            .O(N__5495),
            .I(N__5464));
    InMux I__1250 (
            .O(N__5494),
            .I(N__5464));
    InMux I__1249 (
            .O(N__5493),
            .I(N__5464));
    InMux I__1248 (
            .O(N__5492),
            .I(N__5464));
    InMux I__1247 (
            .O(N__5491),
            .I(N__5464));
    LocalMux I__1246 (
            .O(N__5488),
            .I(N__5461));
    LocalMux I__1245 (
            .O(N__5485),
            .I(N__5450));
    LocalMux I__1244 (
            .O(N__5482),
            .I(N__5450));
    LocalMux I__1243 (
            .O(N__5479),
            .I(N__5445));
    LocalMux I__1242 (
            .O(N__5464),
            .I(N__5445));
    Span4Mux_s2_v I__1241 (
            .O(N__5461),
            .I(N__5440));
    InMux I__1240 (
            .O(N__5460),
            .I(N__5437));
    InMux I__1239 (
            .O(N__5459),
            .I(N__5432));
    InMux I__1238 (
            .O(N__5458),
            .I(N__5432));
    InMux I__1237 (
            .O(N__5457),
            .I(N__5427));
    InMux I__1236 (
            .O(N__5456),
            .I(N__5427));
    InMux I__1235 (
            .O(N__5455),
            .I(N__5424));
    Span4Mux_s2_v I__1234 (
            .O(N__5450),
            .I(N__5419));
    Span4Mux_h I__1233 (
            .O(N__5445),
            .I(N__5416));
    InMux I__1232 (
            .O(N__5444),
            .I(N__5411));
    InMux I__1231 (
            .O(N__5443),
            .I(N__5411));
    Span4Mux_h I__1230 (
            .O(N__5440),
            .I(N__5406));
    LocalMux I__1229 (
            .O(N__5437),
            .I(N__5406));
    LocalMux I__1228 (
            .O(N__5432),
            .I(N__5401));
    LocalMux I__1227 (
            .O(N__5427),
            .I(N__5401));
    LocalMux I__1226 (
            .O(N__5424),
            .I(N__5398));
    InMux I__1225 (
            .O(N__5423),
            .I(N__5393));
    InMux I__1224 (
            .O(N__5422),
            .I(N__5393));
    Odrv4 I__1223 (
            .O(N__5419),
            .I(uart_data_rdy_c));
    Odrv4 I__1222 (
            .O(N__5416),
            .I(uart_data_rdy_c));
    LocalMux I__1221 (
            .O(N__5411),
            .I(uart_data_rdy_c));
    Odrv4 I__1220 (
            .O(N__5406),
            .I(uart_data_rdy_c));
    Odrv4 I__1219 (
            .O(N__5401),
            .I(uart_data_rdy_c));
    Odrv4 I__1218 (
            .O(N__5398),
            .I(uart_data_rdy_c));
    LocalMux I__1217 (
            .O(N__5393),
            .I(uart_data_rdy_c));
    InMux I__1216 (
            .O(N__5378),
            .I(N__5373));
    InMux I__1215 (
            .O(N__5377),
            .I(N__5369));
    InMux I__1214 (
            .O(N__5376),
            .I(N__5365));
    LocalMux I__1213 (
            .O(N__5373),
            .I(N__5355));
    InMux I__1212 (
            .O(N__5372),
            .I(N__5352));
    LocalMux I__1211 (
            .O(N__5369),
            .I(N__5349));
    InMux I__1210 (
            .O(N__5368),
            .I(N__5346));
    LocalMux I__1209 (
            .O(N__5365),
            .I(N__5343));
    InMux I__1208 (
            .O(N__5364),
            .I(N__5338));
    InMux I__1207 (
            .O(N__5363),
            .I(N__5338));
    InMux I__1206 (
            .O(N__5362),
            .I(N__5331));
    InMux I__1205 (
            .O(N__5361),
            .I(N__5331));
    InMux I__1204 (
            .O(N__5360),
            .I(N__5331));
    InMux I__1203 (
            .O(N__5359),
            .I(N__5328));
    InMux I__1202 (
            .O(N__5358),
            .I(N__5325));
    Span4Mux_v I__1201 (
            .O(N__5355),
            .I(N__5318));
    LocalMux I__1200 (
            .O(N__5352),
            .I(N__5318));
    Span4Mux_v I__1199 (
            .O(N__5349),
            .I(N__5318));
    LocalMux I__1198 (
            .O(N__5346),
            .I(N__5309));
    Span4Mux_v I__1197 (
            .O(N__5343),
            .I(N__5309));
    LocalMux I__1196 (
            .O(N__5338),
            .I(N__5309));
    LocalMux I__1195 (
            .O(N__5331),
            .I(N__5309));
    LocalMux I__1194 (
            .O(N__5328),
            .I(reset_system));
    LocalMux I__1193 (
            .O(N__5325),
            .I(reset_system));
    Odrv4 I__1192 (
            .O(N__5318),
            .I(reset_system));
    Odrv4 I__1191 (
            .O(N__5309),
            .I(reset_system));
    SRMux I__1190 (
            .O(N__5300),
            .I(N__5297));
    LocalMux I__1189 (
            .O(N__5297),
            .I(N__5293));
    SRMux I__1188 (
            .O(N__5296),
            .I(N__5290));
    Span4Mux_s2_v I__1187 (
            .O(N__5293),
            .I(N__5287));
    LocalMux I__1186 (
            .O(N__5290),
            .I(N__5284));
    Odrv4 I__1185 (
            .O(N__5287),
            .I(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ));
    Odrv4 I__1184 (
            .O(N__5284),
            .I(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ));
    CascadeMux I__1183 (
            .O(N__5279),
            .I(N__5275));
    InMux I__1182 (
            .O(N__5278),
            .I(N__5271));
    InMux I__1181 (
            .O(N__5275),
            .I(N__5266));
    InMux I__1180 (
            .O(N__5274),
            .I(N__5266));
    LocalMux I__1179 (
            .O(N__5271),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    LocalMux I__1178 (
            .O(N__5266),
            .I(\uart_frame_decoder.state_1Z0Z_4 ));
    IoInMux I__1177 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__1176 (
            .O(N__5258),
            .I(N__5255));
    IoSpan4Mux I__1175 (
            .O(N__5255),
            .I(N__5252));
    IoSpan4Mux I__1174 (
            .O(N__5252),
            .I(N__5249));
    Odrv4 I__1173 (
            .O(N__5249),
            .I(uart_frame_decoder_N_307_i));
    CascadeMux I__1172 (
            .O(N__5246),
            .I(N__5241));
    InMux I__1171 (
            .O(N__5245),
            .I(N__5238));
    InMux I__1170 (
            .O(N__5244),
            .I(N__5233));
    InMux I__1169 (
            .O(N__5241),
            .I(N__5233));
    LocalMux I__1168 (
            .O(N__5238),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    LocalMux I__1167 (
            .O(N__5233),
            .I(\uart_frame_decoder.state_1Z0Z_8 ));
    IoInMux I__1166 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__1165 (
            .O(N__5225),
            .I(N__5222));
    Span4Mux_s3_v I__1164 (
            .O(N__5222),
            .I(N__5219));
    Odrv4 I__1163 (
            .O(N__5219),
            .I(uart_frame_decoder_N_308_i));
    InMux I__1162 (
            .O(N__5216),
            .I(N__5212));
    InMux I__1161 (
            .O(N__5215),
            .I(N__5208));
    LocalMux I__1160 (
            .O(N__5212),
            .I(N__5203));
    InMux I__1159 (
            .O(N__5211),
            .I(N__5200));
    LocalMux I__1158 (
            .O(N__5208),
            .I(N__5197));
    InMux I__1157 (
            .O(N__5207),
            .I(N__5192));
    InMux I__1156 (
            .O(N__5206),
            .I(N__5192));
    Odrv4 I__1155 (
            .O(N__5203),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__1154 (
            .O(N__5200),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    Odrv4 I__1153 (
            .O(N__5197),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    LocalMux I__1152 (
            .O(N__5192),
            .I(\uart_frame_decoder.state_1Z0Z_1 ));
    CascadeMux I__1151 (
            .O(N__5183),
            .I(N__5177));
    InMux I__1150 (
            .O(N__5182),
            .I(N__5172));
    InMux I__1149 (
            .O(N__5181),
            .I(N__5172));
    InMux I__1148 (
            .O(N__5180),
            .I(N__5167));
    InMux I__1147 (
            .O(N__5177),
            .I(N__5167));
    LocalMux I__1146 (
            .O(N__5172),
            .I(\uart_frame_decoder.state_1Z0Z_9 ));
    LocalMux I__1145 (
            .O(N__5167),
            .I(\uart_frame_decoder.state_1Z0Z_9 ));
    CascadeMux I__1144 (
            .O(N__5162),
            .I(\uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_ ));
    CascadeMux I__1143 (
            .O(N__5159),
            .I(N__5154));
    InMux I__1142 (
            .O(N__5158),
            .I(N__5148));
    InMux I__1141 (
            .O(N__5157),
            .I(N__5148));
    InMux I__1140 (
            .O(N__5154),
            .I(N__5143));
    InMux I__1139 (
            .O(N__5153),
            .I(N__5143));
    LocalMux I__1138 (
            .O(N__5148),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    LocalMux I__1137 (
            .O(N__5143),
            .I(\uart_frame_decoder.state_1Z0Z_5 ));
    IoInMux I__1136 (
            .O(N__5138),
            .I(N__5135));
    LocalMux I__1135 (
            .O(N__5135),
            .I(N__5132));
    IoSpan4Mux I__1134 (
            .O(N__5132),
            .I(N__5129));
    Span4Mux_s3_v I__1133 (
            .O(N__5129),
            .I(N__5126));
    Odrv4 I__1132 (
            .O(N__5126),
            .I(uart_frame_decoder_N_305_i));
    CascadeMux I__1131 (
            .O(N__5123),
            .I(N__5119));
    InMux I__1130 (
            .O(N__5122),
            .I(N__5115));
    InMux I__1129 (
            .O(N__5119),
            .I(N__5110));
    InMux I__1128 (
            .O(N__5118),
            .I(N__5110));
    LocalMux I__1127 (
            .O(N__5115),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    LocalMux I__1126 (
            .O(N__5110),
            .I(\uart_frame_decoder.state_1Z0Z_6 ));
    CascadeMux I__1125 (
            .O(N__5105),
            .I(N__5099));
    InMux I__1124 (
            .O(N__5104),
            .I(N__5094));
    InMux I__1123 (
            .O(N__5103),
            .I(N__5094));
    InMux I__1122 (
            .O(N__5102),
            .I(N__5089));
    InMux I__1121 (
            .O(N__5099),
            .I(N__5089));
    LocalMux I__1120 (
            .O(N__5094),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    LocalMux I__1119 (
            .O(N__5089),
            .I(\uart_frame_decoder.state_1Z0Z_7 ));
    InMux I__1118 (
            .O(N__5084),
            .I(N__5081));
    LocalMux I__1117 (
            .O(N__5081),
            .I(\uart_frame_decoder.N_306_1 ));
    InMux I__1116 (
            .O(N__5078),
            .I(N__5075));
    LocalMux I__1115 (
            .O(N__5075),
            .I(N__5070));
    InMux I__1114 (
            .O(N__5074),
            .I(N__5067));
    InMux I__1113 (
            .O(N__5073),
            .I(N__5064));
    Odrv4 I__1112 (
            .O(N__5070),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    LocalMux I__1111 (
            .O(N__5067),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    LocalMux I__1110 (
            .O(N__5064),
            .I(\uart_frame_decoder.state_1Z0Z_2 ));
    CascadeMux I__1109 (
            .O(N__5057),
            .I(N__5052));
    InMux I__1108 (
            .O(N__5056),
            .I(N__5046));
    InMux I__1107 (
            .O(N__5055),
            .I(N__5046));
    InMux I__1106 (
            .O(N__5052),
            .I(N__5041));
    InMux I__1105 (
            .O(N__5051),
            .I(N__5041));
    LocalMux I__1104 (
            .O(N__5046),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    LocalMux I__1103 (
            .O(N__5041),
            .I(\uart_frame_decoder.state_1Z0Z_3 ));
    CascadeMux I__1102 (
            .O(N__5036),
            .I(\uart_frame_decoder.N_306_1_cascade_ ));
    InMux I__1101 (
            .O(N__5033),
            .I(N__5027));
    InMux I__1100 (
            .O(N__5032),
            .I(N__5021));
    InMux I__1099 (
            .O(N__5031),
            .I(N__5021));
    InMux I__1098 (
            .O(N__5030),
            .I(N__5018));
    LocalMux I__1097 (
            .O(N__5027),
            .I(N__5014));
    InMux I__1096 (
            .O(N__5026),
            .I(N__5011));
    LocalMux I__1095 (
            .O(N__5021),
            .I(N__5003));
    LocalMux I__1094 (
            .O(N__5018),
            .I(N__5003));
    InMux I__1093 (
            .O(N__5017),
            .I(N__5000));
    Span4Mux_s1_v I__1092 (
            .O(N__5014),
            .I(N__4995));
    LocalMux I__1091 (
            .O(N__5011),
            .I(N__4995));
    InMux I__1090 (
            .O(N__5010),
            .I(N__4990));
    InMux I__1089 (
            .O(N__5009),
            .I(N__4990));
    InMux I__1088 (
            .O(N__5008),
            .I(N__4987));
    Span4Mux_h I__1087 (
            .O(N__5003),
            .I(N__4982));
    LocalMux I__1086 (
            .O(N__5000),
            .I(N__4982));
    Span4Mux_h I__1085 (
            .O(N__4995),
            .I(N__4979));
    LocalMux I__1084 (
            .O(N__4990),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    LocalMux I__1083 (
            .O(N__4987),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    Odrv4 I__1082 (
            .O(N__4982),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    Odrv4 I__1081 (
            .O(N__4979),
            .I(\uart_frame_decoder.state_1Z0Z_10 ));
    IoInMux I__1080 (
            .O(N__4970),
            .I(N__4967));
    LocalMux I__1079 (
            .O(N__4967),
            .I(N__4964));
    Span12Mux_s3_v I__1078 (
            .O(N__4964),
            .I(N__4961));
    Odrv12 I__1077 (
            .O(N__4961),
            .I(uart_frame_decoder_N_306_i));
    InMux I__1076 (
            .O(N__4958),
            .I(\uart_frame_decoder.un1_WDT_cry_14 ));
    CascadeMux I__1075 (
            .O(N__4955),
            .I(N__4950));
    InMux I__1074 (
            .O(N__4954),
            .I(N__4947));
    InMux I__1073 (
            .O(N__4953),
            .I(N__4942));
    InMux I__1072 (
            .O(N__4950),
            .I(N__4942));
    LocalMux I__1071 (
            .O(N__4947),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    LocalMux I__1070 (
            .O(N__4942),
            .I(\uart_frame_decoder.WDTZ0Z_15 ));
    InMux I__1069 (
            .O(N__4937),
            .I(N__4934));
    LocalMux I__1068 (
            .O(N__4934),
            .I(N__4931));
    Odrv4 I__1067 (
            .O(N__4931),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10 ));
    InMux I__1066 (
            .O(N__4928),
            .I(N__4924));
    InMux I__1065 (
            .O(N__4927),
            .I(N__4921));
    LocalMux I__1064 (
            .O(N__4924),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_d_10 ));
    LocalMux I__1063 (
            .O(N__4921),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_d_10 ));
    InMux I__1062 (
            .O(N__4916),
            .I(N__4893));
    InMux I__1061 (
            .O(N__4915),
            .I(N__4893));
    InMux I__1060 (
            .O(N__4914),
            .I(N__4893));
    InMux I__1059 (
            .O(N__4913),
            .I(N__4893));
    InMux I__1058 (
            .O(N__4912),
            .I(N__4893));
    InMux I__1057 (
            .O(N__4911),
            .I(N__4893));
    InMux I__1056 (
            .O(N__4910),
            .I(N__4893));
    InMux I__1055 (
            .O(N__4909),
            .I(N__4888));
    InMux I__1054 (
            .O(N__4908),
            .I(N__4888));
    LocalMux I__1053 (
            .O(N__4893),
            .I(\uart_frame_decoder.N_85 ));
    LocalMux I__1052 (
            .O(N__4888),
            .I(\uart_frame_decoder.N_85 ));
    ClkMux I__1051 (
            .O(N__4883),
            .I(N__4808));
    ClkMux I__1050 (
            .O(N__4882),
            .I(N__4808));
    ClkMux I__1049 (
            .O(N__4881),
            .I(N__4808));
    ClkMux I__1048 (
            .O(N__4880),
            .I(N__4808));
    ClkMux I__1047 (
            .O(N__4879),
            .I(N__4808));
    ClkMux I__1046 (
            .O(N__4878),
            .I(N__4808));
    ClkMux I__1045 (
            .O(N__4877),
            .I(N__4808));
    ClkMux I__1044 (
            .O(N__4876),
            .I(N__4808));
    ClkMux I__1043 (
            .O(N__4875),
            .I(N__4808));
    ClkMux I__1042 (
            .O(N__4874),
            .I(N__4808));
    ClkMux I__1041 (
            .O(N__4873),
            .I(N__4808));
    ClkMux I__1040 (
            .O(N__4872),
            .I(N__4808));
    ClkMux I__1039 (
            .O(N__4871),
            .I(N__4808));
    ClkMux I__1038 (
            .O(N__4870),
            .I(N__4808));
    ClkMux I__1037 (
            .O(N__4869),
            .I(N__4808));
    ClkMux I__1036 (
            .O(N__4868),
            .I(N__4808));
    ClkMux I__1035 (
            .O(N__4867),
            .I(N__4808));
    ClkMux I__1034 (
            .O(N__4866),
            .I(N__4808));
    ClkMux I__1033 (
            .O(N__4865),
            .I(N__4808));
    ClkMux I__1032 (
            .O(N__4864),
            .I(N__4808));
    ClkMux I__1031 (
            .O(N__4863),
            .I(N__4808));
    ClkMux I__1030 (
            .O(N__4862),
            .I(N__4808));
    ClkMux I__1029 (
            .O(N__4861),
            .I(N__4808));
    ClkMux I__1028 (
            .O(N__4860),
            .I(N__4808));
    ClkMux I__1027 (
            .O(N__4859),
            .I(N__4808));
    GlobalMux I__1026 (
            .O(N__4808),
            .I(N__4805));
    gio2CtrlBuf I__1025 (
            .O(N__4805),
            .I(clk_system_c_g));
    InMux I__1024 (
            .O(N__4802),
            .I(N__4797));
    InMux I__1023 (
            .O(N__4801),
            .I(N__4794));
    InMux I__1022 (
            .O(N__4800),
            .I(N__4791));
    LocalMux I__1021 (
            .O(N__4797),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__1020 (
            .O(N__4794),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__1019 (
            .O(N__4791),
            .I(\uart_frame_decoder.WDTZ0Z_7 ));
    InMux I__1018 (
            .O(N__4784),
            .I(\uart_frame_decoder.un1_WDT_cry_6 ));
    CascadeMux I__1017 (
            .O(N__4781),
            .I(N__4776));
    InMux I__1016 (
            .O(N__4780),
            .I(N__4773));
    InMux I__1015 (
            .O(N__4779),
            .I(N__4770));
    InMux I__1014 (
            .O(N__4776),
            .I(N__4767));
    LocalMux I__1013 (
            .O(N__4773),
            .I(N__4764));
    LocalMux I__1012 (
            .O(N__4770),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__1011 (
            .O(N__4767),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    Odrv4 I__1010 (
            .O(N__4764),
            .I(\uart_frame_decoder.WDTZ0Z_8 ));
    InMux I__1009 (
            .O(N__4757),
            .I(bfn_12_3_0_));
    InMux I__1008 (
            .O(N__4754),
            .I(N__4749));
    InMux I__1007 (
            .O(N__4753),
            .I(N__4746));
    InMux I__1006 (
            .O(N__4752),
            .I(N__4743));
    LocalMux I__1005 (
            .O(N__4749),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__1004 (
            .O(N__4746),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__1003 (
            .O(N__4743),
            .I(\uart_frame_decoder.WDTZ0Z_9 ));
    InMux I__1002 (
            .O(N__4736),
            .I(\uart_frame_decoder.un1_WDT_cry_8 ));
    CascadeMux I__1001 (
            .O(N__4733),
            .I(N__4728));
    InMux I__1000 (
            .O(N__4732),
            .I(N__4724));
    InMux I__999 (
            .O(N__4731),
            .I(N__4719));
    InMux I__998 (
            .O(N__4728),
            .I(N__4719));
    InMux I__997 (
            .O(N__4727),
            .I(N__4716));
    LocalMux I__996 (
            .O(N__4724),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__995 (
            .O(N__4719),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__994 (
            .O(N__4716),
            .I(\uart_frame_decoder.WDTZ0Z_10 ));
    InMux I__993 (
            .O(N__4709),
            .I(\uart_frame_decoder.un1_WDT_cry_9 ));
    InMux I__992 (
            .O(N__4706),
            .I(N__4701));
    InMux I__991 (
            .O(N__4705),
            .I(N__4698));
    InMux I__990 (
            .O(N__4704),
            .I(N__4695));
    LocalMux I__989 (
            .O(N__4701),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__988 (
            .O(N__4698),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__987 (
            .O(N__4695),
            .I(\uart_frame_decoder.WDTZ0Z_11 ));
    InMux I__986 (
            .O(N__4688),
            .I(\uart_frame_decoder.un1_WDT_cry_10 ));
    InMux I__985 (
            .O(N__4685),
            .I(N__4680));
    InMux I__984 (
            .O(N__4684),
            .I(N__4677));
    InMux I__983 (
            .O(N__4683),
            .I(N__4674));
    LocalMux I__982 (
            .O(N__4680),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__981 (
            .O(N__4677),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__980 (
            .O(N__4674),
            .I(\uart_frame_decoder.WDTZ0Z_12 ));
    InMux I__979 (
            .O(N__4667),
            .I(\uart_frame_decoder.un1_WDT_cry_11 ));
    CascadeMux I__978 (
            .O(N__4664),
            .I(N__4658));
    InMux I__977 (
            .O(N__4663),
            .I(N__4655));
    InMux I__976 (
            .O(N__4662),
            .I(N__4648));
    InMux I__975 (
            .O(N__4661),
            .I(N__4648));
    InMux I__974 (
            .O(N__4658),
            .I(N__4648));
    LocalMux I__973 (
            .O(N__4655),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__972 (
            .O(N__4648),
            .I(\uart_frame_decoder.WDTZ0Z_13 ));
    InMux I__971 (
            .O(N__4643),
            .I(\uart_frame_decoder.un1_WDT_cry_12 ));
    InMux I__970 (
            .O(N__4640),
            .I(N__4634));
    InMux I__969 (
            .O(N__4639),
            .I(N__4634));
    LocalMux I__968 (
            .O(N__4634),
            .I(N__4627));
    InMux I__967 (
            .O(N__4633),
            .I(N__4624));
    InMux I__966 (
            .O(N__4632),
            .I(N__4617));
    InMux I__965 (
            .O(N__4631),
            .I(N__4617));
    InMux I__964 (
            .O(N__4630),
            .I(N__4617));
    Span4Mux_s1_v I__963 (
            .O(N__4627),
            .I(N__4614));
    LocalMux I__962 (
            .O(N__4624),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__961 (
            .O(N__4617),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    Odrv4 I__960 (
            .O(N__4614),
            .I(\uart_frame_decoder.WDTZ0Z_14 ));
    InMux I__959 (
            .O(N__4607),
            .I(\uart_frame_decoder.un1_WDT_cry_13 ));
    InMux I__958 (
            .O(N__4604),
            .I(N__4601));
    LocalMux I__957 (
            .O(N__4601),
            .I(N__4597));
    CascadeMux I__956 (
            .O(N__4600),
            .I(N__4594));
    Span4Mux_h I__955 (
            .O(N__4597),
            .I(N__4591));
    InMux I__954 (
            .O(N__4594),
            .I(N__4588));
    Odrv4 I__953 (
            .O(N__4591),
            .I(\uart.data_AuxZ0Z_4 ));
    LocalMux I__952 (
            .O(N__4588),
            .I(\uart.data_AuxZ0Z_4 ));
    InMux I__951 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__950 (
            .O(N__4580),
            .I(N__4577));
    Odrv4 I__949 (
            .O(N__4577),
            .I(uart_data_4));
    InMux I__948 (
            .O(N__4574),
            .I(N__4571));
    LocalMux I__947 (
            .O(N__4571),
            .I(N__4567));
    InMux I__946 (
            .O(N__4570),
            .I(N__4564));
    Odrv12 I__945 (
            .O(N__4567),
            .I(\uart.data_AuxZ0Z_6 ));
    LocalMux I__944 (
            .O(N__4564),
            .I(\uart.data_AuxZ0Z_6 ));
    InMux I__943 (
            .O(N__4559),
            .I(N__4556));
    LocalMux I__942 (
            .O(N__4556),
            .I(N__4553));
    Span4Mux_s2_v I__941 (
            .O(N__4553),
            .I(N__4550));
    Odrv4 I__940 (
            .O(N__4550),
            .I(uart_data_6));
    CEMux I__939 (
            .O(N__4547),
            .I(N__4543));
    CEMux I__938 (
            .O(N__4546),
            .I(N__4540));
    LocalMux I__937 (
            .O(N__4543),
            .I(N__4537));
    LocalMux I__936 (
            .O(N__4540),
            .I(N__4534));
    Odrv4 I__935 (
            .O(N__4537),
            .I(\uart.state_1_sqmuxa_0 ));
    Odrv4 I__934 (
            .O(N__4534),
            .I(\uart.state_1_sqmuxa_0 ));
    SRMux I__933 (
            .O(N__4529),
            .I(N__4525));
    SRMux I__932 (
            .O(N__4528),
            .I(N__4522));
    LocalMux I__931 (
            .O(N__4525),
            .I(N__4519));
    LocalMux I__930 (
            .O(N__4522),
            .I(N__4516));
    Span4Mux_s3_v I__929 (
            .O(N__4519),
            .I(N__4512));
    Span4Mux_h I__928 (
            .O(N__4516),
            .I(N__4509));
    InMux I__927 (
            .O(N__4515),
            .I(N__4506));
    Odrv4 I__926 (
            .O(N__4512),
            .I(\uart.timer_Count_RNIS4183Z0Z_7 ));
    Odrv4 I__925 (
            .O(N__4509),
            .I(\uart.timer_Count_RNIS4183Z0Z_7 ));
    LocalMux I__924 (
            .O(N__4506),
            .I(\uart.timer_Count_RNIS4183Z0Z_7 ));
    InMux I__923 (
            .O(N__4499),
            .I(N__4495));
    CascadeMux I__922 (
            .O(N__4498),
            .I(N__4492));
    LocalMux I__921 (
            .O(N__4495),
            .I(N__4489));
    InMux I__920 (
            .O(N__4492),
            .I(N__4486));
    Odrv4 I__919 (
            .O(N__4489),
            .I(\uart_frame_decoder.WDT8_0_i ));
    LocalMux I__918 (
            .O(N__4486),
            .I(\uart_frame_decoder.WDT8_0_i ));
    InMux I__917 (
            .O(N__4481),
            .I(N__4478));
    LocalMux I__916 (
            .O(N__4478),
            .I(\uart_frame_decoder.WDTZ0Z_0 ));
    InMux I__915 (
            .O(N__4475),
            .I(N__4472));
    LocalMux I__914 (
            .O(N__4472),
            .I(\uart_frame_decoder.WDTZ0Z_1 ));
    InMux I__913 (
            .O(N__4469),
            .I(\uart_frame_decoder.un1_WDT_cry_0 ));
    InMux I__912 (
            .O(N__4466),
            .I(N__4463));
    LocalMux I__911 (
            .O(N__4463),
            .I(\uart_frame_decoder.WDTZ0Z_2 ));
    InMux I__910 (
            .O(N__4460),
            .I(\uart_frame_decoder.un1_WDT_cry_1 ));
    InMux I__909 (
            .O(N__4457),
            .I(N__4454));
    LocalMux I__908 (
            .O(N__4454),
            .I(\uart_frame_decoder.WDTZ0Z_3 ));
    InMux I__907 (
            .O(N__4451),
            .I(\uart_frame_decoder.un1_WDT_cry_2 ));
    InMux I__906 (
            .O(N__4448),
            .I(N__4443));
    InMux I__905 (
            .O(N__4447),
            .I(N__4438));
    InMux I__904 (
            .O(N__4446),
            .I(N__4438));
    LocalMux I__903 (
            .O(N__4443),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__902 (
            .O(N__4438),
            .I(\uart_frame_decoder.WDTZ0Z_4 ));
    InMux I__901 (
            .O(N__4433),
            .I(\uart_frame_decoder.un1_WDT_cry_3 ));
    CascadeMux I__900 (
            .O(N__4430),
            .I(N__4427));
    InMux I__899 (
            .O(N__4427),
            .I(N__4422));
    InMux I__898 (
            .O(N__4426),
            .I(N__4419));
    InMux I__897 (
            .O(N__4425),
            .I(N__4416));
    LocalMux I__896 (
            .O(N__4422),
            .I(N__4413));
    LocalMux I__895 (
            .O(N__4419),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__894 (
            .O(N__4416),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    Odrv4 I__893 (
            .O(N__4413),
            .I(\uart_frame_decoder.WDTZ0Z_5 ));
    InMux I__892 (
            .O(N__4406),
            .I(\uart_frame_decoder.un1_WDT_cry_4 ));
    CascadeMux I__891 (
            .O(N__4403),
            .I(N__4398));
    InMux I__890 (
            .O(N__4402),
            .I(N__4395));
    InMux I__889 (
            .O(N__4401),
            .I(N__4392));
    InMux I__888 (
            .O(N__4398),
            .I(N__4389));
    LocalMux I__887 (
            .O(N__4395),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__886 (
            .O(N__4392),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__885 (
            .O(N__4389),
            .I(\uart_frame_decoder.WDTZ0Z_6 ));
    InMux I__884 (
            .O(N__4382),
            .I(\uart_frame_decoder.un1_WDT_cry_5 ));
    InMux I__883 (
            .O(N__4379),
            .I(N__4376));
    LocalMux I__882 (
            .O(N__4376),
            .I(\uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ));
    CascadeMux I__881 (
            .O(N__4373),
            .I(\uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_ ));
    CascadeMux I__880 (
            .O(N__4370),
            .I(\uart_frame_decoder.WDT8lt13_cascade_ ));
    InMux I__879 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__878 (
            .O(N__4364),
            .I(\uart_frame_decoder.state_1_ns_i_i_a2_0_0 ));
    CascadeMux I__877 (
            .O(N__4361),
            .I(N__4358));
    InMux I__876 (
            .O(N__4358),
            .I(N__4352));
    InMux I__875 (
            .O(N__4357),
            .I(N__4352));
    LocalMux I__874 (
            .O(N__4352),
            .I(\uart_frame_decoder.WDT8lt13 ));
    CascadeMux I__873 (
            .O(N__4349),
            .I(N__4346));
    InMux I__872 (
            .O(N__4346),
            .I(N__4342));
    InMux I__871 (
            .O(N__4345),
            .I(N__4339));
    LocalMux I__870 (
            .O(N__4342),
            .I(\uart_frame_decoder.WDT8lto15 ));
    LocalMux I__869 (
            .O(N__4339),
            .I(\uart_frame_decoder.WDT8lto15 ));
    InMux I__868 (
            .O(N__4334),
            .I(N__4331));
    LocalMux I__867 (
            .O(N__4331),
            .I(\uart_frame_decoder.N_80 ));
    CascadeMux I__866 (
            .O(N__4328),
            .I(N__4325));
    InMux I__865 (
            .O(N__4325),
            .I(N__4321));
    InMux I__864 (
            .O(N__4324),
            .I(N__4316));
    LocalMux I__863 (
            .O(N__4321),
            .I(N__4313));
    InMux I__862 (
            .O(N__4320),
            .I(N__4308));
    InMux I__861 (
            .O(N__4319),
            .I(N__4308));
    LocalMux I__860 (
            .O(N__4316),
            .I(N__4305));
    Span4Mux_h I__859 (
            .O(N__4313),
            .I(N__4302));
    LocalMux I__858 (
            .O(N__4308),
            .I(\uart.timer_CountZ0Z_0 ));
    Odrv4 I__857 (
            .O(N__4305),
            .I(\uart.timer_CountZ0Z_0 ));
    Odrv4 I__856 (
            .O(N__4302),
            .I(\uart.timer_CountZ0Z_0 ));
    SRMux I__855 (
            .O(N__4295),
            .I(N__4291));
    SRMux I__854 (
            .O(N__4294),
            .I(N__4288));
    LocalMux I__853 (
            .O(N__4291),
            .I(\uart.timer_Count_1_sqmuxa_i ));
    LocalMux I__852 (
            .O(N__4288),
            .I(\uart.timer_Count_1_sqmuxa_i ));
    CascadeMux I__851 (
            .O(N__4283),
            .I(N__4280));
    InMux I__850 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__849 (
            .O(N__4277),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ));
    CascadeMux I__848 (
            .O(N__4274),
            .I(N__4271));
    InMux I__847 (
            .O(N__4271),
            .I(N__4264));
    InMux I__846 (
            .O(N__4270),
            .I(N__4264));
    InMux I__845 (
            .O(N__4269),
            .I(N__4261));
    LocalMux I__844 (
            .O(N__4264),
            .I(\uart_frame_decoder.N_99 ));
    LocalMux I__843 (
            .O(N__4261),
            .I(\uart_frame_decoder.N_99 ));
    InMux I__842 (
            .O(N__4256),
            .I(N__4252));
    InMux I__841 (
            .O(N__4255),
            .I(N__4249));
    LocalMux I__840 (
            .O(N__4252),
            .I(\uart_frame_decoder.N_92 ));
    LocalMux I__839 (
            .O(N__4249),
            .I(\uart_frame_decoder.N_92 ));
    InMux I__838 (
            .O(N__4244),
            .I(N__4241));
    LocalMux I__837 (
            .O(N__4241),
            .I(N__4237));
    CascadeMux I__836 (
            .O(N__4240),
            .I(N__4234));
    Span4Mux_v I__835 (
            .O(N__4237),
            .I(N__4231));
    InMux I__834 (
            .O(N__4234),
            .I(N__4228));
    Odrv4 I__833 (
            .O(N__4231),
            .I(\uart.data_AuxZ0Z_1 ));
    LocalMux I__832 (
            .O(N__4228),
            .I(\uart.data_AuxZ0Z_1 ));
    InMux I__831 (
            .O(N__4223),
            .I(N__4220));
    LocalMux I__830 (
            .O(N__4220),
            .I(N__4217));
    Odrv4 I__829 (
            .O(N__4217),
            .I(uart_data_1));
    CascadeMux I__828 (
            .O(N__4214),
            .I(\uart_frame_decoder.N_4_0_cascade_ ));
    InMux I__827 (
            .O(N__4211),
            .I(N__4208));
    LocalMux I__826 (
            .O(N__4208),
            .I(\uart_frame_decoder.g0_1_0_1 ));
    InMux I__825 (
            .O(N__4205),
            .I(N__4202));
    LocalMux I__824 (
            .O(N__4202),
            .I(\uart_frame_decoder.g0_1_a3_3 ));
    CascadeMux I__823 (
            .O(N__4199),
            .I(\uart_frame_decoder.WDT8lto15_cascade_ ));
    InMux I__822 (
            .O(N__4196),
            .I(N__4193));
    LocalMux I__821 (
            .O(N__4193),
            .I(\uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10 ));
    InMux I__820 (
            .O(N__4190),
            .I(N__4187));
    LocalMux I__819 (
            .O(N__4187),
            .I(\uart_frame_decoder.state_1_ns_i_i_a2_1_1_0 ));
    InMux I__818 (
            .O(N__4184),
            .I(N__4179));
    InMux I__817 (
            .O(N__4183),
            .I(N__4174));
    InMux I__816 (
            .O(N__4182),
            .I(N__4174));
    LocalMux I__815 (
            .O(N__4179),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    LocalMux I__814 (
            .O(N__4174),
            .I(\uart_frame_decoder.state_1Z0Z_0 ));
    CascadeMux I__813 (
            .O(N__4169),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_ ));
    InMux I__812 (
            .O(N__4166),
            .I(N__4163));
    LocalMux I__811 (
            .O(N__4163),
            .I(\uart_frame_decoder.N_35_i_1 ));
    CascadeMux I__810 (
            .O(N__4160),
            .I(N__4157));
    InMux I__809 (
            .O(N__4157),
            .I(N__4152));
    InMux I__808 (
            .O(N__4156),
            .I(N__4149));
    InMux I__807 (
            .O(N__4155),
            .I(N__4145));
    LocalMux I__806 (
            .O(N__4152),
            .I(N__4142));
    LocalMux I__805 (
            .O(N__4149),
            .I(N__4139));
    InMux I__804 (
            .O(N__4148),
            .I(N__4136));
    LocalMux I__803 (
            .O(N__4145),
            .I(\uart.timer_CountZ0Z_1 ));
    Odrv4 I__802 (
            .O(N__4142),
            .I(\uart.timer_CountZ0Z_1 ));
    Odrv12 I__801 (
            .O(N__4139),
            .I(\uart.timer_CountZ0Z_1 ));
    LocalMux I__800 (
            .O(N__4136),
            .I(\uart.timer_CountZ0Z_1 ));
    CascadeMux I__799 (
            .O(N__4127),
            .I(N__4124));
    InMux I__798 (
            .O(N__4124),
            .I(N__4121));
    LocalMux I__797 (
            .O(N__4121),
            .I(\uart_frame_decoder.count8_axb_1 ));
    CascadeMux I__796 (
            .O(N__4118),
            .I(N__4115));
    InMux I__795 (
            .O(N__4115),
            .I(N__4112));
    LocalMux I__794 (
            .O(N__4112),
            .I(\uart_frame_decoder.count_i_2 ));
    InMux I__793 (
            .O(N__4109),
            .I(\uart_frame_decoder.count8 ));
    InMux I__792 (
            .O(N__4106),
            .I(N__4103));
    LocalMux I__791 (
            .O(N__4103),
            .I(N__4100));
    Odrv12 I__790 (
            .O(N__4100),
            .I(\uart_frame_decoder.count8_THRU_CO ));
    CascadeMux I__789 (
            .O(N__4097),
            .I(\uart_frame_decoder.count8_THRU_CO_cascade_ ));
    InMux I__788 (
            .O(N__4094),
            .I(N__4088));
    InMux I__787 (
            .O(N__4093),
            .I(N__4088));
    LocalMux I__786 (
            .O(N__4088),
            .I(\uart_frame_decoder.N_37 ));
    CascadeMux I__785 (
            .O(N__4085),
            .I(\uart_frame_decoder.N_37_cascade_ ));
    CascadeMux I__784 (
            .O(N__4082),
            .I(N__4077));
    InMux I__783 (
            .O(N__4081),
            .I(N__4071));
    InMux I__782 (
            .O(N__4080),
            .I(N__4071));
    InMux I__781 (
            .O(N__4077),
            .I(N__4066));
    InMux I__780 (
            .O(N__4076),
            .I(N__4066));
    LocalMux I__779 (
            .O(N__4071),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    LocalMux I__778 (
            .O(N__4066),
            .I(\uart_frame_decoder.countZ0Z_1 ));
    InMux I__777 (
            .O(N__4061),
            .I(N__4056));
    InMux I__776 (
            .O(N__4060),
            .I(N__4051));
    InMux I__775 (
            .O(N__4059),
            .I(N__4051));
    LocalMux I__774 (
            .O(N__4056),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    LocalMux I__773 (
            .O(N__4051),
            .I(\uart_frame_decoder.countZ0Z_2 ));
    InMux I__772 (
            .O(N__4046),
            .I(N__4040));
    InMux I__771 (
            .O(N__4045),
            .I(N__4040));
    LocalMux I__770 (
            .O(N__4040),
            .I(CONSTANT_ONE_NET));
    InMux I__769 (
            .O(N__4037),
            .I(N__4031));
    InMux I__768 (
            .O(N__4036),
            .I(N__4024));
    InMux I__767 (
            .O(N__4035),
            .I(N__4024));
    InMux I__766 (
            .O(N__4034),
            .I(N__4024));
    LocalMux I__765 (
            .O(N__4031),
            .I(\uart_frame_decoder.count8_0 ));
    LocalMux I__764 (
            .O(N__4024),
            .I(\uart_frame_decoder.count8_0 ));
    CascadeMux I__763 (
            .O(N__4019),
            .I(N__4015));
    InMux I__762 (
            .O(N__4018),
            .I(N__4010));
    InMux I__761 (
            .O(N__4015),
            .I(N__4010));
    LocalMux I__760 (
            .O(N__4010),
            .I(\uart_frame_decoder.count8_0_i ));
    InMux I__759 (
            .O(N__4007),
            .I(N__4004));
    LocalMux I__758 (
            .O(N__4004),
            .I(N__3997));
    InMux I__757 (
            .O(N__4003),
            .I(N__3994));
    InMux I__756 (
            .O(N__4002),
            .I(N__3987));
    InMux I__755 (
            .O(N__4001),
            .I(N__3987));
    InMux I__754 (
            .O(N__4000),
            .I(N__3987));
    Odrv4 I__753 (
            .O(N__3997),
            .I(\uart.N_145_0 ));
    LocalMux I__752 (
            .O(N__3994),
            .I(\uart.N_145_0 ));
    LocalMux I__751 (
            .O(N__3987),
            .I(\uart.N_145_0 ));
    InMux I__750 (
            .O(N__3980),
            .I(N__3977));
    LocalMux I__749 (
            .O(N__3977),
            .I(\uart.state_1_sqmuxa ));
    CascadeMux I__748 (
            .O(N__3974),
            .I(\uart.state_1_sqmuxa_cascade_ ));
    InMux I__747 (
            .O(N__3971),
            .I(N__3968));
    LocalMux I__746 (
            .O(N__3968),
            .I(N__3961));
    InMux I__745 (
            .O(N__3967),
            .I(N__3958));
    InMux I__744 (
            .O(N__3966),
            .I(N__3955));
    InMux I__743 (
            .O(N__3965),
            .I(N__3952));
    InMux I__742 (
            .O(N__3964),
            .I(N__3949));
    Span4Mux_v I__741 (
            .O(N__3961),
            .I(N__3946));
    LocalMux I__740 (
            .O(N__3958),
            .I(N__3941));
    LocalMux I__739 (
            .O(N__3955),
            .I(N__3941));
    LocalMux I__738 (
            .O(N__3952),
            .I(\uart.timer_CountZ0Z_2 ));
    LocalMux I__737 (
            .O(N__3949),
            .I(\uart.timer_CountZ0Z_2 ));
    Odrv4 I__736 (
            .O(N__3946),
            .I(\uart.timer_CountZ0Z_2 ));
    Odrv4 I__735 (
            .O(N__3941),
            .I(\uart.timer_CountZ0Z_2 ));
    InMux I__734 (
            .O(N__3932),
            .I(\uart.un4_timer_Count_1_cry_1 ));
    InMux I__733 (
            .O(N__3929),
            .I(N__3926));
    LocalMux I__732 (
            .O(N__3926),
            .I(N__3921));
    InMux I__731 (
            .O(N__3925),
            .I(N__3916));
    InMux I__730 (
            .O(N__3924),
            .I(N__3913));
    Span4Mux_h I__729 (
            .O(N__3921),
            .I(N__3910));
    InMux I__728 (
            .O(N__3920),
            .I(N__3907));
    InMux I__727 (
            .O(N__3919),
            .I(N__3904));
    LocalMux I__726 (
            .O(N__3916),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__725 (
            .O(N__3913),
            .I(\uart.timer_CountZ0Z_3 ));
    Odrv4 I__724 (
            .O(N__3910),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__723 (
            .O(N__3907),
            .I(\uart.timer_CountZ0Z_3 ));
    LocalMux I__722 (
            .O(N__3904),
            .I(\uart.timer_CountZ0Z_3 ));
    InMux I__721 (
            .O(N__3893),
            .I(\uart.un4_timer_Count_1_cry_2 ));
    InMux I__720 (
            .O(N__3890),
            .I(N__3887));
    LocalMux I__719 (
            .O(N__3887),
            .I(N__3881));
    CascadeMux I__718 (
            .O(N__3886),
            .I(N__3877));
    InMux I__717 (
            .O(N__3885),
            .I(N__3874));
    InMux I__716 (
            .O(N__3884),
            .I(N__3871));
    Span4Mux_h I__715 (
            .O(N__3881),
            .I(N__3868));
    InMux I__714 (
            .O(N__3880),
            .I(N__3865));
    InMux I__713 (
            .O(N__3877),
            .I(N__3862));
    LocalMux I__712 (
            .O(N__3874),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__711 (
            .O(N__3871),
            .I(\uart.timer_CountZ0Z_4 ));
    Odrv4 I__710 (
            .O(N__3868),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__709 (
            .O(N__3865),
            .I(\uart.timer_CountZ0Z_4 ));
    LocalMux I__708 (
            .O(N__3862),
            .I(\uart.timer_CountZ0Z_4 ));
    InMux I__707 (
            .O(N__3851),
            .I(\uart.un4_timer_Count_1_cry_3 ));
    InMux I__706 (
            .O(N__3848),
            .I(N__3844));
    InMux I__705 (
            .O(N__3847),
            .I(N__3838));
    LocalMux I__704 (
            .O(N__3844),
            .I(N__3835));
    InMux I__703 (
            .O(N__3843),
            .I(N__3828));
    InMux I__702 (
            .O(N__3842),
            .I(N__3828));
    InMux I__701 (
            .O(N__3841),
            .I(N__3828));
    LocalMux I__700 (
            .O(N__3838),
            .I(\uart.timer_CountZ0Z_5 ));
    Odrv4 I__699 (
            .O(N__3835),
            .I(\uart.timer_CountZ0Z_5 ));
    LocalMux I__698 (
            .O(N__3828),
            .I(\uart.timer_CountZ0Z_5 ));
    InMux I__697 (
            .O(N__3821),
            .I(\uart.un4_timer_Count_1_cry_4 ));
    InMux I__696 (
            .O(N__3818),
            .I(N__3814));
    InMux I__695 (
            .O(N__3817),
            .I(N__3809));
    LocalMux I__694 (
            .O(N__3814),
            .I(N__3806));
    InMux I__693 (
            .O(N__3813),
            .I(N__3801));
    InMux I__692 (
            .O(N__3812),
            .I(N__3801));
    LocalMux I__691 (
            .O(N__3809),
            .I(\uart.timer_CountZ0Z_6 ));
    Odrv4 I__690 (
            .O(N__3806),
            .I(\uart.timer_CountZ0Z_6 ));
    LocalMux I__689 (
            .O(N__3801),
            .I(\uart.timer_CountZ0Z_6 ));
    InMux I__688 (
            .O(N__3794),
            .I(\uart.un4_timer_Count_1_cry_5 ));
    InMux I__687 (
            .O(N__3791),
            .I(\uart.un4_timer_Count_1_cry_6 ));
    InMux I__686 (
            .O(N__3788),
            .I(N__3784));
    InMux I__685 (
            .O(N__3787),
            .I(N__3781));
    LocalMux I__684 (
            .O(N__3784),
            .I(N__3774));
    LocalMux I__683 (
            .O(N__3781),
            .I(N__3774));
    CascadeMux I__682 (
            .O(N__3780),
            .I(N__3767));
    InMux I__681 (
            .O(N__3779),
            .I(N__3764));
    Span4Mux_s1_v I__680 (
            .O(N__3774),
            .I(N__3761));
    InMux I__679 (
            .O(N__3773),
            .I(N__3754));
    InMux I__678 (
            .O(N__3772),
            .I(N__3754));
    InMux I__677 (
            .O(N__3771),
            .I(N__3754));
    InMux I__676 (
            .O(N__3770),
            .I(N__3749));
    InMux I__675 (
            .O(N__3767),
            .I(N__3749));
    LocalMux I__674 (
            .O(N__3764),
            .I(\uart.timer_CountZ0Z_7 ));
    Odrv4 I__673 (
            .O(N__3761),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__672 (
            .O(N__3754),
            .I(\uart.timer_CountZ0Z_7 ));
    LocalMux I__671 (
            .O(N__3749),
            .I(\uart.timer_CountZ0Z_7 ));
    InMux I__670 (
            .O(N__3740),
            .I(N__3737));
    LocalMux I__669 (
            .O(N__3737),
            .I(uart_data_3));
    CascadeMux I__668 (
            .O(N__3734),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_ ));
    InMux I__667 (
            .O(N__3731),
            .I(N__3725));
    InMux I__666 (
            .O(N__3730),
            .I(N__3725));
    LocalMux I__665 (
            .O(N__3725),
            .I(uart_data_2));
    InMux I__664 (
            .O(N__3722),
            .I(N__3716));
    InMux I__663 (
            .O(N__3721),
            .I(N__3716));
    LocalMux I__662 (
            .O(N__3716),
            .I(uart_data_5));
    CascadeMux I__661 (
            .O(N__3713),
            .I(N__3710));
    InMux I__660 (
            .O(N__3710),
            .I(N__3704));
    InMux I__659 (
            .O(N__3709),
            .I(N__3704));
    LocalMux I__658 (
            .O(N__3704),
            .I(uart_data_7));
    InMux I__657 (
            .O(N__3701),
            .I(N__3695));
    InMux I__656 (
            .O(N__3700),
            .I(N__3695));
    LocalMux I__655 (
            .O(N__3695),
            .I(uart_data_0));
    InMux I__654 (
            .O(N__3692),
            .I(N__3689));
    LocalMux I__653 (
            .O(N__3689),
            .I(\uart_frame_decoder.N_79_4 ));
    CascadeMux I__652 (
            .O(N__3686),
            .I(\uart_frame_decoder.N_79_4_cascade_ ));
    CascadeMux I__651 (
            .O(N__3683),
            .I(N__3678));
    CascadeMux I__650 (
            .O(N__3682),
            .I(N__3673));
    InMux I__649 (
            .O(N__3681),
            .I(N__3665));
    InMux I__648 (
            .O(N__3678),
            .I(N__3662));
    InMux I__647 (
            .O(N__3677),
            .I(N__3659));
    InMux I__646 (
            .O(N__3676),
            .I(N__3656));
    InMux I__645 (
            .O(N__3673),
            .I(N__3653));
    InMux I__644 (
            .O(N__3672),
            .I(N__3647));
    InMux I__643 (
            .O(N__3671),
            .I(N__3638));
    InMux I__642 (
            .O(N__3670),
            .I(N__3638));
    InMux I__641 (
            .O(N__3669),
            .I(N__3638));
    InMux I__640 (
            .O(N__3668),
            .I(N__3638));
    LocalMux I__639 (
            .O(N__3665),
            .I(N__3635));
    LocalMux I__638 (
            .O(N__3662),
            .I(N__3626));
    LocalMux I__637 (
            .O(N__3659),
            .I(N__3626));
    LocalMux I__636 (
            .O(N__3656),
            .I(N__3626));
    LocalMux I__635 (
            .O(N__3653),
            .I(N__3626));
    InMux I__634 (
            .O(N__3652),
            .I(N__3619));
    InMux I__633 (
            .O(N__3651),
            .I(N__3619));
    InMux I__632 (
            .O(N__3650),
            .I(N__3619));
    LocalMux I__631 (
            .O(N__3647),
            .I(N__3616));
    LocalMux I__630 (
            .O(N__3638),
            .I(N__3613));
    Span4Mux_s1_v I__629 (
            .O(N__3635),
            .I(N__3608));
    Span4Mux_v I__628 (
            .O(N__3626),
            .I(N__3608));
    LocalMux I__627 (
            .O(N__3619),
            .I(uart_input_sync));
    Odrv4 I__626 (
            .O(N__3616),
            .I(uart_input_sync));
    Odrv4 I__625 (
            .O(N__3613),
            .I(uart_input_sync));
    Odrv4 I__624 (
            .O(N__3608),
            .I(uart_input_sync));
    CascadeMux I__623 (
            .O(N__3599),
            .I(\uart.data_8_0_cascade_ ));
    InMux I__622 (
            .O(N__3596),
            .I(N__3593));
    LocalMux I__621 (
            .O(N__3593),
            .I(\uart.state_srsts_0_a3_1_4 ));
    CascadeMux I__620 (
            .O(N__3590),
            .I(\uart.N_152_0_cascade_ ));
    InMux I__619 (
            .O(N__3587),
            .I(N__3584));
    LocalMux I__618 (
            .O(N__3584),
            .I(\uart.N_167 ));
    InMux I__617 (
            .O(N__3581),
            .I(N__3578));
    LocalMux I__616 (
            .O(N__3578),
            .I(\uart.N_159 ));
    CascadeMux I__615 (
            .O(N__3575),
            .I(\uart.N_167_cascade_ ));
    InMux I__614 (
            .O(N__3572),
            .I(N__3568));
    InMux I__613 (
            .O(N__3571),
            .I(N__3562));
    LocalMux I__612 (
            .O(N__3568),
            .I(N__3559));
    InMux I__611 (
            .O(N__3567),
            .I(N__3556));
    InMux I__610 (
            .O(N__3566),
            .I(N__3553));
    InMux I__609 (
            .O(N__3565),
            .I(N__3550));
    LocalMux I__608 (
            .O(N__3562),
            .I(\uart.N_180 ));
    Odrv4 I__607 (
            .O(N__3559),
            .I(\uart.N_180 ));
    LocalMux I__606 (
            .O(N__3556),
            .I(\uart.N_180 ));
    LocalMux I__605 (
            .O(N__3553),
            .I(\uart.N_180 ));
    LocalMux I__604 (
            .O(N__3550),
            .I(\uart.N_180 ));
    InMux I__603 (
            .O(N__3539),
            .I(N__3536));
    LocalMux I__602 (
            .O(N__3536),
            .I(N__3531));
    InMux I__601 (
            .O(N__3535),
            .I(N__3526));
    InMux I__600 (
            .O(N__3534),
            .I(N__3526));
    Odrv4 I__599 (
            .O(N__3531),
            .I(\uart.N_152_0 ));
    LocalMux I__598 (
            .O(N__3526),
            .I(\uart.N_152_0 ));
    InMux I__597 (
            .O(N__3521),
            .I(N__3517));
    InMux I__596 (
            .O(N__3520),
            .I(N__3514));
    LocalMux I__595 (
            .O(N__3517),
            .I(N__3506));
    LocalMux I__594 (
            .O(N__3514),
            .I(N__3506));
    CascadeMux I__593 (
            .O(N__3513),
            .I(N__3502));
    InMux I__592 (
            .O(N__3512),
            .I(N__3497));
    InMux I__591 (
            .O(N__3511),
            .I(N__3494));
    Span4Mux_s1_v I__590 (
            .O(N__3506),
            .I(N__3491));
    InMux I__589 (
            .O(N__3505),
            .I(N__3488));
    InMux I__588 (
            .O(N__3502),
            .I(N__3483));
    InMux I__587 (
            .O(N__3501),
            .I(N__3483));
    InMux I__586 (
            .O(N__3500),
            .I(N__3480));
    LocalMux I__585 (
            .O(N__3497),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__584 (
            .O(N__3494),
            .I(\uart.stateZ0Z_4 ));
    Odrv4 I__583 (
            .O(N__3491),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__582 (
            .O(N__3488),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__581 (
            .O(N__3483),
            .I(\uart.stateZ0Z_4 ));
    LocalMux I__580 (
            .O(N__3480),
            .I(\uart.stateZ0Z_4 ));
    CascadeMux I__579 (
            .O(N__3467),
            .I(\uart_frame_decoder.N_43_cascade_ ));
    CascadeMux I__578 (
            .O(N__3464),
            .I(\uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_ ));
    CascadeMux I__577 (
            .O(N__3461),
            .I(\uart_frame_decoder.N_81_cascade_ ));
    CascadeMux I__576 (
            .O(N__3458),
            .I(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ));
    SRMux I__575 (
            .O(N__3455),
            .I(N__3450));
    SRMux I__574 (
            .O(N__3454),
            .I(N__3447));
    SRMux I__573 (
            .O(N__3453),
            .I(N__3444));
    LocalMux I__572 (
            .O(N__3450),
            .I(N__3439));
    LocalMux I__571 (
            .O(N__3447),
            .I(N__3439));
    LocalMux I__570 (
            .O(N__3444),
            .I(N__3436));
    Span4Mux_v I__569 (
            .O(N__3439),
            .I(N__3433));
    Span4Mux_h I__568 (
            .O(N__3436),
            .I(N__3430));
    Span4Mux_h I__567 (
            .O(N__3433),
            .I(N__3427));
    Odrv4 I__566 (
            .O(N__3430),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    Odrv4 I__565 (
            .O(N__3427),
            .I(\uart.state_RNIAFHLZ0Z_4 ));
    InMux I__564 (
            .O(N__3422),
            .I(N__3417));
    InMux I__563 (
            .O(N__3421),
            .I(N__3412));
    InMux I__562 (
            .O(N__3420),
            .I(N__3412));
    LocalMux I__561 (
            .O(N__3417),
            .I(\uart.stateZ0Z_1 ));
    LocalMux I__560 (
            .O(N__3412),
            .I(\uart.stateZ0Z_1 ));
    CascadeMux I__559 (
            .O(N__3407),
            .I(\uart.N_151_cascade_ ));
    CascadeMux I__558 (
            .O(N__3404),
            .I(N__3400));
    InMux I__557 (
            .O(N__3403),
            .I(N__3397));
    InMux I__556 (
            .O(N__3400),
            .I(N__3393));
    LocalMux I__555 (
            .O(N__3397),
            .I(N__3389));
    InMux I__554 (
            .O(N__3396),
            .I(N__3386));
    LocalMux I__553 (
            .O(N__3393),
            .I(N__3383));
    InMux I__552 (
            .O(N__3392),
            .I(N__3380));
    Odrv12 I__551 (
            .O(N__3389),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__550 (
            .O(N__3386),
            .I(\uart.stateZ0Z_2 ));
    Odrv4 I__549 (
            .O(N__3383),
            .I(\uart.stateZ0Z_2 ));
    LocalMux I__548 (
            .O(N__3380),
            .I(\uart.stateZ0Z_2 ));
    InMux I__547 (
            .O(N__3371),
            .I(N__3366));
    CascadeMux I__546 (
            .O(N__3370),
            .I(N__3363));
    CascadeMux I__545 (
            .O(N__3369),
            .I(N__3357));
    LocalMux I__544 (
            .O(N__3366),
            .I(N__3353));
    InMux I__543 (
            .O(N__3363),
            .I(N__3349));
    InMux I__542 (
            .O(N__3362),
            .I(N__3346));
    InMux I__541 (
            .O(N__3361),
            .I(N__3343));
    InMux I__540 (
            .O(N__3360),
            .I(N__3338));
    InMux I__539 (
            .O(N__3357),
            .I(N__3338));
    InMux I__538 (
            .O(N__3356),
            .I(N__3335));
    Span4Mux_h I__537 (
            .O(N__3353),
            .I(N__3331));
    InMux I__536 (
            .O(N__3352),
            .I(N__3328));
    LocalMux I__535 (
            .O(N__3349),
            .I(N__3317));
    LocalMux I__534 (
            .O(N__3346),
            .I(N__3317));
    LocalMux I__533 (
            .O(N__3343),
            .I(N__3317));
    LocalMux I__532 (
            .O(N__3338),
            .I(N__3317));
    LocalMux I__531 (
            .O(N__3335),
            .I(N__3317));
    InMux I__530 (
            .O(N__3334),
            .I(N__3314));
    Odrv4 I__529 (
            .O(N__3331),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__528 (
            .O(N__3328),
            .I(\uart.stateZ0Z_3 ));
    Odrv4 I__527 (
            .O(N__3317),
            .I(\uart.stateZ0Z_3 ));
    LocalMux I__526 (
            .O(N__3314),
            .I(\uart.stateZ0Z_3 ));
    InMux I__525 (
            .O(N__3305),
            .I(N__3302));
    LocalMux I__524 (
            .O(N__3302),
            .I(N__3299));
    Span4Mux_s1_v I__523 (
            .O(N__3299),
            .I(N__3296));
    Odrv4 I__522 (
            .O(N__3296),
            .I(\uart.state_srsts_i_1_1_3 ));
    CascadeMux I__521 (
            .O(N__3293),
            .I(\uart.N_166_cascade_ ));
    CascadeMux I__520 (
            .O(N__3290),
            .I(\uart.state_srsts_0_1_0_cascade_ ));
    InMux I__519 (
            .O(N__3287),
            .I(N__3284));
    LocalMux I__518 (
            .O(N__3284),
            .I(N__3280));
    InMux I__517 (
            .O(N__3283),
            .I(N__3277));
    Odrv4 I__516 (
            .O(N__3280),
            .I(\uart.stateZ0Z_0 ));
    LocalMux I__515 (
            .O(N__3277),
            .I(\uart.stateZ0Z_0 ));
    CascadeMux I__514 (
            .O(N__3272),
            .I(N__3269));
    InMux I__513 (
            .O(N__3269),
            .I(N__3266));
    LocalMux I__512 (
            .O(N__3266),
            .I(N__3263));
    Odrv4 I__511 (
            .O(N__3263),
            .I(\uart_frame_decoder.N_43 ));
    InMux I__510 (
            .O(N__3260),
            .I(N__3256));
    CascadeMux I__509 (
            .O(N__3259),
            .I(N__3253));
    LocalMux I__508 (
            .O(N__3256),
            .I(N__3250));
    InMux I__507 (
            .O(N__3253),
            .I(N__3247));
    Odrv4 I__506 (
            .O(N__3250),
            .I(\uart.data_AuxZ0Z_7 ));
    LocalMux I__505 (
            .O(N__3247),
            .I(\uart.data_AuxZ0Z_7 ));
    CascadeMux I__504 (
            .O(N__3242),
            .I(\uart.timer_Count10lto5_0_0_cascade_ ));
    InMux I__503 (
            .O(N__3239),
            .I(N__3234));
    InMux I__502 (
            .O(N__3238),
            .I(N__3231));
    InMux I__501 (
            .O(N__3237),
            .I(N__3228));
    LocalMux I__500 (
            .O(N__3234),
            .I(\uart.N_177 ));
    LocalMux I__499 (
            .O(N__3231),
            .I(\uart.N_177 ));
    LocalMux I__498 (
            .O(N__3228),
            .I(\uart.N_177 ));
    CascadeMux I__497 (
            .O(N__3221),
            .I(\uart.N_168_cascade_ ));
    InMux I__496 (
            .O(N__3218),
            .I(N__3214));
    InMux I__495 (
            .O(N__3217),
            .I(N__3211));
    LocalMux I__494 (
            .O(N__3214),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__493 (
            .O(N__3211),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__492 (
            .O(N__3206),
            .I(N__3202));
    InMux I__491 (
            .O(N__3205),
            .I(N__3199));
    LocalMux I__490 (
            .O(N__3202),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__489 (
            .O(N__3199),
            .I(\reset_module_System.countZ0Z_17 ));
    CascadeMux I__488 (
            .O(N__3194),
            .I(\reset_module_System.reset6_3_cascade_ ));
    InMux I__487 (
            .O(N__3191),
            .I(N__3188));
    LocalMux I__486 (
            .O(N__3188),
            .I(\reset_module_System.reset6_13 ));
    InMux I__485 (
            .O(N__3185),
            .I(N__3181));
    InMux I__484 (
            .O(N__3184),
            .I(N__3178));
    LocalMux I__483 (
            .O(N__3181),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__482 (
            .O(N__3178),
            .I(\reset_module_System.countZ0Z_12 ));
    InMux I__481 (
            .O(N__3173),
            .I(N__3167));
    CascadeMux I__480 (
            .O(N__3172),
            .I(N__3164));
    InMux I__479 (
            .O(N__3171),
            .I(N__3161));
    InMux I__478 (
            .O(N__3170),
            .I(N__3158));
    LocalMux I__477 (
            .O(N__3167),
            .I(N__3155));
    InMux I__476 (
            .O(N__3164),
            .I(N__3152));
    LocalMux I__475 (
            .O(N__3161),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__474 (
            .O(N__3158),
            .I(\reset_module_System.countZ0Z_0 ));
    Odrv12 I__473 (
            .O(N__3155),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__472 (
            .O(N__3152),
            .I(\reset_module_System.countZ0Z_0 ));
    CascadeMux I__471 (
            .O(N__3143),
            .I(\reset_module_System.reset6_17_cascade_ ));
    InMux I__470 (
            .O(N__3140),
            .I(N__3137));
    LocalMux I__469 (
            .O(N__3137),
            .I(\reset_module_System.reset6_11 ));
    InMux I__468 (
            .O(N__3134),
            .I(N__3119));
    InMux I__467 (
            .O(N__3133),
            .I(N__3119));
    InMux I__466 (
            .O(N__3132),
            .I(N__3119));
    InMux I__465 (
            .O(N__3131),
            .I(N__3119));
    InMux I__464 (
            .O(N__3130),
            .I(N__3119));
    LocalMux I__463 (
            .O(N__3119),
            .I(\reset_module_System.reset6_19 ));
    CascadeMux I__462 (
            .O(N__3116),
            .I(\uart.N_169_cascade_ ));
    CascadeMux I__461 (
            .O(N__3113),
            .I(\uart.state_srsts_i_1_3_cascade_ ));
    InMux I__460 (
            .O(N__3110),
            .I(N__3106));
    InMux I__459 (
            .O(N__3109),
            .I(N__3103));
    LocalMux I__458 (
            .O(N__3106),
            .I(\uart.data_AuxZ0Z_0 ));
    LocalMux I__457 (
            .O(N__3103),
            .I(\uart.data_AuxZ0Z_0 ));
    InMux I__456 (
            .O(N__3098),
            .I(N__3094));
    CascadeMux I__455 (
            .O(N__3097),
            .I(N__3091));
    LocalMux I__454 (
            .O(N__3094),
            .I(N__3088));
    InMux I__453 (
            .O(N__3091),
            .I(N__3085));
    Odrv4 I__452 (
            .O(N__3088),
            .I(\uart.data_AuxZ0Z_2 ));
    LocalMux I__451 (
            .O(N__3085),
            .I(\uart.data_AuxZ0Z_2 ));
    InMux I__450 (
            .O(N__3080),
            .I(N__3076));
    InMux I__449 (
            .O(N__3079),
            .I(N__3073));
    LocalMux I__448 (
            .O(N__3076),
            .I(N__3070));
    LocalMux I__447 (
            .O(N__3073),
            .I(\uart.data_AuxZ0Z_3 ));
    Odrv4 I__446 (
            .O(N__3070),
            .I(\uart.data_AuxZ0Z_3 ));
    InMux I__445 (
            .O(N__3065),
            .I(N__3062));
    LocalMux I__444 (
            .O(N__3062),
            .I(N__3058));
    InMux I__443 (
            .O(N__3061),
            .I(N__3055));
    Odrv4 I__442 (
            .O(N__3058),
            .I(\uart.data_AuxZ0Z_5 ));
    LocalMux I__441 (
            .O(N__3055),
            .I(\uart.data_AuxZ0Z_5 ));
    InMux I__440 (
            .O(N__3050),
            .I(N__3047));
    LocalMux I__439 (
            .O(N__3047),
            .I(N__3043));
    InMux I__438 (
            .O(N__3046),
            .I(N__3040));
    Odrv4 I__437 (
            .O(N__3043),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__436 (
            .O(N__3040),
            .I(\reset_module_System.countZ0Z_16 ));
    InMux I__435 (
            .O(N__3035),
            .I(N__3031));
    InMux I__434 (
            .O(N__3034),
            .I(N__3028));
    LocalMux I__433 (
            .O(N__3031),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__432 (
            .O(N__3028),
            .I(\reset_module_System.countZ0Z_4 ));
    CascadeMux I__431 (
            .O(N__3023),
            .I(N__3020));
    InMux I__430 (
            .O(N__3020),
            .I(N__3016));
    InMux I__429 (
            .O(N__3019),
            .I(N__3013));
    LocalMux I__428 (
            .O(N__3016),
            .I(N__3010));
    LocalMux I__427 (
            .O(N__3013),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__426 (
            .O(N__3010),
            .I(\reset_module_System.countZ0Z_18 ));
    CascadeMux I__425 (
            .O(N__3005),
            .I(\reset_module_System.reset6_14_cascade_ ));
    InMux I__424 (
            .O(N__3002),
            .I(N__2998));
    InMux I__423 (
            .O(N__3001),
            .I(N__2995));
    LocalMux I__422 (
            .O(N__2998),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__421 (
            .O(N__2995),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__420 (
            .O(N__2990),
            .I(N__2986));
    InMux I__419 (
            .O(N__2989),
            .I(N__2983));
    LocalMux I__418 (
            .O(N__2986),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__417 (
            .O(N__2983),
            .I(\reset_module_System.countZ0Z_3 ));
    CascadeMux I__416 (
            .O(N__2978),
            .I(N__2975));
    InMux I__415 (
            .O(N__2975),
            .I(N__2971));
    InMux I__414 (
            .O(N__2974),
            .I(N__2968));
    LocalMux I__413 (
            .O(N__2971),
            .I(N__2965));
    LocalMux I__412 (
            .O(N__2968),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__411 (
            .O(N__2965),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__410 (
            .O(N__2960),
            .I(N__2956));
    InMux I__409 (
            .O(N__2959),
            .I(N__2953));
    LocalMux I__408 (
            .O(N__2956),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__407 (
            .O(N__2953),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__406 (
            .O(N__2948),
            .I(N__2944));
    InMux I__405 (
            .O(N__2947),
            .I(N__2941));
    LocalMux I__404 (
            .O(N__2944),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__403 (
            .O(N__2941),
            .I(\reset_module_System.countZ0Z_7 ));
    CascadeMux I__402 (
            .O(N__2936),
            .I(N__2932));
    InMux I__401 (
            .O(N__2935),
            .I(N__2929));
    InMux I__400 (
            .O(N__2932),
            .I(N__2926));
    LocalMux I__399 (
            .O(N__2929),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__398 (
            .O(N__2926),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__397 (
            .O(N__2921),
            .I(N__2917));
    InMux I__396 (
            .O(N__2920),
            .I(N__2914));
    LocalMux I__395 (
            .O(N__2917),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__394 (
            .O(N__2914),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__393 (
            .O(N__2909),
            .I(N__2906));
    LocalMux I__392 (
            .O(N__2906),
            .I(N__2903));
    Span4Mux_h I__391 (
            .O(N__2903),
            .I(N__2900));
    Odrv4 I__390 (
            .O(N__2900),
            .I(\reset_module_System.count_1_1 ));
    InMux I__389 (
            .O(N__2897),
            .I(N__2894));
    LocalMux I__388 (
            .O(N__2894),
            .I(N__2889));
    InMux I__387 (
            .O(N__2893),
            .I(N__2886));
    InMux I__386 (
            .O(N__2892),
            .I(N__2883));
    Odrv12 I__385 (
            .O(N__2889),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__384 (
            .O(N__2886),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__383 (
            .O(N__2883),
            .I(\reset_module_System.countZ0Z_1 ));
    CascadeMux I__382 (
            .O(N__2876),
            .I(N__2872));
    CascadeMux I__381 (
            .O(N__2875),
            .I(N__2869));
    InMux I__380 (
            .O(N__2872),
            .I(N__2855));
    InMux I__379 (
            .O(N__2869),
            .I(N__2855));
    InMux I__378 (
            .O(N__2868),
            .I(N__2855));
    InMux I__377 (
            .O(N__2867),
            .I(N__2855));
    InMux I__376 (
            .O(N__2866),
            .I(N__2855));
    LocalMux I__375 (
            .O(N__2855),
            .I(N__2852));
    Span4Mux_h I__374 (
            .O(N__2852),
            .I(N__2849));
    Odrv4 I__373 (
            .O(N__2849),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__372 (
            .O(N__2846),
            .I(N__2843));
    InMux I__371 (
            .O(N__2843),
            .I(N__2831));
    InMux I__370 (
            .O(N__2842),
            .I(N__2831));
    InMux I__369 (
            .O(N__2841),
            .I(N__2831));
    InMux I__368 (
            .O(N__2840),
            .I(N__2831));
    LocalMux I__367 (
            .O(N__2831),
            .I(\reset_module_System.reset6_14 ));
    InMux I__366 (
            .O(N__2828),
            .I(N__2825));
    LocalMux I__365 (
            .O(N__2825),
            .I(\reset_module_System.count_1_2 ));
    CascadeMux I__364 (
            .O(N__2822),
            .I(N__2819));
    InMux I__363 (
            .O(N__2819),
            .I(N__2815));
    InMux I__362 (
            .O(N__2818),
            .I(N__2812));
    LocalMux I__361 (
            .O(N__2815),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__360 (
            .O(N__2812),
            .I(\reset_module_System.countZ0Z_2 ));
    InMux I__359 (
            .O(N__2807),
            .I(N__2803));
    InMux I__358 (
            .O(N__2806),
            .I(N__2800));
    LocalMux I__357 (
            .O(N__2803),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__356 (
            .O(N__2800),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__355 (
            .O(N__2795),
            .I(N__2791));
    InMux I__354 (
            .O(N__2794),
            .I(N__2788));
    LocalMux I__353 (
            .O(N__2791),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__352 (
            .O(N__2788),
            .I(\reset_module_System.countZ0Z_10 ));
    CascadeMux I__351 (
            .O(N__2783),
            .I(N__2778));
    InMux I__350 (
            .O(N__2782),
            .I(N__2771));
    InMux I__349 (
            .O(N__2781),
            .I(N__2764));
    InMux I__348 (
            .O(N__2778),
            .I(N__2764));
    InMux I__347 (
            .O(N__2777),
            .I(N__2764));
    InMux I__346 (
            .O(N__2776),
            .I(N__2757));
    InMux I__345 (
            .O(N__2775),
            .I(N__2757));
    InMux I__344 (
            .O(N__2774),
            .I(N__2757));
    LocalMux I__343 (
            .O(N__2771),
            .I(\uart.un1_state_2_0 ));
    LocalMux I__342 (
            .O(N__2764),
            .I(\uart.un1_state_2_0 ));
    LocalMux I__341 (
            .O(N__2757),
            .I(\uart.un1_state_2_0 ));
    InMux I__340 (
            .O(N__2750),
            .I(N__2747));
    LocalMux I__339 (
            .O(N__2747),
            .I(\uart.data_Auxce_0_0_4 ));
    InMux I__338 (
            .O(N__2744),
            .I(N__2741));
    LocalMux I__337 (
            .O(N__2741),
            .I(\uart.data_Auxce_0_0_0 ));
    InMux I__336 (
            .O(N__2738),
            .I(N__2735));
    LocalMux I__335 (
            .O(N__2735),
            .I(\uart.data_Auxce_0_1 ));
    InMux I__334 (
            .O(N__2732),
            .I(N__2729));
    LocalMux I__333 (
            .O(N__2729),
            .I(N__2726));
    Odrv4 I__332 (
            .O(N__2726),
            .I(\uart.data_Auxce_0_0_2 ));
    InMux I__331 (
            .O(N__2723),
            .I(N__2714));
    InMux I__330 (
            .O(N__2722),
            .I(N__2714));
    InMux I__329 (
            .O(N__2721),
            .I(N__2714));
    LocalMux I__328 (
            .O(N__2714),
            .I(\uart.un1_state_5_0 ));
    CascadeMux I__327 (
            .O(N__2711),
            .I(N__2701));
    CascadeMux I__326 (
            .O(N__2710),
            .I(N__2698));
    InMux I__325 (
            .O(N__2709),
            .I(N__2693));
    InMux I__324 (
            .O(N__2708),
            .I(N__2682));
    InMux I__323 (
            .O(N__2707),
            .I(N__2682));
    InMux I__322 (
            .O(N__2706),
            .I(N__2682));
    InMux I__321 (
            .O(N__2705),
            .I(N__2682));
    InMux I__320 (
            .O(N__2704),
            .I(N__2682));
    InMux I__319 (
            .O(N__2701),
            .I(N__2677));
    InMux I__318 (
            .O(N__2698),
            .I(N__2677));
    InMux I__317 (
            .O(N__2697),
            .I(N__2672));
    InMux I__316 (
            .O(N__2696),
            .I(N__2672));
    LocalMux I__315 (
            .O(N__2693),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__314 (
            .O(N__2682),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__313 (
            .O(N__2677),
            .I(\uart.bit_CountZ0Z_2 ));
    LocalMux I__312 (
            .O(N__2672),
            .I(\uart.bit_CountZ0Z_2 ));
    CascadeMux I__311 (
            .O(N__2663),
            .I(N__2658));
    CascadeMux I__310 (
            .O(N__2662),
            .I(N__2653));
    CascadeMux I__309 (
            .O(N__2661),
            .I(N__2645));
    InMux I__308 (
            .O(N__2658),
            .I(N__2633));
    InMux I__307 (
            .O(N__2657),
            .I(N__2633));
    InMux I__306 (
            .O(N__2656),
            .I(N__2633));
    InMux I__305 (
            .O(N__2653),
            .I(N__2633));
    InMux I__304 (
            .O(N__2652),
            .I(N__2633));
    InMux I__303 (
            .O(N__2651),
            .I(N__2628));
    InMux I__302 (
            .O(N__2650),
            .I(N__2628));
    InMux I__301 (
            .O(N__2649),
            .I(N__2623));
    InMux I__300 (
            .O(N__2648),
            .I(N__2623));
    InMux I__299 (
            .O(N__2645),
            .I(N__2618));
    InMux I__298 (
            .O(N__2644),
            .I(N__2618));
    LocalMux I__297 (
            .O(N__2633),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__296 (
            .O(N__2628),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__295 (
            .O(N__2623),
            .I(\uart.bit_CountZ0Z_1 ));
    LocalMux I__294 (
            .O(N__2618),
            .I(\uart.bit_CountZ0Z_1 ));
    InMux I__293 (
            .O(N__2609),
            .I(N__2587));
    InMux I__292 (
            .O(N__2608),
            .I(N__2587));
    InMux I__291 (
            .O(N__2607),
            .I(N__2587));
    InMux I__290 (
            .O(N__2606),
            .I(N__2587));
    InMux I__289 (
            .O(N__2605),
            .I(N__2587));
    InMux I__288 (
            .O(N__2604),
            .I(N__2582));
    InMux I__287 (
            .O(N__2603),
            .I(N__2582));
    InMux I__286 (
            .O(N__2602),
            .I(N__2575));
    InMux I__285 (
            .O(N__2601),
            .I(N__2575));
    InMux I__284 (
            .O(N__2600),
            .I(N__2575));
    InMux I__283 (
            .O(N__2599),
            .I(N__2570));
    InMux I__282 (
            .O(N__2598),
            .I(N__2570));
    LocalMux I__281 (
            .O(N__2587),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__280 (
            .O(N__2582),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__279 (
            .O(N__2575),
            .I(\uart.bit_CountZ0Z_0 ));
    LocalMux I__278 (
            .O(N__2570),
            .I(\uart.bit_CountZ0Z_0 ));
    CascadeMux I__277 (
            .O(N__2561),
            .I(N__2558));
    InMux I__276 (
            .O(N__2558),
            .I(N__2555));
    LocalMux I__275 (
            .O(N__2555),
            .I(\uart.data_Auxce_0_3 ));
    InMux I__274 (
            .O(N__2552),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__273 (
            .O(N__2549),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__272 (
            .O(N__2546),
            .I(\reset_module_System.count_1_cry_20 ));
    CascadeMux I__271 (
            .O(N__2543),
            .I(N__2539));
    InMux I__270 (
            .O(N__2542),
            .I(N__2536));
    InMux I__269 (
            .O(N__2539),
            .I(N__2533));
    LocalMux I__268 (
            .O(N__2536),
            .I(\reset_module_System.countZ0Z_21 ));
    LocalMux I__267 (
            .O(N__2533),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__266 (
            .O(N__2528),
            .I(N__2525));
    LocalMux I__265 (
            .O(N__2525),
            .I(\uart.data_Auxce_0_5 ));
    InMux I__264 (
            .O(N__2522),
            .I(N__2519));
    LocalMux I__263 (
            .O(N__2519),
            .I(N__2516));
    Odrv4 I__262 (
            .O(N__2516),
            .I(\uart.timer_Count_RNI9M0NZ0Z_1 ));
    CascadeMux I__261 (
            .O(N__2513),
            .I(\uart.timer_Count_RNILKMA1Z0Z_0_cascade_ ));
    CascadeMux I__260 (
            .O(N__2510),
            .I(\uart.un1_state_2_0_cascade_ ));
    InMux I__259 (
            .O(N__2507),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__258 (
            .O(N__2504),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__257 (
            .O(N__2501),
            .I(N__2497));
    InMux I__256 (
            .O(N__2500),
            .I(N__2494));
    LocalMux I__255 (
            .O(N__2497),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__254 (
            .O(N__2494),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__253 (
            .O(N__2489),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__252 (
            .O(N__2486),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__251 (
            .O(N__2483),
            .I(N__2479));
    InMux I__250 (
            .O(N__2482),
            .I(N__2476));
    LocalMux I__249 (
            .O(N__2479),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__248 (
            .O(N__2476),
            .I(\reset_module_System.countZ0Z_15 ));
    InMux I__247 (
            .O(N__2471),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__246 (
            .O(N__2468),
            .I(\reset_module_System.count_1_cry_15 ));
    InMux I__245 (
            .O(N__2465),
            .I(bfn_8_3_0_));
    InMux I__244 (
            .O(N__2462),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__243 (
            .O(N__2459),
            .I(N__2455));
    InMux I__242 (
            .O(N__2458),
            .I(N__2452));
    LocalMux I__241 (
            .O(N__2455),
            .I(\reset_module_System.countZ0Z_19 ));
    LocalMux I__240 (
            .O(N__2452),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__239 (
            .O(N__2447),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__238 (
            .O(N__2444),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__237 (
            .O(N__2441),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__236 (
            .O(N__2438),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__235 (
            .O(N__2435),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__234 (
            .O(N__2432),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__233 (
            .O(N__2429),
            .I(\reset_module_System.count_1_cry_7 ));
    InMux I__232 (
            .O(N__2426),
            .I(bfn_8_2_0_));
    InMux I__231 (
            .O(N__2423),
            .I(\reset_module_System.count_1_cry_9 ));
    CascadeMux I__230 (
            .O(N__2420),
            .I(\uart.N_133_0_cascade_ ));
    InMux I__229 (
            .O(N__2417),
            .I(N__2413));
    InMux I__228 (
            .O(N__2416),
            .I(N__2410));
    LocalMux I__227 (
            .O(N__2413),
            .I(\uart.N_133_0 ));
    LocalMux I__226 (
            .O(N__2410),
            .I(\uart.N_133_0 ));
    CascadeMux I__225 (
            .O(N__2405),
            .I(\uart.data_Auxce_0_6_cascade_ ));
    InMux I__224 (
            .O(N__2402),
            .I(N__2399));
    LocalMux I__223 (
            .O(N__2399),
            .I(N__2396));
    Odrv4 I__222 (
            .O(N__2396),
            .I(\uart.CO1_0 ));
    IoInMux I__221 (
            .O(N__2393),
            .I(N__2390));
    LocalMux I__220 (
            .O(N__2390),
            .I(N__2387));
    Span4Mux_s0_v I__219 (
            .O(N__2387),
            .I(N__2384));
    Sp12to4 I__218 (
            .O(N__2384),
            .I(N__2380));
    CascadeMux I__217 (
            .O(N__2383),
            .I(N__2377));
    Span12Mux_h I__216 (
            .O(N__2380),
            .I(N__2374));
    InMux I__215 (
            .O(N__2377),
            .I(N__2371));
    Odrv12 I__214 (
            .O(N__2374),
            .I(frame_decoder_dv_c));
    LocalMux I__213 (
            .O(N__2371),
            .I(frame_decoder_dv_c));
    InMux I__212 (
            .O(N__2366),
            .I(N__2362));
    IoInMux I__211 (
            .O(N__2365),
            .I(N__2359));
    LocalMux I__210 (
            .O(N__2362),
            .I(N__2356));
    LocalMux I__209 (
            .O(N__2359),
            .I(N__2353));
    Span4Mux_h I__208 (
            .O(N__2356),
            .I(N__2350));
    IoSpan4Mux I__207 (
            .O(N__2353),
            .I(N__2347));
    Odrv4 I__206 (
            .O(N__2350),
            .I(uart_input_c));
    Odrv4 I__205 (
            .O(N__2347),
            .I(uart_input_c));
    InMux I__204 (
            .O(N__2342),
            .I(N__2339));
    LocalMux I__203 (
            .O(N__2339),
            .I(\uart_sync.aux_0__0_Z0Z_0 ));
    InMux I__202 (
            .O(N__2336),
            .I(N__2333));
    LocalMux I__201 (
            .O(N__2333),
            .I(\uart_sync.aux_1__0_Z0Z_0 ));
    InMux I__200 (
            .O(N__2330),
            .I(N__2327));
    LocalMux I__199 (
            .O(N__2327),
            .I(\uart_sync.aux_2__0_Z0Z_0 ));
    InMux I__198 (
            .O(N__2324),
            .I(N__2321));
    LocalMux I__197 (
            .O(N__2321),
            .I(\uart_sync.aux_3__0_Z0Z_0 ));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(\uart_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_12_3_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_5_1_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_5_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__3173),
            .in2(_gnd_net_),
            .in3(N__2897),
            .lcout(\reset_module_System.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.source_data_valid_LC_7_1_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.source_data_valid_LC_7_1_2 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \uart_frame_decoder.source_data_valid_LC_7_1_2  (
            .in0(N__5033),
            .in1(N__5501),
            .in2(N__2383),
            .in3(N__4106),
            .lcout(frame_decoder_dv_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4883),
            .ce(),
            .sr(N__5551));
    defparam \uart_sync.aux_2__0__0_LC_7_2_0 .C_ON=1'b0;
    defparam \uart_sync.aux_2__0__0_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_2__0__0_LC_7_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_2__0__0_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2336),
            .lcout(\uart_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4881),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.aux_0__0__0_LC_7_2_1 .C_ON=1'b0;
    defparam \uart_sync.aux_0__0__0_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_0__0__0_LC_7_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_0__0__0_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2366),
            .lcout(\uart_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4881),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.Q_0__0_LC_7_2_2 .C_ON=1'b0;
    defparam \uart_sync.Q_0__0_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_sync.Q_0__0_LC_7_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.Q_0__0_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2324),
            .lcout(uart_input_sync),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4881),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.aux_1__0__0_LC_7_2_4 .C_ON=1'b0;
    defparam \uart_sync.aux_1__0__0_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_1__0__0_LC_7_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_1__0__0_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2342),
            .lcout(\uart_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4881),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_sync.aux_3__0__0_LC_7_2_5 .C_ON=1'b0;
    defparam \uart_sync.aux_3__0__0_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_sync.aux_3__0__0_LC_7_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_sync.aux_3__0__0_LC_7_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2330),
            .lcout(\uart_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4881),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_7_2_7 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_7_2_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_7_2_7  (
            .in0(N__2458),
            .in1(N__2483),
            .in2(N__2543),
            .in3(N__2501),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_5_LC_7_3_1 .C_ON=1'b0;
    defparam \uart.data_Aux_5_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_5_LC_7_3_1 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \uart.data_Aux_5_LC_7_3_1  (
            .in0(N__3650),
            .in1(N__3061),
            .in2(N__2783),
            .in3(N__2528),
            .lcout(\uart.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4878),
            .ce(),
            .sr(N__3455));
    defparam \uart.data_Aux_7_LC_7_3_2 .C_ON=1'b0;
    defparam \uart.data_Aux_7_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_7_LC_7_3_2 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \uart.data_Aux_7_LC_7_3_2  (
            .in0(N__3238),
            .in1(N__2781),
            .in2(N__3259),
            .in3(N__3652),
            .lcout(\uart.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4878),
            .ce(),
            .sr(N__3455));
    defparam \uart.data_Aux_2_LC_7_3_4 .C_ON=1'b0;
    defparam \uart.data_Aux_2_LC_7_3_4 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_2_LC_7_3_4 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \uart.data_Aux_2_LC_7_3_4  (
            .in0(N__2732),
            .in1(N__2777),
            .in2(N__3097),
            .in3(N__3651),
            .lcout(\uart.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4878),
            .ce(),
            .sr(N__3455));
    defparam \uart.bit_Count_0_LC_7_4_2 .C_ON=1'b0;
    defparam \uart.bit_Count_0_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_0_LC_7_4_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \uart.bit_Count_0_LC_7_4_2  (
            .in0(N__2601),
            .in1(N__2416),
            .in2(_gnd_net_),
            .in3(N__2721),
            .lcout(\uart.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4875),
            .ce(),
            .sr(N__5550));
    defparam \uart.state_RNI4ENK_3_LC_7_4_3 .C_ON=1'b0;
    defparam \uart.state_RNI4ENK_3_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNI4ENK_3_LC_7_4_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \uart.state_RNI4ENK_3_LC_7_4_3  (
            .in0(N__2648),
            .in1(N__3371),
            .in2(N__2710),
            .in3(N__2600),
            .lcout(\uart.N_133_0 ),
            .ltout(\uart.N_133_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_1_LC_7_4_4 .C_ON=1'b0;
    defparam \uart.bit_Count_1_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_1_LC_7_4_4 .LUT_INIT=16'b0110000011001100;
    LogicCell40 \uart.bit_Count_1_LC_7_4_4  (
            .in0(N__2602),
            .in1(N__2649),
            .in2(N__2420),
            .in3(N__2722),
            .lcout(\uart.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4875),
            .ce(),
            .sr(N__5550));
    defparam \uart.bit_Count_2_LC_7_4_7 .C_ON=1'b0;
    defparam \uart.bit_Count_2_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \uart.bit_Count_2_LC_7_4_7 .LUT_INIT=16'b0111100001010000;
    LogicCell40 \uart.bit_Count_2_LC_7_4_7  (
            .in0(N__2723),
            .in1(N__2402),
            .in2(N__2711),
            .in3(N__2417),
            .lcout(\uart.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4875),
            .ce(),
            .sr(N__5550));
    defparam \uart.data_Aux_RNO_0_6_LC_7_5_0 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_6_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_6_LC_7_5_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart.data_Aux_RNO_0_6_LC_7_5_0  (
            .in0(N__2651),
            .in1(N__2709),
            .in2(_gnd_net_),
            .in3(N__2604),
            .lcout(),
            .ltout(\uart.data_Auxce_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_6_LC_7_5_1 .C_ON=1'b0;
    defparam \uart.data_Aux_6_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_6_LC_7_5_1 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \uart.data_Aux_6_LC_7_5_1  (
            .in0(N__4570),
            .in1(N__2782),
            .in2(N__2405),
            .in3(N__3672),
            .lcout(\uart.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4871),
            .ce(),
            .sr(N__3454));
    defparam \uart.bit_Count_RNO_0_2_LC_7_5_3 .C_ON=1'b0;
    defparam \uart.bit_Count_RNO_0_2_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNO_0_2_LC_7_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart.bit_Count_RNO_0_2_LC_7_5_3  (
            .in0(N__2603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2650),
            .lcout(\uart.CO1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_8_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__2892),
            .in2(N__3172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_8_1_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2822),
            .in3(N__2447),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_8_1_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_8_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__2990),
            .in2(_gnd_net_),
            .in3(N__2444),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_8_1_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_8_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__3034),
            .in2(_gnd_net_),
            .in3(N__2441),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_8_1_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_8_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__2921),
            .in2(_gnd_net_),
            .in3(N__2438),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_8_1_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_8_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__3002),
            .in2(_gnd_net_),
            .in3(N__2435),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_8_1_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_8_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__2948),
            .in2(_gnd_net_),
            .in3(N__2432),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_8_1_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_8_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(N__2960),
            .in2(_gnd_net_),
            .in3(N__2429),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__4882),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_8_2_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_8_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__2935),
            .in2(_gnd_net_),
            .in3(N__2426),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_8_2_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_8_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__2795),
            .in2(_gnd_net_),
            .in3(N__2423),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_8_2_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_8_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__2807),
            .in2(_gnd_net_),
            .in3(N__2507),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_8_2_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_8_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__3184),
            .in2(_gnd_net_),
            .in3(N__2504),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_8_2_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_8_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__2500),
            .in2(_gnd_net_),
            .in3(N__2489),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_8_2_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_8_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__3218),
            .in2(_gnd_net_),
            .in3(N__2486),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_8_2_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_8_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__2482),
            .in2(_gnd_net_),
            .in3(N__2471),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_8_2_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_8_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__3046),
            .in2(_gnd_net_),
            .in3(N__2468),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__4879),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_8_3_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_8_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__3206),
            .in2(_gnd_net_),
            .in3(N__2465),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__4876),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_8_3_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_8_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__3019),
            .in2(_gnd_net_),
            .in3(N__2462),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__4876),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_8_3_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_8_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_19_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__2459),
            .in2(_gnd_net_),
            .in3(N__2552),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__4876),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_8_3_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_8_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__2549),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__4876),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_8_3_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_8_3_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \reset_module_System.count_21_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__2542),
            .in2(_gnd_net_),
            .in3(N__2546),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4876),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.bit_Count_RNIETHE_2_LC_8_3_5 .C_ON=1'b0;
    defparam \uart.bit_Count_RNIETHE_2_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \uart.bit_Count_RNIETHE_2_LC_8_3_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart.bit_Count_RNIETHE_2_LC_8_3_5  (
            .in0(N__2696),
            .in1(N__2644),
            .in2(_gnd_net_),
            .in3(N__2598),
            .lcout(\uart.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_5_LC_8_3_6 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_5_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_5_LC_8_3_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart.data_Aux_RNO_0_5_LC_8_3_6  (
            .in0(N__2599),
            .in1(_gnd_net_),
            .in2(N__2661),
            .in3(N__2697),
            .lcout(\uart.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNI9M0N_1_LC_8_3_7 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI9M0N_1_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI9M0N_1_LC_8_3_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \uart.timer_Count_RNI9M0N_1_LC_8_3_7  (
            .in0(N__3334),
            .in1(N__3505),
            .in2(_gnd_net_),
            .in3(N__4156),
            .lcout(\uart.timer_Count_RNI9M0NZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNILKMA1_0_LC_8_4_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNILKMA1_0_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNILKMA1_0_LC_8_4_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uart.timer_Count_RNILKMA1_0_LC_8_4_1  (
            .in0(N__3929),
            .in1(N__3971),
            .in2(N__4328),
            .in3(N__3890),
            .lcout(),
            .ltout(\uart.timer_Count_RNILKMA1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNILC8T2_3_LC_8_4_2 .C_ON=1'b0;
    defparam \uart.state_RNILC8T2_3_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNILC8T2_3_LC_8_4_2 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \uart.state_RNILC8T2_3_LC_8_4_2  (
            .in0(N__2522),
            .in1(N__3361),
            .in2(N__2513),
            .in3(N__4003),
            .lcout(\uart.un1_state_2_0 ),
            .ltout(\uart.un1_state_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_0_LC_8_4_3 .C_ON=1'b0;
    defparam \uart.data_Aux_0_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_0_LC_8_4_3 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \uart.data_Aux_0_LC_8_4_3  (
            .in0(N__3109),
            .in1(N__2744),
            .in2(N__2510),
            .in3(N__3670),
            .lcout(\uart.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4872),
            .ce(),
            .sr(N__3453));
    defparam \uart.data_Aux_1_LC_8_4_4 .C_ON=1'b0;
    defparam \uart.data_Aux_1_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_1_LC_8_4_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart.data_Aux_1_LC_8_4_4  (
            .in0(N__3668),
            .in1(N__2738),
            .in2(N__4240),
            .in3(N__2774),
            .lcout(\uart.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4872),
            .ce(),
            .sr(N__3453));
    defparam \uart.data_Aux_3_LC_8_4_6 .C_ON=1'b0;
    defparam \uart.data_Aux_3_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_3_LC_8_4_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \uart.data_Aux_3_LC_8_4_6  (
            .in0(N__3669),
            .in1(N__3080),
            .in2(N__2561),
            .in3(N__2775),
            .lcout(\uart.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4872),
            .ce(),
            .sr(N__3453));
    defparam \uart.data_Aux_4_LC_8_4_7 .C_ON=1'b0;
    defparam \uart.data_Aux_4_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_Aux_4_LC_8_4_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart.data_Aux_4_LC_8_4_7  (
            .in0(N__2776),
            .in1(N__2750),
            .in2(N__4600),
            .in3(N__3671),
            .lcout(\uart.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4872),
            .ce(),
            .sr(N__3453));
    defparam \uart.data_Aux_RNO_0_4_LC_8_5_1 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_4_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_4_LC_8_5_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart.data_Aux_RNO_0_4_LC_8_5_1  (
            .in0(N__2609),
            .in1(_gnd_net_),
            .in2(N__2663),
            .in3(N__2708),
            .lcout(\uart.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_0_LC_8_5_2 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_0_LC_8_5_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart.data_Aux_RNO_0_0_LC_8_5_2  (
            .in0(N__2704),
            .in1(N__2652),
            .in2(_gnd_net_),
            .in3(N__2605),
            .lcout(\uart.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_1_LC_8_5_3 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_1_LC_8_5_3 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart.data_Aux_RNO_0_1_LC_8_5_3  (
            .in0(N__2606),
            .in1(_gnd_net_),
            .in2(N__2662),
            .in3(N__2705),
            .lcout(\uart.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_2_LC_8_5_4 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_2_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_2_LC_8_5_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart.data_Aux_RNO_0_2_LC_8_5_4  (
            .in0(N__2706),
            .in1(N__2656),
            .in2(_gnd_net_),
            .in3(N__2607),
            .lcout(\uart.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIA73N2_4_LC_8_5_5 .C_ON=1'b0;
    defparam \uart.state_RNIA73N2_4_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIA73N2_4_LC_8_5_5 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \uart.state_RNIA73N2_4_LC_8_5_5  (
            .in0(N__3362),
            .in1(N__3511),
            .in2(_gnd_net_),
            .in3(N__3565),
            .lcout(\uart.un1_state_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_Aux_RNO_0_3_LC_8_5_6 .C_ON=1'b0;
    defparam \uart.data_Aux_RNO_0_3_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \uart.data_Aux_RNO_0_3_LC_8_5_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart.data_Aux_RNO_0_3_LC_8_5_6  (
            .in0(N__2707),
            .in1(N__2657),
            .in2(_gnd_net_),
            .in3(N__2608),
            .lcout(\uart.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_9_1_0 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_9_1_0 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \reset_module_System.count_0_LC_9_1_0  (
            .in0(N__3171),
            .in1(N__2841),
            .in2(N__2876),
            .in3(N__3133),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4880),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI10J41_1_LC_9_1_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI10J41_1_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI10J41_1_LC_9_1_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \reset_module_System.count_RNI10J41_1_LC_9_1_1  (
            .in0(N__3050),
            .in1(N__3035),
            .in2(N__3023),
            .in3(N__2893),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(\reset_module_System.reset6_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_LC_9_1_2 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_9_1_2 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \reset_module_System.reset_LC_9_1_2  (
            .in0(N__2867),
            .in1(_gnd_net_),
            .in2(N__3005),
            .in3(N__3131),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4880),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_9_1_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_9_1_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_9_1_3  (
            .in0(N__3001),
            .in1(N__2989),
            .in2(N__2978),
            .in3(N__2818),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.reset_iso_LC_9_1_4 .C_ON=1'b0;
    defparam \reset_module_System.reset_iso_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_iso_LC_9_1_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_iso_LC_9_1_4  (
            .in0(N__2868),
            .in1(N__2840),
            .in2(_gnd_net_),
            .in3(N__3132),
            .lcout(reset_module_System_reset_iso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4880),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_9_1_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_9_1_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_9_1_5  (
            .in0(N__2959),
            .in1(N__2947),
            .in2(N__2936),
            .in3(N__2920),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_9_1_6 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_9_1_6 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \reset_module_System.count_1_LC_9_1_6  (
            .in0(N__2909),
            .in1(N__2842),
            .in2(N__2875),
            .in3(N__3134),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4880),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_9_1_7 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_9_1_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \reset_module_System.count_2_LC_9_1_7  (
            .in0(N__3130),
            .in1(N__2866),
            .in2(N__2846),
            .in3(N__2828),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4880),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIP8RT_10_LC_9_2_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIP8RT_10_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIP8RT_10_LC_9_2_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \reset_module_System.count_RNIP8RT_10_LC_9_2_2  (
            .in0(N__2806),
            .in1(N__2794),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\reset_module_System.reset6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI53692_14_LC_9_2_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI53692_14_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI53692_14_LC_9_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI53692_14_LC_9_2_3  (
            .in0(N__3217),
            .in1(N__3205),
            .in2(N__3194),
            .in3(N__3191),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIN3HK3_12_LC_9_2_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIN3HK3_12_LC_9_2_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIN3HK3_12_LC_9_2_4  (
            .in0(N__3185),
            .in1(N__3170),
            .in2(N__3143),
            .in3(N__3140),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_1_3_LC_9_2_5 .C_ON=1'b0;
    defparam \uart.state_RNO_1_3_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_3_LC_9_2_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart.state_RNO_1_3_LC_9_2_5  (
            .in0(N__3352),
            .in1(N__3787),
            .in2(N__3404),
            .in3(N__3818),
            .lcout(),
            .ltout(\uart.N_169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_3_LC_9_2_6 .C_ON=1'b0;
    defparam \uart.state_RNO_0_3_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_3_LC_9_2_6 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart.state_RNO_0_3_LC_9_2_6  (
            .in0(N__3848),
            .in1(N__3305),
            .in2(N__3116),
            .in3(N__5359),
            .lcout(),
            .ltout(\uart.state_srsts_i_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_3_LC_9_2_7 .C_ON=1'b0;
    defparam \uart.state_3_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \uart.state_3_LC_9_2_7 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \uart.state_3_LC_9_2_7  (
            .in0(N__3239),
            .in1(N__3403),
            .in2(N__3113),
            .in3(N__3572),
            .lcout(\uart.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4877),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_esr_0_LC_9_3_0 .C_ON=1'b0;
    defparam \uart.data_esr_0_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_0_LC_9_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_0_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3110),
            .lcout(uart_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4873),
            .ce(N__4547),
            .sr(N__4529));
    defparam \uart.data_esr_2_LC_9_3_2 .C_ON=1'b0;
    defparam \uart.data_esr_2_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_2_LC_9_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_2_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3098),
            .lcout(uart_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4873),
            .ce(N__4547),
            .sr(N__4529));
    defparam \uart.data_esr_3_LC_9_3_3 .C_ON=1'b0;
    defparam \uart.data_esr_3_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_3_LC_9_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_3_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3079),
            .lcout(uart_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4873),
            .ce(N__4547),
            .sr(N__4529));
    defparam \uart.data_esr_5_LC_9_3_5 .C_ON=1'b0;
    defparam \uart.data_esr_5_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_5_LC_9_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_5_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3065),
            .lcout(uart_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4873),
            .ce(N__4547),
            .sr(N__4529));
    defparam \uart.data_esr_7_LC_9_3_7 .C_ON=1'b0;
    defparam \uart.data_esr_7_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_7_LC_9_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_7_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3260),
            .lcout(uart_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4873),
            .ce(N__4547),
            .sr(N__4529));
    defparam \uart.timer_Count_RNI22NA1_6_LC_9_4_0 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI22NA1_6_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI22NA1_6_LC_9_4_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \uart.timer_Count_RNI22NA1_6_LC_9_4_0  (
            .in0(N__3880),
            .in1(N__3813),
            .in2(N__3780),
            .in3(N__3842),
            .lcout(),
            .ltout(\uart.timer_Count10lto5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIT4OA2_2_LC_9_4_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIT4OA2_2_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIT4OA2_2_LC_9_4_1 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \uart.timer_Count_RNIT4OA2_2_LC_9_4_1  (
            .in0(N__3843),
            .in1(N__3920),
            .in2(N__3242),
            .in3(N__3967),
            .lcout(\uart.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_4_2 .C_ON=1'b0;
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNI1HBL_6_LC_9_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.timer_Count_RNI1HBL_6_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__3841),
            .in2(_gnd_net_),
            .in3(N__3812),
            .lcout(\uart.N_145_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_1_LC_9_4_3 .C_ON=1'b0;
    defparam \uart.state_1_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \uart.state_1_LC_9_4_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart.state_1_LC_9_4_3  (
            .in0(N__5362),
            .in1(N__3422),
            .in2(N__3683),
            .in3(N__3287),
            .lcout(\uart.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4868),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIMO1Q_4_LC_9_4_4 .C_ON=1'b0;
    defparam \uart.state_RNIMO1Q_4_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIMO1Q_4_LC_9_4_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart.state_RNIMO1Q_4_LC_9_4_4  (
            .in0(N__3770),
            .in1(N__3500),
            .in2(_gnd_net_),
            .in3(N__5360),
            .lcout(\uart.state_srsts_0_a3_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_4_LC_9_4_5 .C_ON=1'b0;
    defparam \uart.state_RNO_0_4_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_4_LC_9_4_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uart.state_RNO_0_4_LC_9_4_5  (
            .in0(N__5361),
            .in1(N__3237),
            .in2(N__3370),
            .in3(N__3566),
            .lcout(),
            .ltout(\uart.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_4_LC_9_4_6 .C_ON=1'b0;
    defparam \uart.state_4_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \uart.state_4_LC_9_4_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart.state_4_LC_9_4_6  (
            .in0(N__3587),
            .in1(_gnd_net_),
            .in2(N__3221),
            .in3(_gnd_net_),
            .lcout(\uart.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4868),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIB0BC_2_LC_9_4_7 .C_ON=1'b0;
    defparam \uart.state_RNIB0BC_2_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIB0BC_2_LC_9_4_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart.state_RNIB0BC_2_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(N__3392),
            .in2(_gnd_net_),
            .in3(N__3356),
            .lcout(\uart.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIAFHL_4_LC_9_5_3 .C_ON=1'b0;
    defparam \uart.state_RNIAFHL_4_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIAFHL_4_LC_9_5_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart.state_RNIAFHL_4_LC_9_5_3  (
            .in0(N__3360),
            .in1(N__3512),
            .in2(_gnd_net_),
            .in3(N__5376),
            .lcout(\uart.state_RNIAFHLZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_2_LC_9_5_4 .C_ON=1'b0;
    defparam \uart.state_RNO_0_2_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_2_LC_9_5_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \uart.state_RNO_0_2_LC_9_5_4  (
            .in0(N__3420),
            .in1(N__3396),
            .in2(_gnd_net_),
            .in3(N__3676),
            .lcout(),
            .ltout(\uart.N_151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_2_LC_9_5_5 .C_ON=1'b0;
    defparam \uart.state_2_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \uart.state_2_LC_9_5_5 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \uart.state_2_LC_9_5_5  (
            .in0(N__5378),
            .in1(N__3421),
            .in2(N__3407),
            .in3(N__3571),
            .lcout(\uart.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4866),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_2_3_LC_9_5_7 .C_ON=1'b0;
    defparam \uart.state_RNO_2_3_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_2_3_LC_9_5_7 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uart.state_RNO_2_3_LC_9_5_7  (
            .in0(N__3924),
            .in1(N__3964),
            .in2(N__3369),
            .in3(N__3884),
            .lcout(\uart.state_srsts_i_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_1_0_LC_10_1_0 .C_ON=1'b0;
    defparam \uart.state_RNO_1_0_LC_10_1_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_1_0_LC_10_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart.state_RNO_1_0_LC_10_1_0  (
            .in0(_gnd_net_),
            .in1(N__3788),
            .in2(_gnd_net_),
            .in3(N__3520),
            .lcout(),
            .ltout(\uart.N_166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNO_0_0_LC_10_1_1 .C_ON=1'b0;
    defparam \uart.state_RNO_0_0_LC_10_1_1 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNO_0_0_LC_10_1_1 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \uart.state_RNO_0_0_LC_10_1_1  (
            .in0(N__3283),
            .in1(N__3681),
            .in2(N__3293),
            .in3(N__5358),
            .lcout(),
            .ltout(\uart.state_srsts_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_0_LC_10_1_2 .C_ON=1'b0;
    defparam \uart.state_0_LC_10_1_2 .SEQ_MODE=4'b1000;
    defparam \uart.state_0_LC_10_1_2 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \uart.state_0_LC_10_1_2  (
            .in0(N__3521),
            .in1(N__3539),
            .in2(N__3290),
            .in3(N__4007),
            .lcout(\uart.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4874),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_1_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_1_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_1_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_2_LC_10_1_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_2_LC_10_1_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_2_LC_10_1_4 .LUT_INIT=16'b0000000010100110;
    LogicCell40 \uart_frame_decoder.count_2_LC_10_1_4  (
            .in0(N__4061),
            .in1(N__4081),
            .in2(N__3272),
            .in3(N__4094),
            .lcout(\uart_frame_decoder.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4874),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_10_1_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_10_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNIV5MS_0_LC_10_1_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uart_frame_decoder.count_RNIV5MS_0_LC_10_1_5  (
            .in0(N__5030),
            .in1(N__5455),
            .in2(_gnd_net_),
            .in3(N__4037),
            .lcout(\uart_frame_decoder.N_43 ),
            .ltout(\uart_frame_decoder.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_1_LC_10_1_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_1_LC_10_1_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_1_LC_10_1_6 .LUT_INIT=16'b0000000011000011;
    LogicCell40 \uart_frame_decoder.count_1_LC_10_1_6  (
            .in0(_gnd_net_),
            .in1(N__4080),
            .in2(N__3467),
            .in3(N__4093),
            .lcout(\uart_frame_decoder.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4874),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIMBMF_1_LC_10_2_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIMBMF_1_LC_10_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIMBMF_1_LC_10_2_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_RNIMBMF_1_LC_10_2_4  (
            .in0(_gnd_net_),
            .in1(N__5026),
            .in2(_gnd_net_),
            .in3(N__5215),
            .lcout(\uart_frame_decoder.state_1_ns_i_i_a2_1_1_0 ),
            .ltout(\uart_frame_decoder.state_1_ns_i_i_a2_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_10_2_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_10_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_1_0_LC_10_2_5 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_1_0_LC_10_2_5  (
            .in0(N__3692),
            .in1(N__4269),
            .in2(N__3464),
            .in3(N__4255),
            .lcout(),
            .ltout(\uart_frame_decoder.N_81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_0_LC_10_2_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_0_LC_10_2_6 .SEQ_MODE=4'b1001;
    defparam \uart_frame_decoder.state_1_0_LC_10_2_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_frame_decoder.state_1_0_LC_10_2_6  (
            .in0(N__4166),
            .in1(N__4927),
            .in2(N__3461),
            .in3(N__4334),
            .lcout(\uart_frame_decoder.state_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4869),
            .ce(),
            .sr(N__5536));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_10_3_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_10_3_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_0_1_2_LC_10_3_0  (
            .in0(_gnd_net_),
            .in1(N__3721),
            .in2(_gnd_net_),
            .in3(N__3700),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_10_3_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI5BVV_1_LC_10_3_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_frame_decoder.state_1_RNI5BVV_1_LC_10_3_1  (
            .in0(N__5207),
            .in1(N__3709),
            .in2(N__3458),
            .in3(N__3730),
            .lcout(\uart_frame_decoder.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_10_3_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_3_0_LC_10_3_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_frame_decoder.state_1_RNO_3_0_LC_10_3_2  (
            .in0(N__4182),
            .in1(N__5206),
            .in2(_gnd_net_),
            .in3(N__5422),
            .lcout(\uart_frame_decoder.state_1_ns_i_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.data_rdy_LC_10_3_3 .C_ON=1'b0;
    defparam \uart.data_rdy_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_rdy_LC_10_3_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart.data_rdy_LC_10_3_3  (
            .in0(N__3980),
            .in1(N__3677),
            .in2(_gnd_net_),
            .in3(N__5368),
            .lcout(uart_data_rdy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4867),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_0_2_LC_10_3_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_0_2_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_0_2_LC_10_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_0_2_LC_10_3_4  (
            .in0(_gnd_net_),
            .in1(N__5423),
            .in2(_gnd_net_),
            .in3(N__4583),
            .lcout(),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_1_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_10_3_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_10_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_1_2_LC_10_3_5  (
            .in0(N__4559),
            .in1(N__3740),
            .in2(N__3734),
            .in3(N__4223),
            .lcout(\uart_frame_decoder.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_10_3_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_10_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_frame_decoder.state_1_ns_0_i_a2_0_4_1_LC_10_3_6  (
            .in0(N__3731),
            .in1(N__3722),
            .in2(N__3713),
            .in3(N__3701),
            .lcout(\uart_frame_decoder.N_79_4 ),
            .ltout(\uart_frame_decoder.N_79_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_10_3_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_1_LC_10_3_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_1_LC_10_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3686),
            .in3(N__4183),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNI78E91_4_LC_10_4_0 .C_ON=1'b0;
    defparam \uart.state_RNI78E91_4_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNI78E91_4_LC_10_4_0 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \uart.state_RNI78E91_4_LC_10_4_0  (
            .in0(N__3501),
            .in1(N__3771),
            .in2(N__3682),
            .in3(N__4000),
            .lcout(),
            .ltout(\uart.data_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIS4183_7_LC_10_4_1 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIS4183_7_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIS4183_7_LC_10_4_1 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \uart.timer_Count_RNIS4183_7_LC_10_4_1  (
            .in0(N__3772),
            .in1(N__5363),
            .in2(N__3599),
            .in3(N__3534),
            .lcout(\uart.timer_Count_RNIS4183Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_RNIMLMA1_1_LC_10_4_3 .C_ON=1'b0;
    defparam \uart.timer_Count_RNIMLMA1_1_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \uart.timer_Count_RNIMLMA1_1_LC_10_4_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uart.timer_Count_RNIMLMA1_1_LC_10_4_3  (
            .in0(N__4148),
            .in1(N__3966),
            .in2(N__3886),
            .in3(N__3919),
            .lcout(\uart.N_152_0 ),
            .ltout(\uart.N_152_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIDV3Q2_4_LC_10_4_4 .C_ON=1'b0;
    defparam \uart.state_RNIDV3Q2_4_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIDV3Q2_4_LC_10_4_4 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \uart.state_RNIDV3Q2_4_LC_10_4_4  (
            .in0(_gnd_net_),
            .in1(N__3596),
            .in2(N__3590),
            .in3(N__4001),
            .lcout(\uart.N_167 ),
            .ltout(\uart.N_167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIIHDQ5_2_LC_10_4_5 .C_ON=1'b0;
    defparam \uart.state_RNIIHDQ5_2_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIIHDQ5_2_LC_10_4_5 .LUT_INIT=16'b1100111111001110;
    LogicCell40 \uart.state_RNIIHDQ5_2_LC_10_4_5  (
            .in0(N__3581),
            .in1(N__5364),
            .in2(N__3575),
            .in3(N__3567),
            .lcout(\uart.timer_Count_1_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNIGITG2_4_LC_10_4_6 .C_ON=1'b0;
    defparam \uart.state_RNIGITG2_4_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNIGITG2_4_LC_10_4_6 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \uart.state_RNIGITG2_4_LC_10_4_6  (
            .in0(N__3535),
            .in1(N__3773),
            .in2(N__3513),
            .in3(N__4002),
            .lcout(\uart.state_1_sqmuxa ),
            .ltout(\uart.state_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.state_RNICNUO5_4_LC_10_4_7 .C_ON=1'b0;
    defparam \uart.state_RNICNUO5_4_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \uart.state_RNICNUO5_4_LC_10_4_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart.state_RNICNUO5_4_LC_10_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3974),
            .in3(N__4515),
            .lcout(\uart.state_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_10_5_0 .C_ON=1'b1;
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \uart.un4_timer_Count_1_cry_1_c_LC_10_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart.un4_timer_Count_1_cry_1_c_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__4324),
            .in2(N__4160),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\uart.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_2_LC_10_5_1 .C_ON=1'b1;
    defparam \uart.timer_Count_2_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_2_LC_10_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_2_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__3965),
            .in2(_gnd_net_),
            .in3(N__3932),
            .lcout(\uart.timer_CountZ0Z_2 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_1 ),
            .carryout(\uart.un4_timer_Count_1_cry_2 ),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart.timer_Count_3_LC_10_5_2 .C_ON=1'b1;
    defparam \uart.timer_Count_3_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_3_LC_10_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_3_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__3925),
            .in2(_gnd_net_),
            .in3(N__3893),
            .lcout(\uart.timer_CountZ0Z_3 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_2 ),
            .carryout(\uart.un4_timer_Count_1_cry_3 ),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart.timer_Count_4_LC_10_5_3 .C_ON=1'b1;
    defparam \uart.timer_Count_4_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_4_LC_10_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_4_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__3885),
            .in2(_gnd_net_),
            .in3(N__3851),
            .lcout(\uart.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_3 ),
            .carryout(\uart.un4_timer_Count_1_cry_4 ),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart.timer_Count_5_LC_10_5_4 .C_ON=1'b1;
    defparam \uart.timer_Count_5_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_5_LC_10_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_5_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__3847),
            .in2(_gnd_net_),
            .in3(N__3821),
            .lcout(\uart.timer_CountZ0Z_5 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_4 ),
            .carryout(\uart.un4_timer_Count_1_cry_5 ),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart.timer_Count_6_LC_10_5_5 .C_ON=1'b1;
    defparam \uart.timer_Count_6_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_6_LC_10_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart.timer_Count_6_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__3817),
            .in2(_gnd_net_),
            .in3(N__3794),
            .lcout(\uart.timer_CountZ0Z_6 ),
            .ltout(),
            .carryin(\uart.un4_timer_Count_1_cry_5 ),
            .carryout(\uart.un4_timer_Count_1_cry_6 ),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart.timer_Count_7_LC_10_5_6 .C_ON=1'b0;
    defparam \uart.timer_Count_7_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_7_LC_10_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart.timer_Count_7_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(N__3779),
            .in2(_gnd_net_),
            .in3(N__3791),
            .lcout(\uart.timer_CountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4862),
            .ce(),
            .sr(N__4294));
    defparam \uart_frame_decoder.count8_cry_0_c_LC_11_1_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_LC_11_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_LC_11_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(\uart_frame_decoder.count8_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_11_1_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_1_c_inv_LC_11_1_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_1_c_inv_LC_11_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4127),
            .in3(N__4076),
            .lcout(\uart_frame_decoder.count8_axb_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_0 ),
            .carryout(\uart_frame_decoder.count8_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_11_1_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_inv_LC_11_1_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_inv_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(N__4046),
            .in2(N__4118),
            .in3(N__4059),
            .lcout(\uart_frame_decoder.count_i_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.count8_cry_1 ),
            .carryout(\uart_frame_decoder.count8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_11_1_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_THRU_LUT4_0_LC_11_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_frame_decoder.count8_THRU_LUT4_0_LC_11_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4109),
            .lcout(\uart_frame_decoder.count8_THRU_CO ),
            .ltout(\uart_frame_decoder.count8_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_11_1_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_11_1_4 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \uart_frame_decoder.count8_cry_2_c_RNICKS21_LC_11_1_4  (
            .in0(N__5031),
            .in1(N__5458),
            .in2(N__4097),
            .in3(N__5372),
            .lcout(\uart_frame_decoder.N_37 ),
            .ltout(\uart_frame_decoder.N_37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_0_LC_11_1_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_0_LC_11_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.count_0_LC_11_1_5 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uart_frame_decoder.count_0_LC_11_1_5  (
            .in0(N__5459),
            .in1(N__5032),
            .in2(N__4085),
            .in3(N__4036),
            .lcout(\uart_frame_decoder.count8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4870),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count_RNIHPR51_2_LC_11_1_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.count_RNIHPR51_2_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count_RNIHPR51_2_LC_11_1_6 .LUT_INIT=16'b0000010111111111;
    LogicCell40 \uart_frame_decoder.count_RNIHPR51_2_LC_11_1_6  (
            .in0(N__4035),
            .in1(_gnd_net_),
            .in2(N__4082),
            .in3(N__4060),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_o2_0_tz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_11_1_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.count8_cry_0_c_inv_LC_11_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_frame_decoder.count8_cry_0_c_inv_LC_11_1_7  (
            .in0(N__4045),
            .in1(N__4018),
            .in2(_gnd_net_),
            .in3(N__4034),
            .lcout(\uart_frame_decoder.count8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIOAVK1_5_LC_11_2_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIOAVK1_5_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIOAVK1_5_LC_11_2_0 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \uart_frame_decoder.WDT_RNIOAVK1_5_LC_11_2_0  (
            .in0(N__4800),
            .in1(N__4727),
            .in2(N__4430),
            .in3(N__4205),
            .lcout(),
            .ltout(\uart_frame_decoder.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIGSL62_15_LC_11_2_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIGSL62_15_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIGSL62_15_LC_11_2_1 .LUT_INIT=16'b1111011101010101;
    LogicCell40 \uart_frame_decoder.WDT_RNIGSL62_15_LC_11_2_1  (
            .in0(N__4953),
            .in1(N__4661),
            .in2(N__4214),
            .in3(N__4211),
            .lcout(\uart_frame_decoder.WDT8_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIEKPB_11_LC_11_2_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIEKPB_11_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIEKPB_11_LC_11_2_2 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \uart_frame_decoder.WDT_RNIEKPB_11_LC_11_2_2  (
            .in0(N__4704),
            .in1(N__4683),
            .in2(N__4664),
            .in3(N__4639),
            .lcout(\uart_frame_decoder.g0_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIRBB11_4_LC_11_2_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIRBB11_4_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIRBB11_4_LC_11_2_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_frame_decoder.WDT_RNIRBB11_4_LC_11_2_3  (
            .in0(N__4780),
            .in1(N__4446),
            .in2(N__4403),
            .in3(N__4752),
            .lcout(\uart_frame_decoder.g0_1_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_11_2_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIQAB11_4_LC_11_2_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_frame_decoder.WDT_RNIQAB11_4_LC_11_2_4  (
            .in0(N__4447),
            .in1(N__4425),
            .in2(N__4781),
            .in3(N__4753),
            .lcout(\uart_frame_decoder.WDT_RNIQAB11Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIVBR8_15_LC_11_2_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIVBR8_15_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIVBR8_15_LC_11_2_5 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \uart_frame_decoder.WDT_RNIVBR8_15_LC_11_2_5  (
            .in0(N__4640),
            .in1(_gnd_net_),
            .in2(N__4955),
            .in3(N__4662),
            .lcout(\uart_frame_decoder.WDT8lto15 ),
            .ltout(\uart_frame_decoder.WDT8lto15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNILEPU1_10_LC_11_2_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNILEPU1_10_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNILEPU1_10_LC_11_2_6 .LUT_INIT=16'b1000110000000100;
    LogicCell40 \uart_frame_decoder.state_1_RNILEPU1_10_LC_11_2_6  (
            .in0(N__5456),
            .in1(N__5017),
            .in2(N__4199),
            .in3(N__4196),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10 ),
            .ltout(\uart_frame_decoder.state_1_ns_0_i_a2_0_0_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_11_2_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_2_0_LC_11_2_7 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \uart_frame_decoder.state_1_RNO_2_0_LC_11_2_7  (
            .in0(N__4190),
            .in1(N__4184),
            .in2(N__4169),
            .in3(N__5457),
            .lcout(\uart_frame_decoder.N_35_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_1_LC_11_3_1 .C_ON=1'b0;
    defparam \uart.timer_Count_1_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_1_LC_11_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart.timer_Count_1_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__4320),
            .in2(_gnd_net_),
            .in3(N__4155),
            .lcout(\uart.timer_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4865),
            .ce(),
            .sr(N__4295));
    defparam \uart_frame_decoder.WDT_RNISS5H_11_LC_11_3_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNISS5H_11_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNISS5H_11_LC_11_3_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \uart_frame_decoder.WDT_RNISS5H_11_LC_11_3_2  (
            .in0(N__4684),
            .in1(N__4705),
            .in2(N__4733),
            .in3(N__4401),
            .lcout(),
            .ltout(\uart_frame_decoder.WDT_RNISS5HZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIEDQT1_7_LC_11_3_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIEDQT1_7_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIEDQT1_7_LC_11_3_3 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \uart_frame_decoder.WDT_RNIEDQT1_7_LC_11_3_3  (
            .in0(N__4379),
            .in1(N__4731),
            .in2(N__4373),
            .in3(N__4801),
            .lcout(\uart_frame_decoder.WDT8lt13 ),
            .ltout(\uart_frame_decoder.WDT8lt13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNIKVEI2_14_LC_11_3_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNIKVEI2_14_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNIKVEI2_14_LC_11_3_4 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \uart_frame_decoder.WDT_RNIKVEI2_14_LC_11_3_4  (
            .in0(N__5443),
            .in1(N__4345),
            .in2(N__4370),
            .in3(N__4631),
            .lcout(\uart_frame_decoder.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.WDT_RNI85RG2_14_LC_11_3_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_RNI85RG2_14_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.WDT_RNI85RG2_14_LC_11_3_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uart_frame_decoder.WDT_RNI85RG2_14_LC_11_3_5  (
            .in0(N__4630),
            .in1(N__5008),
            .in2(N__4361),
            .in3(N__5444),
            .lcout(\uart_frame_decoder.state_1_ns_0_i_a2_0_d_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_11_3_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNO_0_0_LC_11_3_6 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \uart_frame_decoder.state_1_RNO_0_0_LC_11_3_6  (
            .in0(N__4367),
            .in1(N__4357),
            .in2(N__4349),
            .in3(N__4632),
            .lcout(\uart_frame_decoder.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart.timer_Count_0_LC_11_3_7 .C_ON=1'b0;
    defparam \uart.timer_Count_0_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \uart.timer_Count_0_LC_11_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart.timer_Count_0_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4319),
            .lcout(\uart.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4865),
            .ce(),
            .sr(N__4295));
    defparam \uart_frame_decoder.state_1_1_LC_11_4_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_1_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_1_LC_11_4_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uart_frame_decoder.state_1_1_LC_11_4_1  (
            .in0(N__5211),
            .in1(N__4270),
            .in2(N__4283),
            .in3(N__4908),
            .lcout(\uart_frame_decoder.state_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4863),
            .ce(),
            .sr(N__5549));
    defparam \uart_frame_decoder.state_1_2_LC_11_4_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_2_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_2_LC_11_4_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_2_LC_11_4_2  (
            .in0(N__4909),
            .in1(N__5074),
            .in2(N__4274),
            .in3(N__4256),
            .lcout(\uart_frame_decoder.state_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4863),
            .ce(),
            .sr(N__5549));
    defparam \uart.data_esr_1_LC_11_5_2 .C_ON=1'b0;
    defparam \uart.data_esr_1_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_1_LC_11_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart.data_esr_1_LC_11_5_2  (
            .in0(N__4244),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uart_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4860),
            .ce(N__4546),
            .sr(N__4528));
    defparam \uart.data_esr_4_LC_11_5_3 .C_ON=1'b0;
    defparam \uart.data_esr_4_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_4_LC_11_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_4_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4604),
            .lcout(uart_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4860),
            .ce(N__4546),
            .sr(N__4528));
    defparam \uart.data_esr_6_LC_11_5_7 .C_ON=1'b0;
    defparam \uart.data_esr_6_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \uart.data_esr_6_LC_11_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart.data_esr_6_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4574),
            .lcout(uart_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4860),
            .ce(N__4546),
            .sr(N__4528));
    defparam \uart_frame_decoder.WDT_0_LC_12_2_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_0_LC_12_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_0_LC_12_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_0_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__4481),
            .in2(N__4498),
            .in3(N__4499),
            .lcout(\uart_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_1_LC_12_2_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_1_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_1_LC_12_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_1_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__4475),
            .in2(_gnd_net_),
            .in3(N__4469),
            .lcout(\uart_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_2_LC_12_2_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_2_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_2_LC_12_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_2_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__4466),
            .in2(_gnd_net_),
            .in3(N__4460),
            .lcout(\uart_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_3_LC_12_2_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_3_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_3_LC_12_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_3_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(N__4457),
            .in2(_gnd_net_),
            .in3(N__4451),
            .lcout(\uart_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_4_LC_12_2_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_4_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_4_LC_12_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_4_LC_12_2_4  (
            .in0(_gnd_net_),
            .in1(N__4448),
            .in2(_gnd_net_),
            .in3(N__4433),
            .lcout(\uart_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_5_LC_12_2_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_5_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_5_LC_12_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_5_LC_12_2_5  (
            .in0(_gnd_net_),
            .in1(N__4426),
            .in2(_gnd_net_),
            .in3(N__4406),
            .lcout(\uart_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_6_LC_12_2_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_6_LC_12_2_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_6_LC_12_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_6_LC_12_2_6  (
            .in0(_gnd_net_),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__4382),
            .lcout(\uart_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_7_LC_12_2_7 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_7_LC_12_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_7_LC_12_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_7_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(N__4802),
            .in2(_gnd_net_),
            .in3(N__4784),
            .lcout(\uart_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__4864),
            .ce(),
            .sr(N__5300));
    defparam \uart_frame_decoder.WDT_8_LC_12_3_0 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_8_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_8_LC_12_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_8_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__4779),
            .in2(_gnd_net_),
            .in3(N__4757),
            .lcout(\uart_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\uart_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_9_LC_12_3_1 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_9_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_9_LC_12_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_9_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__4754),
            .in2(_gnd_net_),
            .in3(N__4736),
            .lcout(\uart_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_10_LC_12_3_2 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_10_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_10_LC_12_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_10_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__4732),
            .in2(_gnd_net_),
            .in3(N__4709),
            .lcout(\uart_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_11_LC_12_3_3 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_11_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_11_LC_12_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_11_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__4706),
            .in2(_gnd_net_),
            .in3(N__4688),
            .lcout(\uart_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_12_LC_12_3_4 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_12_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_12_LC_12_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_12_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__4685),
            .in2(_gnd_net_),
            .in3(N__4667),
            .lcout(\uart_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_13_LC_12_3_5 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_13_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_13_LC_12_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_13_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__4663),
            .in2(_gnd_net_),
            .in3(N__4643),
            .lcout(\uart_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_14_LC_12_3_6 .C_ON=1'b1;
    defparam \uart_frame_decoder.WDT_14_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_14_LC_12_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_frame_decoder.WDT_14_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__4633),
            .in2(_gnd_net_),
            .in3(N__4607),
            .lcout(\uart_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\uart_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\uart_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.WDT_15_LC_12_3_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.WDT_15_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.WDT_15_LC_12_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_frame_decoder.WDT_15_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__4954),
            .in2(_gnd_net_),
            .in3(N__4958),
            .lcout(\uart_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4861),
            .ce(),
            .sr(N__5296));
    defparam \uart_frame_decoder.state_1_10_LC_12_4_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_10_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_10_LC_12_4_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \uart_frame_decoder.state_1_10_LC_12_4_0  (
            .in0(N__4937),
            .in1(N__5495),
            .in2(N__5183),
            .in3(N__4928),
            .lcout(\uart_frame_decoder.state_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_3_LC_12_4_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_3_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_3_LC_12_4_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_3_LC_12_4_1  (
            .in0(N__5491),
            .in1(N__5073),
            .in2(N__5057),
            .in3(N__4910),
            .lcout(\uart_frame_decoder.state_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_4_LC_12_4_2 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_4_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_4_LC_12_4_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uart_frame_decoder.state_1_4_LC_12_4_2  (
            .in0(N__4911),
            .in1(N__5496),
            .in2(N__5279),
            .in3(N__5051),
            .lcout(\uart_frame_decoder.state_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_5_LC_12_4_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_5_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_5_LC_12_4_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_5_LC_12_4_3  (
            .in0(N__5492),
            .in1(N__5274),
            .in2(N__5159),
            .in3(N__4912),
            .lcout(\uart_frame_decoder.state_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_6_LC_12_4_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_6_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_6_LC_12_4_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uart_frame_decoder.state_1_6_LC_12_4_4  (
            .in0(N__4913),
            .in1(N__5497),
            .in2(N__5123),
            .in3(N__5153),
            .lcout(\uart_frame_decoder.state_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_7_LC_12_4_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_7_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_7_LC_12_4_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uart_frame_decoder.state_1_7_LC_12_4_5  (
            .in0(N__5493),
            .in1(N__5118),
            .in2(N__5105),
            .in3(N__4914),
            .lcout(\uart_frame_decoder.state_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_8_LC_12_4_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_8_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_8_LC_12_4_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uart_frame_decoder.state_1_8_LC_12_4_6  (
            .in0(N__4915),
            .in1(N__5102),
            .in2(N__5504),
            .in3(N__5244),
            .lcout(\uart_frame_decoder.state_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.state_1_9_LC_12_4_7 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_9_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_frame_decoder.state_1_9_LC_12_4_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uart_frame_decoder.state_1_9_LC_12_4_7  (
            .in0(N__5494),
            .in1(N__5180),
            .in2(N__5246),
            .in3(N__4916),
            .lcout(\uart_frame_decoder.state_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4859),
            .ce(),
            .sr(N__5552));
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_13_3_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_13_3_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_frame_decoder.source_data_valid_2_sqmuxa_i_LC_13_3_6  (
            .in0(_gnd_net_),
            .in1(N__5460),
            .in2(_gnd_net_),
            .in3(N__5377),
            .lcout(\uart_frame_decoder.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIUQR11_4_LC_13_4_0 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIUQR11_4_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIUQR11_4_LC_13_4_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \uart_frame_decoder.state_1_RNIUQR11_4_LC_13_4_0  (
            .in0(N__5278),
            .in1(N__5084),
            .in2(_gnd_net_),
            .in3(N__5158),
            .lcout(uart_frame_decoder_N_307_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI8L5O_8_LC_13_4_1 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI8L5O_8_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI8L5O_8_LC_13_4_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uart_frame_decoder.state_1_RNI8L5O_8_LC_13_4_1  (
            .in0(N__5009),
            .in1(N__5245),
            .in2(_gnd_net_),
            .in3(N__5182),
            .lcout(uart_frame_decoder_N_308_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNICQTG_7_LC_13_4_3 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNICQTG_7_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNICQTG_7_LC_13_4_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_frame_decoder.state_1_RNICQTG_7_LC_13_4_3  (
            .in0(_gnd_net_),
            .in1(N__5103),
            .in2(_gnd_net_),
            .in3(N__5216),
            .lcout(),
            .ltout(\uart_frame_decoder.un14_i_a2_0_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNI3NAA1_3_LC_13_4_4 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNI3NAA1_3_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNI3NAA1_3_LC_13_4_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \uart_frame_decoder.state_1_RNI3NAA1_3_LC_13_4_4  (
            .in0(N__5181),
            .in1(N__5055),
            .in2(N__5162),
            .in3(N__5157),
            .lcout(uart_frame_decoder_N_305_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNIHVTG_6_LC_13_4_5 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNIHVTG_6_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNIHVTG_6_LC_13_4_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart_frame_decoder.state_1_RNIHVTG_6_LC_13_4_5  (
            .in0(N__5122),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5104),
            .lcout(\uart_frame_decoder.N_306_1 ),
            .ltout(\uart_frame_decoder.N_306_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_frame_decoder.state_1_RNID8391_2_LC_13_4_6 .C_ON=1'b0;
    defparam \uart_frame_decoder.state_1_RNID8391_2_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \uart_frame_decoder.state_1_RNID8391_2_LC_13_4_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \uart_frame_decoder.state_1_RNID8391_2_LC_13_4_6  (
            .in0(N__5078),
            .in1(N__5056),
            .in2(N__5036),
            .in3(N__5010),
            .lcout(uart_frame_decoder_N_306_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // Pc2Drone
