// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 16 2019 22:03:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "Pc2drone" view "INTERFACE"

module Pc2drone (
    uart_input_pc,
    debug_CH5_31B,
    debug_CH3_20A,
    debug_CH0_16A,
    uart_input_drone,
    ppm_output,
    debug_CH6_5B,
    debug_CH2_18A,
    debug_CH4_2A,
    debug_CH1_0A,
    clk_system);

    input uart_input_pc;
    output debug_CH5_31B;
    output debug_CH3_20A;
    output debug_CH0_16A;
    input uart_input_drone;
    output ppm_output;
    output debug_CH6_5B;
    output debug_CH2_18A;
    output debug_CH4_2A;
    output debug_CH1_0A;
    input clk_system;

    wire N__52031;
    wire N__52030;
    wire N__52029;
    wire N__52020;
    wire N__52019;
    wire N__52018;
    wire N__52011;
    wire N__52010;
    wire N__52009;
    wire N__52002;
    wire N__52001;
    wire N__52000;
    wire N__51993;
    wire N__51992;
    wire N__51991;
    wire N__51984;
    wire N__51983;
    wire N__51982;
    wire N__51975;
    wire N__51974;
    wire N__51973;
    wire N__51966;
    wire N__51965;
    wire N__51964;
    wire N__51957;
    wire N__51956;
    wire N__51955;
    wire N__51948;
    wire N__51947;
    wire N__51946;
    wire N__51939;
    wire N__51938;
    wire N__51937;
    wire N__51920;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51908;
    wire N__51907;
    wire N__51904;
    wire N__51901;
    wire N__51898;
    wire N__51895;
    wire N__51892;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51872;
    wire N__51869;
    wire N__51866;
    wire N__51863;
    wire N__51860;
    wire N__51857;
    wire N__51856;
    wire N__51855;
    wire N__51852;
    wire N__51849;
    wire N__51846;
    wire N__51841;
    wire N__51836;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51824;
    wire N__51823;
    wire N__51822;
    wire N__51819;
    wire N__51816;
    wire N__51813;
    wire N__51808;
    wire N__51803;
    wire N__51800;
    wire N__51797;
    wire N__51796;
    wire N__51795;
    wire N__51792;
    wire N__51789;
    wire N__51786;
    wire N__51781;
    wire N__51776;
    wire N__51773;
    wire N__51770;
    wire N__51767;
    wire N__51764;
    wire N__51761;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51750;
    wire N__51747;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51731;
    wire N__51728;
    wire N__51725;
    wire N__51722;
    wire N__51719;
    wire N__51716;
    wire N__51713;
    wire N__51712;
    wire N__51711;
    wire N__51708;
    wire N__51703;
    wire N__51700;
    wire N__51699;
    wire N__51696;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51680;
    wire N__51679;
    wire N__51678;
    wire N__51677;
    wire N__51676;
    wire N__51675;
    wire N__51672;
    wire N__51671;
    wire N__51670;
    wire N__51669;
    wire N__51668;
    wire N__51667;
    wire N__51666;
    wire N__51665;
    wire N__51664;
    wire N__51663;
    wire N__51662;
    wire N__51661;
    wire N__51660;
    wire N__51659;
    wire N__51658;
    wire N__51657;
    wire N__51652;
    wire N__51645;
    wire N__51640;
    wire N__51629;
    wire N__51618;
    wire N__51613;
    wire N__51610;
    wire N__51607;
    wire N__51602;
    wire N__51595;
    wire N__51592;
    wire N__51587;
    wire N__51582;
    wire N__51575;
    wire N__51572;
    wire N__51569;
    wire N__51566;
    wire N__51563;
    wire N__51562;
    wire N__51561;
    wire N__51558;
    wire N__51555;
    wire N__51552;
    wire N__51547;
    wire N__51542;
    wire N__51541;
    wire N__51540;
    wire N__51539;
    wire N__51538;
    wire N__51537;
    wire N__51536;
    wire N__51535;
    wire N__51534;
    wire N__51533;
    wire N__51532;
    wire N__51531;
    wire N__51530;
    wire N__51529;
    wire N__51528;
    wire N__51527;
    wire N__51526;
    wire N__51525;
    wire N__51524;
    wire N__51523;
    wire N__51522;
    wire N__51521;
    wire N__51520;
    wire N__51519;
    wire N__51518;
    wire N__51517;
    wire N__51516;
    wire N__51515;
    wire N__51514;
    wire N__51513;
    wire N__51512;
    wire N__51511;
    wire N__51510;
    wire N__51509;
    wire N__51508;
    wire N__51507;
    wire N__51506;
    wire N__51505;
    wire N__51504;
    wire N__51503;
    wire N__51502;
    wire N__51501;
    wire N__51500;
    wire N__51499;
    wire N__51498;
    wire N__51497;
    wire N__51496;
    wire N__51495;
    wire N__51494;
    wire N__51493;
    wire N__51492;
    wire N__51491;
    wire N__51490;
    wire N__51489;
    wire N__51488;
    wire N__51487;
    wire N__51486;
    wire N__51485;
    wire N__51484;
    wire N__51483;
    wire N__51482;
    wire N__51481;
    wire N__51480;
    wire N__51479;
    wire N__51478;
    wire N__51477;
    wire N__51476;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51472;
    wire N__51471;
    wire N__51470;
    wire N__51469;
    wire N__51468;
    wire N__51467;
    wire N__51466;
    wire N__51465;
    wire N__51464;
    wire N__51463;
    wire N__51462;
    wire N__51461;
    wire N__51460;
    wire N__51459;
    wire N__51458;
    wire N__51457;
    wire N__51456;
    wire N__51455;
    wire N__51454;
    wire N__51453;
    wire N__51452;
    wire N__51451;
    wire N__51450;
    wire N__51449;
    wire N__51448;
    wire N__51447;
    wire N__51446;
    wire N__51445;
    wire N__51444;
    wire N__51443;
    wire N__51442;
    wire N__51441;
    wire N__51440;
    wire N__51439;
    wire N__51438;
    wire N__51437;
    wire N__51436;
    wire N__51435;
    wire N__51434;
    wire N__51433;
    wire N__51432;
    wire N__51431;
    wire N__51430;
    wire N__51429;
    wire N__51428;
    wire N__51427;
    wire N__51426;
    wire N__51425;
    wire N__51424;
    wire N__51423;
    wire N__51422;
    wire N__51421;
    wire N__51420;
    wire N__51419;
    wire N__51418;
    wire N__51417;
    wire N__51416;
    wire N__51415;
    wire N__51414;
    wire N__51413;
    wire N__51412;
    wire N__51411;
    wire N__51410;
    wire N__51409;
    wire N__51408;
    wire N__51407;
    wire N__51406;
    wire N__51405;
    wire N__51404;
    wire N__51403;
    wire N__51402;
    wire N__51401;
    wire N__51400;
    wire N__51399;
    wire N__51398;
    wire N__51397;
    wire N__51396;
    wire N__51395;
    wire N__51394;
    wire N__51393;
    wire N__51392;
    wire N__51391;
    wire N__51390;
    wire N__51389;
    wire N__51388;
    wire N__51387;
    wire N__51386;
    wire N__51385;
    wire N__51384;
    wire N__51383;
    wire N__51382;
    wire N__51381;
    wire N__51380;
    wire N__51379;
    wire N__51378;
    wire N__51377;
    wire N__51376;
    wire N__51375;
    wire N__51374;
    wire N__51373;
    wire N__51372;
    wire N__51371;
    wire N__51370;
    wire N__51369;
    wire N__51368;
    wire N__51367;
    wire N__51366;
    wire N__51365;
    wire N__51364;
    wire N__51363;
    wire N__51362;
    wire N__51361;
    wire N__51360;
    wire N__51359;
    wire N__51358;
    wire N__51357;
    wire N__51356;
    wire N__51355;
    wire N__51354;
    wire N__51353;
    wire N__51352;
    wire N__51351;
    wire N__51350;
    wire N__51349;
    wire N__51348;
    wire N__51347;
    wire N__51346;
    wire N__51345;
    wire N__51344;
    wire N__51343;
    wire N__51342;
    wire N__51341;
    wire N__51340;
    wire N__51339;
    wire N__51338;
    wire N__51337;
    wire N__51336;
    wire N__51335;
    wire N__51334;
    wire N__51333;
    wire N__51332;
    wire N__51331;
    wire N__51330;
    wire N__51329;
    wire N__51328;
    wire N__51327;
    wire N__51326;
    wire N__51325;
    wire N__51324;
    wire N__51323;
    wire N__51322;
    wire N__51321;
    wire N__51320;
    wire N__51319;
    wire N__51318;
    wire N__51317;
    wire N__51316;
    wire N__51315;
    wire N__51314;
    wire N__51313;
    wire N__51312;
    wire N__51311;
    wire N__51310;
    wire N__51309;
    wire N__51308;
    wire N__51307;
    wire N__51306;
    wire N__50831;
    wire N__50828;
    wire N__50825;
    wire N__50824;
    wire N__50823;
    wire N__50822;
    wire N__50821;
    wire N__50820;
    wire N__50819;
    wire N__50818;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50814;
    wire N__50813;
    wire N__50812;
    wire N__50811;
    wire N__50810;
    wire N__50809;
    wire N__50808;
    wire N__50807;
    wire N__50806;
    wire N__50805;
    wire N__50804;
    wire N__50803;
    wire N__50802;
    wire N__50801;
    wire N__50800;
    wire N__50799;
    wire N__50798;
    wire N__50797;
    wire N__50796;
    wire N__50795;
    wire N__50788;
    wire N__50781;
    wire N__50776;
    wire N__50773;
    wire N__50762;
    wire N__50755;
    wire N__50746;
    wire N__50741;
    wire N__50738;
    wire N__50735;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50717;
    wire N__50716;
    wire N__50715;
    wire N__50714;
    wire N__50713;
    wire N__50712;
    wire N__50711;
    wire N__50710;
    wire N__50709;
    wire N__50708;
    wire N__50707;
    wire N__50706;
    wire N__50705;
    wire N__50704;
    wire N__50703;
    wire N__50702;
    wire N__50701;
    wire N__50700;
    wire N__50699;
    wire N__50698;
    wire N__50697;
    wire N__50696;
    wire N__50695;
    wire N__50694;
    wire N__50693;
    wire N__50692;
    wire N__50691;
    wire N__50690;
    wire N__50687;
    wire N__50684;
    wire N__50681;
    wire N__50678;
    wire N__50675;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50654;
    wire N__50651;
    wire N__50648;
    wire N__50645;
    wire N__50558;
    wire N__50555;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50540;
    wire N__50539;
    wire N__50536;
    wire N__50533;
    wire N__50530;
    wire N__50527;
    wire N__50524;
    wire N__50523;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50504;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50492;
    wire N__50491;
    wire N__50488;
    wire N__50485;
    wire N__50484;
    wire N__50479;
    wire N__50476;
    wire N__50473;
    wire N__50468;
    wire N__50465;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50453;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50445;
    wire N__50442;
    wire N__50439;
    wire N__50436;
    wire N__50431;
    wire N__50426;
    wire N__50423;
    wire N__50420;
    wire N__50417;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50409;
    wire N__50406;
    wire N__50403;
    wire N__50400;
    wire N__50395;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50381;
    wire N__50378;
    wire N__50377;
    wire N__50374;
    wire N__50373;
    wire N__50370;
    wire N__50367;
    wire N__50364;
    wire N__50361;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50342;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50334;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50318;
    wire N__50315;
    wire N__50312;
    wire N__50311;
    wire N__50308;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50283;
    wire N__50278;
    wire N__50273;
    wire N__50270;
    wire N__50267;
    wire N__50264;
    wire N__50261;
    wire N__50258;
    wire N__50255;
    wire N__50252;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50244;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50228;
    wire N__50227;
    wire N__50226;
    wire N__50223;
    wire N__50222;
    wire N__50219;
    wire N__50218;
    wire N__50217;
    wire N__50216;
    wire N__50215;
    wire N__50214;
    wire N__50213;
    wire N__50212;
    wire N__50209;
    wire N__50208;
    wire N__50207;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50203;
    wire N__50202;
    wire N__50197;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50160;
    wire N__50155;
    wire N__50152;
    wire N__50147;
    wire N__50144;
    wire N__50141;
    wire N__50136;
    wire N__50131;
    wire N__50126;
    wire N__50123;
    wire N__50120;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50108;
    wire N__50107;
    wire N__50104;
    wire N__50101;
    wire N__50096;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50086;
    wire N__50081;
    wire N__50078;
    wire N__50075;
    wire N__50072;
    wire N__50069;
    wire N__50066;
    wire N__50063;
    wire N__50060;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50048;
    wire N__50047;
    wire N__50046;
    wire N__50045;
    wire N__50044;
    wire N__50041;
    wire N__50040;
    wire N__50039;
    wire N__50036;
    wire N__50035;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50027;
    wire N__50024;
    wire N__50023;
    wire N__50022;
    wire N__50021;
    wire N__50020;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50012;
    wire N__50009;
    wire N__50006;
    wire N__50003;
    wire N__49996;
    wire N__49989;
    wire N__49986;
    wire N__49985;
    wire N__49982;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49976;
    wire N__49975;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49963;
    wire N__49960;
    wire N__49957;
    wire N__49950;
    wire N__49945;
    wire N__49940;
    wire N__49937;
    wire N__49934;
    wire N__49931;
    wire N__49930;
    wire N__49927;
    wire N__49926;
    wire N__49923;
    wire N__49918;
    wire N__49915;
    wire N__49912;
    wire N__49903;
    wire N__49900;
    wire N__49891;
    wire N__49888;
    wire N__49881;
    wire N__49868;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49858;
    wire N__49855;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49835;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49827;
    wire N__49822;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49807;
    wire N__49802;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49792;
    wire N__49789;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49764;
    wire N__49761;
    wire N__49760;
    wire N__49759;
    wire N__49758;
    wire N__49757;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49748;
    wire N__49747;
    wire N__49746;
    wire N__49743;
    wire N__49738;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49718;
    wire N__49715;
    wire N__49712;
    wire N__49709;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49689;
    wire N__49686;
    wire N__49683;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49658;
    wire N__49655;
    wire N__49652;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49638;
    wire N__49635;
    wire N__49632;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49617;
    wire N__49616;
    wire N__49615;
    wire N__49614;
    wire N__49613;
    wire N__49612;
    wire N__49611;
    wire N__49610;
    wire N__49609;
    wire N__49608;
    wire N__49607;
    wire N__49606;
    wire N__49605;
    wire N__49604;
    wire N__49603;
    wire N__49602;
    wire N__49601;
    wire N__49600;
    wire N__49599;
    wire N__49598;
    wire N__49597;
    wire N__49596;
    wire N__49595;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49588;
    wire N__49587;
    wire N__49586;
    wire N__49585;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49573;
    wire N__49572;
    wire N__49571;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49564;
    wire N__49563;
    wire N__49562;
    wire N__49561;
    wire N__49560;
    wire N__49559;
    wire N__49558;
    wire N__49557;
    wire N__49556;
    wire N__49555;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49551;
    wire N__49550;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49529;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49519;
    wire N__49518;
    wire N__49517;
    wire N__49516;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49512;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49495;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49462;
    wire N__49459;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49441;
    wire N__49438;
    wire N__49435;
    wire N__49432;
    wire N__49429;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49411;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49070;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49052;
    wire N__49049;
    wire N__49046;
    wire N__49043;
    wire N__49042;
    wire N__49039;
    wire N__49038;
    wire N__49035;
    wire N__49034;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49024;
    wire N__49023;
    wire N__49022;
    wire N__49019;
    wire N__49016;
    wire N__49015;
    wire N__49014;
    wire N__49011;
    wire N__49010;
    wire N__49005;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48993;
    wire N__48990;
    wire N__48989;
    wire N__48988;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48980;
    wire N__48979;
    wire N__48978;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48966;
    wire N__48965;
    wire N__48962;
    wire N__48961;
    wire N__48958;
    wire N__48957;
    wire N__48956;
    wire N__48953;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48911;
    wire N__48910;
    wire N__48905;
    wire N__48900;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48886;
    wire N__48881;
    wire N__48876;
    wire N__48869;
    wire N__48864;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48850;
    wire N__48839;
    wire N__48836;
    wire N__48831;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48812;
    wire N__48805;
    wire N__48794;
    wire N__48791;
    wire N__48788;
    wire N__48785;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48774;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48755;
    wire N__48752;
    wire N__48749;
    wire N__48746;
    wire N__48743;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48724;
    wire N__48719;
    wire N__48716;
    wire N__48713;
    wire N__48710;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48693;
    wire N__48690;
    wire N__48683;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48671;
    wire N__48668;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48660;
    wire N__48657;
    wire N__48654;
    wire N__48651;
    wire N__48648;
    wire N__48645;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48612;
    wire N__48609;
    wire N__48606;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48590;
    wire N__48587;
    wire N__48584;
    wire N__48581;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48557;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48535;
    wire N__48530;
    wire N__48527;
    wire N__48524;
    wire N__48521;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48482;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48458;
    wire N__48455;
    wire N__48452;
    wire N__48449;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48434;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48412;
    wire N__48409;
    wire N__48408;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48391;
    wire N__48386;
    wire N__48381;
    wire N__48378;
    wire N__48371;
    wire N__48370;
    wire N__48367;
    wire N__48362;
    wire N__48359;
    wire N__48356;
    wire N__48355;
    wire N__48354;
    wire N__48351;
    wire N__48348;
    wire N__48345;
    wire N__48344;
    wire N__48341;
    wire N__48336;
    wire N__48333;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48314;
    wire N__48311;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48290;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48230;
    wire N__48229;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48211;
    wire N__48210;
    wire N__48209;
    wire N__48208;
    wire N__48207;
    wire N__48206;
    wire N__48203;
    wire N__48200;
    wire N__48199;
    wire N__48194;
    wire N__48193;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48185;
    wire N__48180;
    wire N__48177;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48170;
    wire N__48169;
    wire N__48166;
    wire N__48165;
    wire N__48162;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48136;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48110;
    wire N__48107;
    wire N__48106;
    wire N__48105;
    wire N__48104;
    wire N__48099;
    wire N__48096;
    wire N__48091;
    wire N__48088;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48081;
    wire N__48074;
    wire N__48069;
    wire N__48066;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48047;
    wire N__48044;
    wire N__48043;
    wire N__48042;
    wire N__48041;
    wire N__48040;
    wire N__48037;
    wire N__48032;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47990;
    wire N__47989;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47971;
    wire N__47966;
    wire N__47963;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47943;
    wire N__47936;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47918;
    wire N__47915;
    wire N__47912;
    wire N__47907;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47886;
    wire N__47885;
    wire N__47884;
    wire N__47883;
    wire N__47880;
    wire N__47875;
    wire N__47872;
    wire N__47865;
    wire N__47860;
    wire N__47853;
    wire N__47846;
    wire N__47843;
    wire N__47842;
    wire N__47839;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47823;
    wire N__47816;
    wire N__47809;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47713;
    wire N__47712;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47645;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47588;
    wire N__47585;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47575;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47552;
    wire N__47549;
    wire N__47548;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47538;
    wire N__47535;
    wire N__47528;
    wire N__47525;
    wire N__47524;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47497;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47477;
    wire N__47474;
    wire N__47471;
    wire N__47468;
    wire N__47467;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47447;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47423;
    wire N__47420;
    wire N__47419;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47392;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47369;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47360;
    wire N__47355;
    wire N__47352;
    wire N__47345;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47324;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47303;
    wire N__47300;
    wire N__47299;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47279;
    wire N__47276;
    wire N__47275;
    wire N__47272;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47249;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47225;
    wire N__47222;
    wire N__47221;
    wire N__47220;
    wire N__47215;
    wire N__47212;
    wire N__47209;
    wire N__47204;
    wire N__47201;
    wire N__47198;
    wire N__47197;
    wire N__47196;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47173;
    wire N__47172;
    wire N__47167;
    wire N__47164;
    wire N__47163;
    wire N__47160;
    wire N__47155;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47114;
    wire N__47111;
    wire N__47108;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47086;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47014;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47002;
    wire N__46997;
    wire N__46996;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46986;
    wire N__46979;
    wire N__46978;
    wire N__46977;
    wire N__46976;
    wire N__46973;
    wire N__46966;
    wire N__46961;
    wire N__46958;
    wire N__46955;
    wire N__46954;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46935;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46889;
    wire N__46886;
    wire N__46883;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46871;
    wire N__46868;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46820;
    wire N__46817;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46796;
    wire N__46795;
    wire N__46792;
    wire N__46789;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46783;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46771;
    wire N__46768;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46760;
    wire N__46755;
    wire N__46754;
    wire N__46753;
    wire N__46752;
    wire N__46749;
    wire N__46746;
    wire N__46745;
    wire N__46742;
    wire N__46733;
    wire N__46730;
    wire N__46725;
    wire N__46720;
    wire N__46713;
    wire N__46708;
    wire N__46705;
    wire N__46700;
    wire N__46693;
    wire N__46690;
    wire N__46679;
    wire N__46678;
    wire N__46677;
    wire N__46670;
    wire N__46667;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46663;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46646;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46636;
    wire N__46633;
    wire N__46632;
    wire N__46631;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46605;
    wire N__46602;
    wire N__46601;
    wire N__46598;
    wire N__46593;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46585;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46577;
    wire N__46574;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46523;
    wire N__46518;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46490;
    wire N__46481;
    wire N__46478;
    wire N__46477;
    wire N__46476;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46410;
    wire N__46405;
    wire N__46402;
    wire N__46397;
    wire N__46396;
    wire N__46395;
    wire N__46394;
    wire N__46391;
    wire N__46390;
    wire N__46389;
    wire N__46388;
    wire N__46387;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46367;
    wire N__46366;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46351;
    wire N__46348;
    wire N__46343;
    wire N__46342;
    wire N__46341;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46333;
    wire N__46332;
    wire N__46329;
    wire N__46328;
    wire N__46325;
    wire N__46322;
    wire N__46321;
    wire N__46312;
    wire N__46311;
    wire N__46310;
    wire N__46309;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46305;
    wire N__46304;
    wire N__46301;
    wire N__46294;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46265;
    wire N__46262;
    wire N__46257;
    wire N__46256;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46248;
    wire N__46245;
    wire N__46244;
    wire N__46243;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46221;
    wire N__46212;
    wire N__46209;
    wire N__46200;
    wire N__46195;
    wire N__46194;
    wire N__46193;
    wire N__46192;
    wire N__46191;
    wire N__46190;
    wire N__46189;
    wire N__46188;
    wire N__46187;
    wire N__46176;
    wire N__46171;
    wire N__46170;
    wire N__46161;
    wire N__46158;
    wire N__46157;
    wire N__46156;
    wire N__46155;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46145;
    wire N__46144;
    wire N__46141;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46106;
    wire N__46097;
    wire N__46094;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46069;
    wire N__46062;
    wire N__46059;
    wire N__46054;
    wire N__46049;
    wire N__46046;
    wire N__46041;
    wire N__46038;
    wire N__46031;
    wire N__46030;
    wire N__46027;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46001;
    wire N__45998;
    wire N__45997;
    wire N__45994;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45977;
    wire N__45974;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45964;
    wire N__45961;
    wire N__45958;
    wire N__45955;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45940;
    wire N__45935;
    wire N__45934;
    wire N__45933;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45925;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45898;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45890;
    wire N__45889;
    wire N__45884;
    wire N__45881;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45842;
    wire N__45841;
    wire N__45840;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45832;
    wire N__45831;
    wire N__45830;
    wire N__45829;
    wire N__45826;
    wire N__45823;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45803;
    wire N__45802;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45756;
    wire N__45753;
    wire N__45748;
    wire N__45731;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45658;
    wire N__45655;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45629;
    wire N__45628;
    wire N__45627;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45601;
    wire N__45598;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45572;
    wire N__45571;
    wire N__45570;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45520;
    wire N__45517;
    wire N__45512;
    wire N__45511;
    wire N__45510;
    wire N__45503;
    wire N__45500;
    wire N__45499;
    wire N__45498;
    wire N__45495;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45478;
    wire N__45477;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45444;
    wire N__45441;
    wire N__45440;
    wire N__45435;
    wire N__45430;
    wire N__45425;
    wire N__45424;
    wire N__45423;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45411;
    wire N__45406;
    wire N__45403;
    wire N__45396;
    wire N__45393;
    wire N__45388;
    wire N__45385;
    wire N__45368;
    wire N__45367;
    wire N__45366;
    wire N__45363;
    wire N__45362;
    wire N__45361;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45353;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45311;
    wire N__45310;
    wire N__45309;
    wire N__45308;
    wire N__45305;
    wire N__45304;
    wire N__45299;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45277;
    wire N__45274;
    wire N__45269;
    wire N__45254;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45226;
    wire N__45221;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45211;
    wire N__45202;
    wire N__45199;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45185;
    wire N__45182;
    wire N__45181;
    wire N__45180;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45164;
    wire N__45161;
    wire N__45160;
    wire N__45159;
    wire N__45158;
    wire N__45157;
    wire N__45156;
    wire N__45153;
    wire N__45152;
    wire N__45149;
    wire N__45148;
    wire N__45145;
    wire N__45144;
    wire N__45141;
    wire N__45140;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45131;
    wire N__45128;
    wire N__45127;
    wire N__45126;
    wire N__45125;
    wire N__45124;
    wire N__45123;
    wire N__45122;
    wire N__45121;
    wire N__45118;
    wire N__45111;
    wire N__45106;
    wire N__45101;
    wire N__45092;
    wire N__45091;
    wire N__45090;
    wire N__45089;
    wire N__45086;
    wire N__45085;
    wire N__45082;
    wire N__45079;
    wire N__45078;
    wire N__45075;
    wire N__45066;
    wire N__45063;
    wire N__45062;
    wire N__45061;
    wire N__45060;
    wire N__45057;
    wire N__45056;
    wire N__45053;
    wire N__45052;
    wire N__45051;
    wire N__45046;
    wire N__45043;
    wire N__45038;
    wire N__45035;
    wire N__45032;
    wire N__45031;
    wire N__45030;
    wire N__45029;
    wire N__45028;
    wire N__45025;
    wire N__45024;
    wire N__45023;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45009;
    wire N__45004;
    wire N__44995;
    wire N__44984;
    wire N__44977;
    wire N__44968;
    wire N__44959;
    wire N__44956;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44930;
    wire N__44927;
    wire N__44926;
    wire N__44925;
    wire N__44924;
    wire N__44923;
    wire N__44922;
    wire N__44921;
    wire N__44920;
    wire N__44919;
    wire N__44918;
    wire N__44917;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44910;
    wire N__44909;
    wire N__44904;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44896;
    wire N__44893;
    wire N__44888;
    wire N__44879;
    wire N__44874;
    wire N__44865;
    wire N__44862;
    wire N__44861;
    wire N__44860;
    wire N__44859;
    wire N__44858;
    wire N__44857;
    wire N__44854;
    wire N__44853;
    wire N__44852;
    wire N__44851;
    wire N__44850;
    wire N__44849;
    wire N__44848;
    wire N__44847;
    wire N__44846;
    wire N__44845;
    wire N__44844;
    wire N__44843;
    wire N__44842;
    wire N__44841;
    wire N__44840;
    wire N__44839;
    wire N__44836;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44832;
    wire N__44831;
    wire N__44830;
    wire N__44829;
    wire N__44828;
    wire N__44827;
    wire N__44826;
    wire N__44819;
    wire N__44816;
    wire N__44811;
    wire N__44806;
    wire N__44801;
    wire N__44796;
    wire N__44793;
    wire N__44788;
    wire N__44787;
    wire N__44786;
    wire N__44783;
    wire N__44772;
    wire N__44757;
    wire N__44748;
    wire N__44739;
    wire N__44726;
    wire N__44725;
    wire N__44724;
    wire N__44723;
    wire N__44722;
    wire N__44711;
    wire N__44708;
    wire N__44703;
    wire N__44700;
    wire N__44689;
    wire N__44684;
    wire N__44679;
    wire N__44670;
    wire N__44669;
    wire N__44668;
    wire N__44667;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44641;
    wire N__44634;
    wire N__44627;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44503;
    wire N__44502;
    wire N__44501;
    wire N__44500;
    wire N__44499;
    wire N__44498;
    wire N__44495;
    wire N__44494;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44490;
    wire N__44489;
    wire N__44488;
    wire N__44477;
    wire N__44474;
    wire N__44473;
    wire N__44464;
    wire N__44455;
    wire N__44452;
    wire N__44449;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44427;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44411;
    wire N__44410;
    wire N__44409;
    wire N__44408;
    wire N__44405;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44383;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44260;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44245;
    wire N__44244;
    wire N__44241;
    wire N__44236;
    wire N__44231;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44219;
    wire N__44216;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44202;
    wire N__44197;
    wire N__44194;
    wire N__44189;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44177;
    wire N__44174;
    wire N__44171;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44163;
    wire N__44158;
    wire N__44155;
    wire N__44150;
    wire N__44147;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44101;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44083;
    wire N__44078;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44054;
    wire N__44051;
    wire N__44048;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44038;
    wire N__44035;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44017;
    wire N__44012;
    wire N__44011;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44003;
    wire N__44000;
    wire N__43995;
    wire N__43992;
    wire N__43987;
    wire N__43982;
    wire N__43979;
    wire N__43978;
    wire N__43977;
    wire N__43974;
    wire N__43969;
    wire N__43966;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43954;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43946;
    wire N__43945;
    wire N__43944;
    wire N__43941;
    wire N__43936;
    wire N__43929;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43903;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43886;
    wire N__43883;
    wire N__43882;
    wire N__43881;
    wire N__43880;
    wire N__43875;
    wire N__43872;
    wire N__43871;
    wire N__43870;
    wire N__43869;
    wire N__43866;
    wire N__43861;
    wire N__43856;
    wire N__43853;
    wire N__43852;
    wire N__43849;
    wire N__43844;
    wire N__43841;
    wire N__43840;
    wire N__43839;
    wire N__43836;
    wire N__43835;
    wire N__43834;
    wire N__43833;
    wire N__43832;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43811;
    wire N__43806;
    wire N__43801;
    wire N__43784;
    wire N__43783;
    wire N__43782;
    wire N__43779;
    wire N__43778;
    wire N__43777;
    wire N__43776;
    wire N__43773;
    wire N__43772;
    wire N__43767;
    wire N__43766;
    wire N__43763;
    wire N__43762;
    wire N__43761;
    wire N__43758;
    wire N__43757;
    wire N__43754;
    wire N__43753;
    wire N__43750;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43739;
    wire N__43736;
    wire N__43729;
    wire N__43728;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43712;
    wire N__43711;
    wire N__43710;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43696;
    wire N__43693;
    wire N__43688;
    wire N__43683;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43662;
    wire N__43655;
    wire N__43646;
    wire N__43643;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43504;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43375;
    wire N__43374;
    wire N__43373;
    wire N__43372;
    wire N__43367;
    wire N__43366;
    wire N__43363;
    wire N__43362;
    wire N__43361;
    wire N__43360;
    wire N__43359;
    wire N__43358;
    wire N__43355;
    wire N__43354;
    wire N__43353;
    wire N__43352;
    wire N__43351;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43331;
    wire N__43326;
    wire N__43323;
    wire N__43318;
    wire N__43311;
    wire N__43310;
    wire N__43309;
    wire N__43308;
    wire N__43305;
    wire N__43300;
    wire N__43287;
    wire N__43280;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43243;
    wire N__43242;
    wire N__43241;
    wire N__43240;
    wire N__43239;
    wire N__43238;
    wire N__43237;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43223;
    wire N__43222;
    wire N__43221;
    wire N__43220;
    wire N__43219;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43204;
    wire N__43201;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43178;
    wire N__43177;
    wire N__43176;
    wire N__43175;
    wire N__43172;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43156;
    wire N__43149;
    wire N__43146;
    wire N__43141;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43125;
    wire N__43122;
    wire N__43117;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43067;
    wire N__43064;
    wire N__43061;
    wire N__43058;
    wire N__43055;
    wire N__43052;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42983;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42829;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42817;
    wire N__42816;
    wire N__42815;
    wire N__42814;
    wire N__42811;
    wire N__42810;
    wire N__42809;
    wire N__42806;
    wire N__42805;
    wire N__42804;
    wire N__42803;
    wire N__42802;
    wire N__42801;
    wire N__42800;
    wire N__42799;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42780;
    wire N__42777;
    wire N__42776;
    wire N__42775;
    wire N__42772;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42764;
    wire N__42761;
    wire N__42756;
    wire N__42751;
    wire N__42744;
    wire N__42737;
    wire N__42734;
    wire N__42727;
    wire N__42726;
    wire N__42723;
    wire N__42716;
    wire N__42713;
    wire N__42704;
    wire N__42699;
    wire N__42696;
    wire N__42695;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42683;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42671;
    wire N__42662;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42641;
    wire N__42640;
    wire N__42639;
    wire N__42634;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42616;
    wire N__42611;
    wire N__42610;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42602;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42571;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42559;
    wire N__42556;
    wire N__42553;
    wire N__42548;
    wire N__42543;
    wire N__42540;
    wire N__42535;
    wire N__42532;
    wire N__42527;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42509;
    wire N__42506;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42437;
    wire N__42434;
    wire N__42431;
    wire N__42428;
    wire N__42425;
    wire N__42424;
    wire N__42423;
    wire N__42422;
    wire N__42421;
    wire N__42420;
    wire N__42419;
    wire N__42412;
    wire N__42409;
    wire N__42402;
    wire N__42395;
    wire N__42392;
    wire N__42389;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42338;
    wire N__42335;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42277;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42257;
    wire N__42254;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42214;
    wire N__42209;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42201;
    wire N__42196;
    wire N__42189;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42175;
    wire N__42174;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42155;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42112;
    wire N__42107;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42087;
    wire N__42086;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42059;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42045;
    wire N__42040;
    wire N__42037;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42020;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__41996;
    wire N__41995;
    wire N__41992;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41975;
    wire N__41972;
    wire N__41971;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41920;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41891;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41815;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41792;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41779;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41759;
    wire N__41756;
    wire N__41753;
    wire N__41750;
    wire N__41747;
    wire N__41746;
    wire N__41745;
    wire N__41742;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41730;
    wire N__41723;
    wire N__41722;
    wire N__41721;
    wire N__41720;
    wire N__41717;
    wire N__41714;
    wire N__41709;
    wire N__41702;
    wire N__41699;
    wire N__41696;
    wire N__41693;
    wire N__41692;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41668;
    wire N__41663;
    wire N__41660;
    wire N__41659;
    wire N__41656;
    wire N__41653;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41602;
    wire N__41599;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41581;
    wire N__41580;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41530;
    wire N__41529;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41485;
    wire N__41484;
    wire N__41481;
    wire N__41476;
    wire N__41473;
    wire N__41468;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41443;
    wire N__41442;
    wire N__41441;
    wire N__41440;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41424;
    wire N__41417;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41409;
    wire N__41406;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41388;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41368;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41353;
    wire N__41350;
    wire N__41345;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41337;
    wire N__41334;
    wire N__41329;
    wire N__41328;
    wire N__41327;
    wire N__41326;
    wire N__41325;
    wire N__41324;
    wire N__41323;
    wire N__41318;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41298;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41275;
    wire N__41274;
    wire N__41271;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41263;
    wire N__41262;
    wire N__41261;
    wire N__41256;
    wire N__41251;
    wire N__41248;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41225;
    wire N__41222;
    wire N__41221;
    wire N__41220;
    wire N__41217;
    wire N__41212;
    wire N__41207;
    wire N__41204;
    wire N__41203;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41175;
    wire N__41168;
    wire N__41167;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41150;
    wire N__41149;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41117;
    wire N__41114;
    wire N__41113;
    wire N__41108;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41087;
    wire N__41084;
    wire N__41083;
    wire N__41082;
    wire N__41081;
    wire N__41078;
    wire N__41077;
    wire N__41074;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41054;
    wire N__41053;
    wire N__41052;
    wire N__41045;
    wire N__41042;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40993;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40967;
    wire N__40964;
    wire N__40963;
    wire N__40962;
    wire N__40959;
    wire N__40954;
    wire N__40951;
    wire N__40946;
    wire N__40943;
    wire N__40942;
    wire N__40941;
    wire N__40938;
    wire N__40933;
    wire N__40928;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40888;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40873;
    wire N__40870;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40796;
    wire N__40793;
    wire N__40790;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40759;
    wire N__40758;
    wire N__40757;
    wire N__40752;
    wire N__40751;
    wire N__40750;
    wire N__40749;
    wire N__40748;
    wire N__40743;
    wire N__40740;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40712;
    wire N__40711;
    wire N__40708;
    wire N__40707;
    wire N__40706;
    wire N__40705;
    wire N__40704;
    wire N__40701;
    wire N__40700;
    wire N__40695;
    wire N__40694;
    wire N__40693;
    wire N__40692;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40682;
    wire N__40677;
    wire N__40676;
    wire N__40673;
    wire N__40670;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40643;
    wire N__40638;
    wire N__40635;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40605;
    wire N__40596;
    wire N__40589;
    wire N__40586;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40575;
    wire N__40570;
    wire N__40567;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40532;
    wire N__40529;
    wire N__40528;
    wire N__40525;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40503;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40465;
    wire N__40464;
    wire N__40461;
    wire N__40456;
    wire N__40451;
    wire N__40448;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40426;
    wire N__40425;
    wire N__40422;
    wire N__40417;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40400;
    wire N__40397;
    wire N__40396;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40379;
    wire N__40378;
    wire N__40375;
    wire N__40370;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40324;
    wire N__40317;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40301;
    wire N__40300;
    wire N__40299;
    wire N__40296;
    wire N__40291;
    wire N__40288;
    wire N__40283;
    wire N__40274;
    wire N__40273;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40262;
    wire N__40261;
    wire N__40258;
    wire N__40257;
    wire N__40256;
    wire N__40255;
    wire N__40254;
    wire N__40251;
    wire N__40250;
    wire N__40247;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40200;
    wire N__40195;
    wire N__40194;
    wire N__40189;
    wire N__40184;
    wire N__40179;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40156;
    wire N__40151;
    wire N__40142;
    wire N__40141;
    wire N__40140;
    wire N__40139;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40122;
    wire N__40121;
    wire N__40116;
    wire N__40111;
    wire N__40110;
    wire N__40107;
    wire N__40106;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40041;
    wire N__40040;
    wire N__40037;
    wire N__40032;
    wire N__40027;
    wire N__40022;
    wire N__40013;
    wire N__40012;
    wire N__40011;
    wire N__40010;
    wire N__40007;
    wire N__40006;
    wire N__40005;
    wire N__40002;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39994;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39983;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39975;
    wire N__39974;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39944;
    wire N__39939;
    wire N__39934;
    wire N__39931;
    wire N__39930;
    wire N__39925;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39853;
    wire N__39848;
    wire N__39845;
    wire N__39844;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39769;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39761;
    wire N__39760;
    wire N__39759;
    wire N__39756;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39713;
    wire N__39710;
    wire N__39707;
    wire N__39706;
    wire N__39699;
    wire N__39698;
    wire N__39697;
    wire N__39692;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39669;
    wire N__39664;
    wire N__39653;
    wire N__39652;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39634;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39626;
    wire N__39625;
    wire N__39620;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39598;
    wire N__39595;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39581;
    wire N__39578;
    wire N__39577;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39541;
    wire N__39538;
    wire N__39527;
    wire N__39526;
    wire N__39525;
    wire N__39522;
    wire N__39519;
    wire N__39516;
    wire N__39513;
    wire N__39512;
    wire N__39509;
    wire N__39504;
    wire N__39501;
    wire N__39500;
    wire N__39499;
    wire N__39498;
    wire N__39497;
    wire N__39492;
    wire N__39489;
    wire N__39488;
    wire N__39487;
    wire N__39484;
    wire N__39483;
    wire N__39478;
    wire N__39475;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39467;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39445;
    wire N__39440;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39405;
    wire N__39394;
    wire N__39391;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39366;
    wire N__39365;
    wire N__39364;
    wire N__39363;
    wire N__39362;
    wire N__39359;
    wire N__39356;
    wire N__39353;
    wire N__39348;
    wire N__39345;
    wire N__39344;
    wire N__39343;
    wire N__39340;
    wire N__39335;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39305;
    wire N__39302;
    wire N__39299;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39267;
    wire N__39262;
    wire N__39251;
    wire N__39250;
    wire N__39247;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39193;
    wire N__39190;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39172;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39157;
    wire N__39152;
    wire N__39149;
    wire N__39148;
    wire N__39145;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39071;
    wire N__39068;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39032;
    wire N__39031;
    wire N__39028;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38975;
    wire N__38974;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38962;
    wire N__38961;
    wire N__38956;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38939;
    wire N__38938;
    wire N__38937;
    wire N__38936;
    wire N__38931;
    wire N__38926;
    wire N__38925;
    wire N__38924;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38900;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38892;
    wire N__38887;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38841;
    wire N__38836;
    wire N__38833;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38815;
    wire N__38810;
    wire N__38807;
    wire N__38806;
    wire N__38803;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38780;
    wire N__38777;
    wire N__38776;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38674;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38614;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38558;
    wire N__38555;
    wire N__38554;
    wire N__38551;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38525;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38498;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38485;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38465;
    wire N__38464;
    wire N__38461;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38443;
    wire N__38440;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38428;
    wire N__38425;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38399;
    wire N__38398;
    wire N__38393;
    wire N__38390;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38380;
    wire N__38375;
    wire N__38372;
    wire N__38371;
    wire N__38370;
    wire N__38365;
    wire N__38362;
    wire N__38361;
    wire N__38360;
    wire N__38357;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38340;
    wire N__38337;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38318;
    wire N__38317;
    wire N__38316;
    wire N__38315;
    wire N__38314;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38285;
    wire N__38284;
    wire N__38281;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38258;
    wire N__38257;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38208;
    wire N__38201;
    wire N__38200;
    wire N__38195;
    wire N__38192;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38180;
    wire N__38179;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38173;
    wire N__38172;
    wire N__38171;
    wire N__38170;
    wire N__38165;
    wire N__38152;
    wire N__38147;
    wire N__38144;
    wire N__38143;
    wire N__38142;
    wire N__38139;
    wire N__38138;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38118;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38100;
    wire N__38097;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38075;
    wire N__38074;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38039;
    wire N__38036;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37996;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37966;
    wire N__37965;
    wire N__37960;
    wire N__37957;
    wire N__37952;
    wire N__37951;
    wire N__37948;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37894;
    wire N__37893;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37864;
    wire N__37859;
    wire N__37856;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37844;
    wire N__37843;
    wire N__37842;
    wire N__37841;
    wire N__37838;
    wire N__37833;
    wire N__37830;
    wire N__37825;
    wire N__37820;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37795;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37756;
    wire N__37755;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37723;
    wire N__37718;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37606;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37552;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37477;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37459;
    wire N__37458;
    wire N__37455;
    wire N__37450;
    wire N__37445;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37432;
    wire N__37429;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37129;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37114;
    wire N__37113;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37062;
    wire N__37059;
    wire N__37052;
    wire N__37049;
    wire N__37048;
    wire N__37045;
    wire N__37044;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37034;
    wire N__37031;
    wire N__37026;
    wire N__37023;
    wire N__37022;
    wire N__37019;
    wire N__37014;
    wire N__37011;
    wire N__37010;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36996;
    wire N__36993;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36971;
    wire N__36970;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36935;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36923;
    wire N__36920;
    wire N__36919;
    wire N__36916;
    wire N__36909;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36884;
    wire N__36881;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36857;
    wire N__36852;
    wire N__36849;
    wire N__36848;
    wire N__36845;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36832;
    wire N__36829;
    wire N__36822;
    wire N__36817;
    wire N__36814;
    wire N__36809;
    wire N__36808;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36789;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36767;
    wire N__36760;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36741;
    wire N__36738;
    wire N__36731;
    wire N__36730;
    wire N__36727;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36628;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36620;
    wire N__36617;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36580;
    wire N__36575;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36548;
    wire N__36545;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36533;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36521;
    wire N__36520;
    wire N__36517;
    wire N__36516;
    wire N__36511;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36485;
    wire N__36484;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36455;
    wire N__36454;
    wire N__36453;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36441;
    wire N__36440;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36416;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36401;
    wire N__36398;
    wire N__36397;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36334;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36196;
    wire N__36193;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36144;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36091;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36067;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36020;
    wire N__36019;
    wire N__36018;
    wire N__36011;
    wire N__36008;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35977;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35962;
    wire N__35957;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35949;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35937;
    wire N__35930;
    wire N__35929;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35897;
    wire N__35896;
    wire N__35895;
    wire N__35894;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35878;
    wire N__35877;
    wire N__35868;
    wire N__35867;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35792;
    wire N__35789;
    wire N__35788;
    wire N__35787;
    wire N__35784;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35758;
    wire N__35753;
    wire N__35750;
    wire N__35749;
    wire N__35748;
    wire N__35747;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35731;
    wire N__35728;
    wire N__35727;
    wire N__35724;
    wire N__35721;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35702;
    wire N__35701;
    wire N__35696;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35665;
    wire N__35664;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35648;
    wire N__35647;
    wire N__35642;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35632;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35620;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35521;
    wire N__35518;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35284;
    wire N__35283;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35269;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35254;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35228;
    wire N__35225;
    wire N__35224;
    wire N__35223;
    wire N__35216;
    wire N__35213;
    wire N__35212;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35196;
    wire N__35189;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35177;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35165;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35150;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35138;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35126;
    wire N__35125;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35108;
    wire N__35105;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35057;
    wire N__35056;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35017;
    wire N__35016;
    wire N__35015;
    wire N__35012;
    wire N__35005;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34940;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34925;
    wire N__34924;
    wire N__34923;
    wire N__34918;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34892;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34848;
    wire N__34847;
    wire N__34842;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34822;
    wire N__34821;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34805;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34790;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34687;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34633;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34610;
    wire N__34609;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34575;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34556;
    wire N__34551;
    wire N__34548;
    wire N__34543;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34503;
    wire N__34502;
    wire N__34497;
    wire N__34494;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34472;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34456;
    wire N__34453;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34413;
    wire N__34406;
    wire N__34403;
    wire N__34402;
    wire N__34401;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34383;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34244;
    wire N__34237;
    wire N__34232;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34208;
    wire N__34205;
    wire N__34204;
    wire N__34201;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34141;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34108;
    wire N__34107;
    wire N__34104;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34088;
    wire N__34085;
    wire N__34084;
    wire N__34083;
    wire N__34080;
    wire N__34075;
    wire N__34072;
    wire N__34067;
    wire N__34066;
    wire N__34065;
    wire N__34062;
    wire N__34057;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__34000;
    wire N__33999;
    wire N__33996;
    wire N__33991;
    wire N__33986;
    wire N__33983;
    wire N__33982;
    wire N__33981;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33926;
    wire N__33923;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33911;
    wire N__33910;
    wire N__33907;
    wire N__33902;
    wire N__33899;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33887;
    wire N__33884;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33761;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33723;
    wire N__33718;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33685;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33666;
    wire N__33665;
    wire N__33664;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33642;
    wire N__33639;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33617;
    wire N__33602;
    wire N__33599;
    wire N__33598;
    wire N__33597;
    wire N__33594;
    wire N__33593;
    wire N__33590;
    wire N__33589;
    wire N__33588;
    wire N__33575;
    wire N__33574;
    wire N__33573;
    wire N__33572;
    wire N__33569;
    wire N__33564;
    wire N__33561;
    wire N__33554;
    wire N__33553;
    wire N__33550;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33519;
    wire N__33514;
    wire N__33511;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33394;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33386;
    wire N__33383;
    wire N__33378;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33347;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33308;
    wire N__33305;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33286;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33256;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33227;
    wire N__33226;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33197;
    wire N__33196;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33173;
    wire N__33172;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33158;
    wire N__33157;
    wire N__33154;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33100;
    wire N__33097;
    wire N__33096;
    wire N__33095;
    wire N__33092;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33054;
    wire N__33049;
    wire N__33046;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33028;
    wire N__33027;
    wire N__33024;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33006;
    wire N__33005;
    wire N__33004;
    wire N__32999;
    wire N__32996;
    wire N__32991;
    wire N__32988;
    wire N__32983;
    wire N__32980;
    wire N__32969;
    wire N__32968;
    wire N__32967;
    wire N__32962;
    wire N__32959;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32936;
    wire N__32933;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32907;
    wire N__32904;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32832;
    wire N__32831;
    wire N__32828;
    wire N__32823;
    wire N__32820;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32776;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32734;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32653;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32617;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32519;
    wire N__32516;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32473;
    wire N__32468;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32416;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32394;
    wire N__32387;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32370;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32342;
    wire N__32341;
    wire N__32340;
    wire N__32339;
    wire N__32336;
    wire N__32335;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32300;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32221;
    wire N__32218;
    wire N__32217;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32196;
    wire N__32189;
    wire N__32188;
    wire N__32185;
    wire N__32180;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32135;
    wire N__32132;
    wire N__32131;
    wire N__32130;
    wire N__32127;
    wire N__32122;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32085;
    wire N__32082;
    wire N__32077;
    wire N__32072;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32047;
    wire N__32046;
    wire N__32043;
    wire N__32038;
    wire N__32033;
    wire N__32030;
    wire N__32029;
    wire N__32028;
    wire N__32027;
    wire N__32026;
    wire N__32025;
    wire N__32024;
    wire N__32023;
    wire N__32022;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31979;
    wire N__31976;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31954;
    wire N__31951;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31943;
    wire N__31940;
    wire N__31933;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31910;
    wire N__31907;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31892;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31870;
    wire N__31867;
    wire N__31856;
    wire N__31855;
    wire N__31854;
    wire N__31853;
    wire N__31852;
    wire N__31851;
    wire N__31844;
    wire N__31843;
    wire N__31842;
    wire N__31839;
    wire N__31834;
    wire N__31833;
    wire N__31830;
    wire N__31825;
    wire N__31820;
    wire N__31817;
    wire N__31808;
    wire N__31807;
    wire N__31804;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31774;
    wire N__31771;
    wire N__31770;
    wire N__31769;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31725;
    wire N__31724;
    wire N__31715;
    wire N__31714;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31703;
    wire N__31702;
    wire N__31701;
    wire N__31700;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31682;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31664;
    wire N__31663;
    wire N__31662;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31642;
    wire N__31641;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31626;
    wire N__31623;
    wire N__31616;
    wire N__31611;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31592;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31517;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31484;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31466;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31445;
    wire N__31444;
    wire N__31443;
    wire N__31442;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31415;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31333;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31310;
    wire N__31307;
    wire N__31306;
    wire N__31305;
    wire N__31304;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31293;
    wire N__31292;
    wire N__31291;
    wire N__31286;
    wire N__31279;
    wire N__31272;
    wire N__31265;
    wire N__31262;
    wire N__31261;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31246;
    wire N__31241;
    wire N__31240;
    wire N__31239;
    wire N__31238;
    wire N__31237;
    wire N__31236;
    wire N__31235;
    wire N__31234;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31177;
    wire N__31174;
    wire N__31171;
    wire N__31168;
    wire N__31167;
    wire N__31164;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31147;
    wire N__31144;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31128;
    wire N__31125;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31101;
    wire N__31100;
    wire N__31099;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31074;
    wire N__31069;
    wire N__31066;
    wire N__31055;
    wire N__31054;
    wire N__31051;
    wire N__31050;
    wire N__31049;
    wire N__31048;
    wire N__31047;
    wire N__31046;
    wire N__31043;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31026;
    wire N__31025;
    wire N__31022;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31011;
    wire N__31010;
    wire N__31009;
    wire N__30996;
    wire N__30991;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30975;
    wire N__30970;
    wire N__30967;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30895;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30854;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30839;
    wire N__30836;
    wire N__30833;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30825;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30761;
    wire N__30758;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30674;
    wire N__30671;
    wire N__30670;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30657;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30638;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30611;
    wire N__30610;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30567;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30547;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30511;
    wire N__30506;
    wire N__30505;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30492;
    wire N__30491;
    wire N__30490;
    wire N__30485;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30469;
    wire N__30466;
    wire N__30461;
    wire N__30460;
    wire N__30459;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30451;
    wire N__30448;
    wire N__30443;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30415;
    wire N__30410;
    wire N__30409;
    wire N__30408;
    wire N__30403;
    wire N__30400;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30354;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30263;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30248;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30236;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30224;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30212;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30197;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30185;
    wire N__30182;
    wire N__30181;
    wire N__30180;
    wire N__30177;
    wire N__30172;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30144;
    wire N__30141;
    wire N__30140;
    wire N__30139;
    wire N__30138;
    wire N__30137;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30114;
    wire N__30101;
    wire N__30098;
    wire N__30097;
    wire N__30096;
    wire N__30089;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30077;
    wire N__30076;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30052;
    wire N__30047;
    wire N__30046;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30036;
    wire N__30033;
    wire N__30032;
    wire N__30031;
    wire N__30030;
    wire N__30027;
    wire N__30020;
    wire N__30011;
    wire N__30008;
    wire N__29999;
    wire N__29998;
    wire N__29997;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29985;
    wire N__29984;
    wire N__29983;
    wire N__29980;
    wire N__29973;
    wire N__29966;
    wire N__29963;
    wire N__29954;
    wire N__29953;
    wire N__29952;
    wire N__29951;
    wire N__29948;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29935;
    wire N__29934;
    wire N__29933;
    wire N__29928;
    wire N__29921;
    wire N__29912;
    wire N__29909;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29821;
    wire N__29820;
    wire N__29819;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29807;
    wire N__29804;
    wire N__29795;
    wire N__29792;
    wire N__29791;
    wire N__29790;
    wire N__29789;
    wire N__29788;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29773;
    wire N__29770;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29722;
    wire N__29721;
    wire N__29718;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29703;
    wire N__29696;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29660;
    wire N__29651;
    wire N__29648;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29636;
    wire N__29633;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29615;
    wire N__29612;
    wire N__29611;
    wire N__29608;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29580;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29449;
    wire N__29448;
    wire N__29445;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29315;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29300;
    wire N__29299;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29267;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29222;
    wire N__29221;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29210;
    wire N__29207;
    wire N__29206;
    wire N__29205;
    wire N__29204;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29196;
    wire N__29195;
    wire N__29192;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29171;
    wire N__29166;
    wire N__29161;
    wire N__29144;
    wire N__29141;
    wire N__29140;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29116;
    wire N__29113;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29099;
    wire N__29098;
    wire N__29097;
    wire N__29094;
    wire N__29089;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29017;
    wire N__29012;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28989;
    wire N__28982;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28974;
    wire N__28969;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28949;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28938;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28925;
    wire N__28916;
    wire N__28913;
    wire N__28912;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28856;
    wire N__28853;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28792;
    wire N__28791;
    wire N__28788;
    wire N__28783;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28770;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28745;
    wire N__28742;
    wire N__28741;
    wire N__28736;
    wire N__28731;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28716;
    wire N__28709;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28613;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28576;
    wire N__28573;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28538;
    wire N__28537;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28501;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28439;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28424;
    wire N__28421;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28409;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28368;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28279;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28147;
    wire N__28146;
    wire N__28143;
    wire N__28138;
    wire N__28137;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28121;
    wire N__28120;
    wire N__28119;
    wire N__28118;
    wire N__28115;
    wire N__28114;
    wire N__28109;
    wire N__28102;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28066;
    wire N__28063;
    wire N__28058;
    wire N__28055;
    wire N__28054;
    wire N__28053;
    wire N__28052;
    wire N__28051;
    wire N__28050;
    wire N__28047;
    wire N__28042;
    wire N__28037;
    wire N__28034;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__28000;
    wire N__27999;
    wire N__27998;
    wire N__27995;
    wire N__27990;
    wire N__27987;
    wire N__27980;
    wire N__27977;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27965;
    wire N__27964;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27947;
    wire N__27946;
    wire N__27943;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27925;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27894;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27870;
    wire N__27863;
    wire N__27856;
    wire N__27855;
    wire N__27854;
    wire N__27849;
    wire N__27844;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27785;
    wire N__27784;
    wire N__27781;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27715;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27700;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27685;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27670;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27655;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27610;
    wire N__27609;
    wire N__27608;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27604;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27578;
    wire N__27577;
    wire N__27574;
    wire N__27569;
    wire N__27568;
    wire N__27567;
    wire N__27564;
    wire N__27551;
    wire N__27546;
    wire N__27541;
    wire N__27538;
    wire N__27537;
    wire N__27536;
    wire N__27535;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27519;
    wire N__27516;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27478;
    wire N__27471;
    wire N__27468;
    wire N__27461;
    wire N__27458;
    wire N__27443;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27430;
    wire N__27425;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27376;
    wire N__27371;
    wire N__27362;
    wire N__27359;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27307;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27255;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27230;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27176;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27158;
    wire N__27155;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26991;
    wire N__26990;
    wire N__26987;
    wire N__26980;
    wire N__26975;
    wire N__26974;
    wire N__26971;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26939;
    wire N__26936;
    wire N__26935;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26917;
    wire N__26916;
    wire N__26915;
    wire N__26914;
    wire N__26913;
    wire N__26904;
    wire N__26903;
    wire N__26902;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26880;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26868;
    wire N__26865;
    wire N__26860;
    wire N__26857;
    wire N__26852;
    wire N__26851;
    wire N__26844;
    wire N__26835;
    wire N__26832;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26764;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26725;
    wire N__26720;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26702;
    wire N__26699;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26673;
    wire N__26668;
    wire N__26663;
    wire N__26660;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26588;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26573;
    wire N__26570;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26558;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26540;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26513;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26498;
    wire N__26495;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26485;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26441;
    wire N__26438;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26249;
    wire N__26246;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26234;
    wire N__26231;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26216;
    wire N__26213;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26201;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26193;
    wire N__26188;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26170;
    wire N__26165;
    wire N__26162;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26143;
    wire N__26142;
    wire N__26141;
    wire N__26138;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26116;
    wire N__26115;
    wire N__26114;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26009;
    wire N__26006;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25933;
    wire N__25930;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25714;
    wire N__25713;
    wire N__25710;
    wire N__25705;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25680;
    wire N__25675;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25660;
    wire N__25659;
    wire N__25656;
    wire N__25651;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25627;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25597;
    wire N__25596;
    wire N__25593;
    wire N__25588;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25576;
    wire N__25575;
    wire N__25574;
    wire N__25573;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25566;
    wire N__25565;
    wire N__25564;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25560;
    wire N__25559;
    wire N__25558;
    wire N__25557;
    wire N__25556;
    wire N__25555;
    wire N__25554;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25498;
    wire N__25497;
    wire N__25496;
    wire N__25487;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25433;
    wire N__25430;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25409;
    wire N__25406;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25394;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25307;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25286;
    wire N__25285;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24977;
    wire N__24974;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24919;
    wire N__24914;
    wire N__24911;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24872;
    wire N__24871;
    wire N__24866;
    wire N__24863;
    wire N__24862;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24844;
    wire N__24843;
    wire N__24840;
    wire N__24835;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24774;
    wire N__24767;
    wire N__24764;
    wire N__24763;
    wire N__24762;
    wire N__24755;
    wire N__24754;
    wire N__24751;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24734;
    wire N__24731;
    wire N__24730;
    wire N__24729;
    wire N__24728;
    wire N__24727;
    wire N__24726;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24653;
    wire N__24652;
    wire N__24651;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24625;
    wire N__24620;
    wire N__24617;
    wire N__24616;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24589;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24545;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24379;
    wire N__24374;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24359;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24341;
    wire N__24338;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24296;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24288;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24263;
    wire N__24262;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24247;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24232;
    wire N__24229;
    wire N__24224;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24216;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24200;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24182;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24163;
    wire N__24160;
    wire N__24155;
    wire N__24152;
    wire N__24151;
    wire N__24150;
    wire N__24147;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24131;
    wire N__24128;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24104;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24056;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24044;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24011;
    wire N__24008;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23989;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23891;
    wire N__23890;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23831;
    wire N__23830;
    wire N__23825;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23797;
    wire N__23792;
    wire N__23789;
    wire N__23788;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23773;
    wire N__23768;
    wire N__23765;
    wire N__23764;
    wire N__23763;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23740;
    wire N__23737;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23713;
    wire N__23710;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23690;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23652;
    wire N__23651;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23593;
    wire N__23592;
    wire N__23589;
    wire N__23584;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23560;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23515;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22681;
    wire N__22680;
    wire N__22677;
    wire N__22676;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22660;
    wire N__22655;
    wire N__22652;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22647;
    wire N__22644;
    wire N__22635;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22629;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22611;
    wire N__22604;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22596;
    wire N__22591;
    wire N__22588;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22426;
    wire N__22425;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22402;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22314;
    wire N__22309;
    wire N__22306;
    wire N__22301;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22243;
    wire N__22240;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22228;
    wire N__22223;
    wire N__22220;
    wire N__22219;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22157;
    wire N__22156;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22114;
    wire N__22113;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22057;
    wire N__22054;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22018;
    wire N__22015;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21902;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21884;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21847;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21815;
    wire N__21812;
    wire N__21811;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21796;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21724;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21631;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21574;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21487;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21434;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21260;
    wire N__21257;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21225;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21170;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21085;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21031;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20990;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20969;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20922;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20887;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20694;
    wire N__20691;
    wire N__20686;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20661;
    wire N__20656;
    wire N__20651;
    wire N__20648;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20617;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20497;
    wire N__20492;
    wire N__20489;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20455;
    wire N__20454;
    wire N__20451;
    wire N__20446;
    wire N__20441;
    wire N__20440;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20393;
    wire N__20390;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20318;
    wire N__20317;
    wire N__20316;
    wire N__20315;
    wire N__20314;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20152;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20122;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20110;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20095;
    wire N__20090;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20044;
    wire N__20039;
    wire N__20036;
    wire N__20035;
    wire N__20034;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20003;
    wire N__20000;
    wire N__19999;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19978;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19942;
    wire N__19941;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19918;
    wire N__19913;
    wire N__19910;
    wire N__19909;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19885;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19840;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19798;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19480;
    wire N__19479;
    wire N__19476;
    wire N__19475;
    wire N__19474;
    wire N__19469;
    wire N__19466;
    wire N__19461;
    wire N__19458;
    wire N__19453;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19441;
    wire N__19438;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19420;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19408;
    wire N__19407;
    wire N__19406;
    wire N__19405;
    wire N__19404;
    wire N__19399;
    wire N__19394;
    wire N__19389;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19336;
    wire N__19335;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19324;
    wire N__19319;
    wire N__19314;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19304;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19296;
    wire N__19289;
    wire N__19284;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19261;
    wire N__19260;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19254;
    wire N__19249;
    wire N__19242;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19225;
    wire N__19222;
    wire N__19217;
    wire N__19212;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19180;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19105;
    wire N__19102;
    wire N__19101;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19089;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire GNDG0;
    wire VCCG0;
    wire \pid_alt.O_1_12 ;
    wire \pid_alt.O_1_15 ;
    wire \pid_alt.O_1_16 ;
    wire \pid_alt.O_1_17 ;
    wire \pid_alt.O_1_19 ;
    wire \pid_alt.O_1_20 ;
    wire \pid_alt.O_1_7 ;
    wire \pid_alt.O_1_22 ;
    wire \pid_alt.O_1_23 ;
    wire \pid_alt.O_1_18 ;
    wire \pid_alt.O_1_24 ;
    wire \pid_alt.O_1_13 ;
    wire \pid_alt.O_1_14 ;
    wire \pid_alt.O_1_10 ;
    wire \pid_alt.O_1_21 ;
    wire \pid_alt.O_2_13 ;
    wire \pid_alt.O_2_21 ;
    wire \pid_alt.O_2_18 ;
    wire \pid_alt.O_2_20 ;
    wire \pid_alt.O_2_22 ;
    wire \pid_alt.O_2_11 ;
    wire \pid_alt.O_2_24 ;
    wire \pid_alt.O_2_7 ;
    wire \pid_alt.O_2_8 ;
    wire \pid_alt.O_2_23 ;
    wire \pid_alt.O_2_10 ;
    wire \pid_alt.O_2_9 ;
    wire \pid_alt.O_2_16 ;
    wire \pid_alt.O_2_17 ;
    wire \pid_alt.O_1_6 ;
    wire \pid_alt.O_2_12 ;
    wire \pid_alt.O_2_19 ;
    wire \pid_alt.O_2_14 ;
    wire \pid_alt.O_2_15 ;
    wire \pid_alt.O_1_5 ;
    wire \pid_side.O_0_9 ;
    wire \pid_side.O_0_19 ;
    wire \pid_side.O_0_14 ;
    wire \pid_side.O_0_8 ;
    wire \pid_side.O_0_10 ;
    wire \pid_side.O_0_23 ;
    wire \pid_side.O_0_15 ;
    wire \pid_side.O_0_18 ;
    wire \pid_side.O_0_11 ;
    wire \pid_side.O_0_6 ;
    wire \pid_side.O_0_17 ;
    wire \pid_side.O_0_16 ;
    wire \pid_side.O_0_12 ;
    wire \pid_side.O_0_20 ;
    wire \pid_side.O_0_21 ;
    wire \pid_side.O_0_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ;
    wire \pid_alt.O_1_4 ;
    wire \pid_alt.O_3_4 ;
    wire \pid_alt.N_1505_i ;
    wire \pid_alt.N_1505_i_cascade_ ;
    wire \pid_alt.un1_pid_prereg_0_axb_2_1 ;
    wire \pid_alt.N_1513_0_cascade_ ;
    wire \pid_alt.N_1505_i_0 ;
    wire \pid_alt.N_3_0 ;
    wire \pid_alt.N_1507_0 ;
    wire \pid_alt.N_5 ;
    wire \pid_alt.N_1511_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_0 ;
    wire \pid_alt.N_1505_i_1 ;
    wire \pid_alt.N_1507_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_1 ;
    wire \pid_alt.error_d_regZ0Z_1 ;
    wire \pid_alt.N_3_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ;
    wire \pid_alt.error_d_regZ0Z_2 ;
    wire \pid_alt.error_d_reg_prevZ0Z_2 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ;
    wire \pid_alt.error_d_reg_prevZ0Z_3 ;
    wire \pid_alt.error_d_regZ0Z_3 ;
    wire \pid_alt.g0_4_0 ;
    wire \pid_alt.O_3_6 ;
    wire \pid_alt.error_p_regZ0Z_2 ;
    wire \pid_alt.O_3_7 ;
    wire \pid_alt.error_p_regZ0Z_3 ;
    wire \pid_alt.O_3_5 ;
    wire \pid_alt.error_p_regZ0Z_1 ;
    wire \pid_alt.O_3_12 ;
    wire \pid_alt.O_3_16 ;
    wire \pid_alt.O_3_17 ;
    wire \pid_alt.O_3_18 ;
    wire \pid_alt.O_3_24 ;
    wire \pid_alt.O_3_20 ;
    wire \pid_alt.O_3_21 ;
    wire \pid_alt.O_3_22 ;
    wire \pid_alt.O_3_23 ;
    wire \pid_alt.O_3_15 ;
    wire \pid_alt.O_3_19 ;
    wire \pid_alt.O_3_14 ;
    wire \pid_alt.O_3_8 ;
    wire \pid_alt.O_3_9 ;
    wire \pid_alt.O_3_10 ;
    wire \pid_alt.O_3_11 ;
    wire \pid_alt.O_3_13 ;
    wire \pid_alt.O_1_8 ;
    wire \pid_alt.O_1_11 ;
    wire alt_kd_6;
    wire alt_kd_2;
    wire alt_kd_7;
    wire alt_kd_5;
    wire alt_kd_1;
    wire \pid_alt.O_1_9 ;
    wire alt_ki_0;
    wire alt_ki_4;
    wire alt_ki_1;
    wire alt_ki_2;
    wire alt_ki_3;
    wire alt_ki_5;
    wire \pid_alt.O_2_5 ;
    wire \pid_alt.O_2_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ;
    wire \pid_alt.error_p_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prevZ0Z_4 ;
    wire \pid_alt.error_d_regZ0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prevZ0Z_9 ;
    wire \pid_alt.error_p_regZ0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ;
    wire \pid_alt.error_d_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_18 ;
    wire \pid_alt.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prevZ0Z_5 ;
    wire \pid_alt.error_d_regZ0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ;
    wire \pid_alt.error_p_regZ0Z_6 ;
    wire \pid_alt.error_d_reg_prevZ0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_6 ;
    wire \pid_side.O_0_24 ;
    wire \pid_side.O_0_13 ;
    wire \dron_frame_decoder_1.drone_altitude_10 ;
    wire \dron_frame_decoder_1.drone_altitude_8 ;
    wire \dron_frame_decoder_1.drone_altitude_9 ;
    wire alt_kp_2;
    wire alt_kp_3;
    wire alt_kp_5;
    wire alt_kp_6;
    wire alt_kd_3;
    wire alt_kd_0;
    wire alt_kd_4;
    wire \pid_alt.O_2_6 ;
    wire \pid_alt.N_850_0_g ;
    wire \pid_alt.error_i_acumm_preregZ0Z_6 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_10 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_9 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_8 ;
    wire bfn_3_14_0_;
    wire \pid_alt.error_i_regZ0Z_1 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_0 ;
    wire \pid_alt.error_i_regZ0Z_2 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_1 ;
    wire \pid_alt.error_i_regZ0Z_3 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_2 ;
    wire \pid_alt.error_i_regZ0Z_4 ;
    wire \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_3 ;
    wire \pid_alt.error_i_regZ0Z_5 ;
    wire \pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_4 ;
    wire \pid_alt.error_i_acummZ0Z_6 ;
    wire \pid_alt.error_i_regZ0Z_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_5 ;
    wire \pid_alt.error_i_regZ0Z_7 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7 ;
    wire \pid_alt.error_i_acummZ0Z_8 ;
    wire \pid_alt.error_i_regZ0Z_8 ;
    wire bfn_3_15_0_;
    wire \pid_alt.error_i_acummZ0Z_9 ;
    wire \pid_alt.error_i_regZ0Z_9 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_8 ;
    wire \pid_alt.error_i_acummZ0Z_10 ;
    wire \pid_alt.error_i_regZ0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9 ;
    wire \pid_alt.error_i_regZ0Z_11 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_10 ;
    wire \pid_alt.error_i_regZ0Z_12 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_11 ;
    wire \pid_alt.error_i_regZ0Z_13 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_12 ;
    wire \pid_alt.error_i_regZ0Z_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_13 ;
    wire \pid_alt.error_i_regZ0Z_15 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_14 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_15 ;
    wire \pid_alt.error_i_regZ0Z_16 ;
    wire bfn_3_16_0_;
    wire \pid_alt.error_i_regZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_16 ;
    wire \pid_alt.error_i_regZ0Z_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_17 ;
    wire \pid_alt.error_i_regZ0Z_19 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_18 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19 ;
    wire \pid_alt.error_i_regZ0Z_20 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ;
    wire \pid_alt.error_p_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prevZ0Z_17 ;
    wire \pid_alt.error_d_regZ0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ;
    wire \pid_alt.error_d_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prevZ0Z_16 ;
    wire \pid_alt.error_p_regZ0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8_cascade_ ;
    wire \Commands_frame_decoder.source_CH1data8 ;
    wire \Commands_frame_decoder.state_ns_i_a2_1_1_0 ;
    wire bfn_3_19_0_;
    wire \pid_alt.error_1 ;
    wire \pid_alt.error_cry_0 ;
    wire \pid_alt.error_2 ;
    wire \pid_alt.error_cry_1 ;
    wire \pid_alt.error_3 ;
    wire \pid_alt.error_cry_2 ;
    wire alt_command_0;
    wire \pid_alt.error_4 ;
    wire \pid_alt.error_cry_3 ;
    wire drone_altitude_i_5;
    wire alt_command_1;
    wire \pid_alt.error_5 ;
    wire \pid_alt.error_cry_4 ;
    wire drone_altitude_i_6;
    wire alt_command_2;
    wire \pid_alt.error_6 ;
    wire \pid_alt.error_cry_5 ;
    wire drone_altitude_i_7;
    wire alt_command_3;
    wire \pid_alt.error_7 ;
    wire \pid_alt.error_cry_6 ;
    wire \pid_alt.error_cry_7 ;
    wire drone_altitude_i_8;
    wire alt_command_4;
    wire \pid_alt.error_8 ;
    wire bfn_3_20_0_;
    wire drone_altitude_i_9;
    wire alt_command_5;
    wire \pid_alt.error_9 ;
    wire \pid_alt.error_cry_8 ;
    wire drone_altitude_i_10;
    wire alt_command_6;
    wire \pid_alt.error_10 ;
    wire \pid_alt.error_cry_9 ;
    wire alt_command_7;
    wire \pid_alt.error_11 ;
    wire \pid_alt.error_cry_10 ;
    wire \pid_alt.error_12 ;
    wire \pid_alt.error_cry_11 ;
    wire \pid_alt.error_13 ;
    wire \pid_alt.error_cry_12 ;
    wire \pid_alt.error_14 ;
    wire \pid_alt.error_cry_13 ;
    wire drone_altitude_15;
    wire \pid_alt.error_cry_14 ;
    wire \pid_alt.error_15 ;
    wire \dron_frame_decoder_1.drone_altitude_11 ;
    wire drone_altitude_i_11;
    wire \pid_alt.error_i_acummZ0Z_11 ;
    wire \pid_alt.error_i_acummZ0Z_7 ;
    wire alt_kp_1;
    wire alt_kp_7;
    wire \Commands_frame_decoder.state_RNIRSI31Z0Z_11 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ;
    wire \Commands_frame_decoder.state_ns_0_a3_3_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ;
    wire \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ;
    wire \pid_alt.error_p_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prevZ0Z_13 ;
    wire \pid_alt.error_d_regZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ;
    wire \pid_alt.error_p_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_14 ;
    wire \pid_alt.error_d_reg_prevZ0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ;
    wire \pid_alt.error_i_acummZ0Z_5 ;
    wire \pid_alt.N_295_cascade_ ;
    wire \pid_alt.error_i_acummZ0Z_1 ;
    wire \pid_alt.error_i_acummZ0Z_2 ;
    wire \pid_alt.error_i_acummZ0Z_3 ;
    wire \pid_alt.m39_i_a2_3 ;
    wire \pid_alt.m39_i_a2_4 ;
    wire \pid_alt.error_i_acumm7lto5 ;
    wire \pid_alt.N_294_cascade_ ;
    wire \pid_alt.N_294 ;
    wire \pid_alt.N_295 ;
    wire \pid_alt.error_i_acumm7lto4 ;
    wire \pid_alt.error_i_acummZ0Z_4 ;
    wire bfn_4_15_0_;
    wire \pid_alt.un1_pid_prereg_0 ;
    wire \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ;
    wire \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_0 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ;
    wire \pid_alt.un1_pid_prereg_0_cry_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ;
    wire \pid_alt.un1_pid_prereg_0_cry_2 ;
    wire \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_3 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ;
    wire \pid_alt.un1_pid_prereg_0_cry_4 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4 ;
    wire \pid_alt.un1_pid_prereg_0_cry_5 ;
    wire \pid_alt.un1_pid_prereg_0_cry_6 ;
    wire bfn_4_16_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ;
    wire \pid_alt.un1_pid_prereg_0_cry_9 ;
    wire \pid_alt.un1_pid_prereg_0_cry_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11 ;
    wire \pid_alt.un1_pid_prereg_0_cry_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_13 ;
    wire \pid_alt.un1_pid_prereg_0_cry_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ;
    wire bfn_4_17_0_;
    wire \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ;
    wire \pid_alt.un1_pid_prereg_0_cry_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ;
    wire \pid_alt.un1_pid_prereg_0_cry_16 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ;
    wire \pid_alt.un1_pid_prereg_0_cry_17 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ;
    wire \pid_alt.un1_pid_prereg_0_cry_18 ;
    wire \pid_alt.un1_pid_prereg_0_cry_19 ;
    wire \pid_alt.un1_pid_prereg_0_cry_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ;
    wire \pid_alt.un1_pid_prereg_0_cry_21 ;
    wire \pid_alt.un1_pid_prereg_0_cry_22 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ;
    wire bfn_4_18_0_;
    wire \pid_alt.un1_pid_prereg_0_cry_23 ;
    wire \pid_alt.error_axbZ0Z_13 ;
    wire drone_altitude_13;
    wire \pid_alt.error_axbZ0Z_14 ;
    wire drone_altitude_14;
    wire \pid_alt.error_axbZ0Z_2 ;
    wire \pid_alt.error_axbZ0Z_3 ;
    wire \pid_alt.error_d_reg_prev_i_0 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_8 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_9 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_10 ;
    wire \pid_alt.error_axbZ0Z_1 ;
    wire drone_altitude_12;
    wire \pid_alt.error_axbZ0Z_12 ;
    wire \pid_side.error_axb_0 ;
    wire bfn_4_21_0_;
    wire \pid_side.error_1 ;
    wire \pid_side.error_cry_0 ;
    wire \pid_side.error_2 ;
    wire \pid_side.error_cry_1 ;
    wire \pid_side.error_3 ;
    wire \pid_side.error_cry_2 ;
    wire \pid_side.error_4 ;
    wire \pid_side.error_cry_3 ;
    wire \pid_side.error_5 ;
    wire \pid_side.error_cry_0_0 ;
    wire \pid_side.error_6 ;
    wire \pid_side.error_cry_1_0 ;
    wire \pid_side.error_7 ;
    wire \pid_side.error_cry_2_0 ;
    wire \pid_side.error_cry_3_0 ;
    wire drone_H_disp_side_i_8;
    wire \pid_side.error_8 ;
    wire bfn_4_22_0_;
    wire drone_H_disp_side_i_9;
    wire \pid_side.error_9 ;
    wire \pid_side.error_cry_4 ;
    wire drone_H_disp_side_i_10;
    wire \pid_side.error_10 ;
    wire \pid_side.error_cry_5 ;
    wire \pid_side.error_11 ;
    wire \pid_side.error_cry_6 ;
    wire \pid_side.error_12 ;
    wire \pid_side.error_cry_7 ;
    wire \pid_side.error_13 ;
    wire \pid_side.error_cry_8 ;
    wire \pid_side.error_14 ;
    wire \pid_side.error_cry_9 ;
    wire \pid_side.error_cry_10 ;
    wire \pid_side.error_15 ;
    wire alt_kp_0;
    wire \Commands_frame_decoder.N_418 ;
    wire \Commands_frame_decoder.N_382_2 ;
    wire \Commands_frame_decoder.N_383_cascade_ ;
    wire \Commands_frame_decoder.state_ns_i_0_0_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_0 ;
    wire \Commands_frame_decoder.stateZ0Z_11 ;
    wire frame_decoder_CH4data_7;
    wire \Commands_frame_decoder.state_ns_i_a2_0_2_0 ;
    wire \Commands_frame_decoder.stateZ0Z_1 ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ;
    wire \Commands_frame_decoder.state_ns_0_a3_0_3_2 ;
    wire \Commands_frame_decoder.stateZ0Z_5 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ;
    wire \pid_alt.error_d_regZ0Z_12 ;
    wire \pid_alt.error_d_reg_prevZ0Z_12 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ;
    wire \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ;
    wire \pid_alt.error_p_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prevZ0Z_10 ;
    wire \pid_alt.error_d_regZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prevZ0Z_11 ;
    wire \pid_alt.error_p_regZ0Z_11 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ;
    wire \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_11 ;
    wire \pid_alt.error_d_regZ0Z_0 ;
    wire \pid_alt.error_d_reg_prevZ0Z_0 ;
    wire \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ;
    wire \pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12 ;
    wire \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ;
    wire \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ;
    wire \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ;
    wire \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ;
    wire \pid_alt.error_i_acumm7lto12 ;
    wire \pid_alt.error_i_acummZ0Z_12 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_3 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_1 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_7 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_2 ;
    wire \pid_alt.un1_reset_1_i_a5_0_7_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_15 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_14 ;
    wire \pid_alt.un1_reset_1_i_a5_0_9 ;
    wire \pid_alt.un1_reset_1_i_a5_0_8 ;
    wire \pid_alt.N_557_cascade_ ;
    wire \pid_alt.un1_reset_1_i_a5_0_10 ;
    wire \pid_alt.N_304_cascade_ ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prevZ0Z_8 ;
    wire \pid_alt.error_d_regZ0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ;
    wire \pid_alt.error_d_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prevZ0Z_7 ;
    wire \pid_alt.error_p_regZ0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ;
    wire \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ;
    wire \pid_alt.pid_preregZ0Z_20 ;
    wire \pid_alt.pid_preregZ0Z_19 ;
    wire \pid_alt.pid_preregZ0Z_22 ;
    wire \pid_alt.pid_preregZ0Z_17 ;
    wire \pid_alt.pid_preregZ0Z_21 ;
    wire \pid_alt.pid_preregZ0Z_15 ;
    wire \pid_alt.pid_preregZ0Z_23 ;
    wire \pid_alt.pid_preregZ0Z_18 ;
    wire \pid_alt.error_p_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ;
    wire \pid_alt.error_d_regZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_19 ;
    wire \pid_alt.error_d_reg_prevZ0Z_20 ;
    wire \pid_alt.error_p_regZ0Z_20 ;
    wire \pid_alt.error_d_regZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1_cascade_ ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ;
    wire \pid_alt.un1_pid_prereg_236_1 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ;
    wire \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_ ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ;
    wire \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ;
    wire drone_altitude_1;
    wire drone_altitude_2;
    wire drone_altitude_3;
    wire \dron_frame_decoder_1.drone_altitude_5 ;
    wire \dron_frame_decoder_1.drone_altitude_6 ;
    wire xy_kp_0;
    wire xy_kp_2;
    wire xy_kp_6;
    wire \dron_frame_decoder_1.drone_altitude_4 ;
    wire drone_altitude_i_4;
    wire \pid_alt.error_i_regZ0Z_0 ;
    wire \pid_alt.error_i_acummZ0Z_0 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_0 ;
    wire drone_H_disp_side_i_13;
    wire drone_H_disp_side_i_6;
    wire side_command_0;
    wire side_command_1;
    wire side_command_2;
    wire side_command_3;
    wire side_command_4;
    wire side_command_5;
    wire side_command_6;
    wire drone_H_disp_side_15;
    wire \Commands_frame_decoder.stateZ0Z_12 ;
    wire \Commands_frame_decoder.stateZ0Z_13 ;
    wire \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ;
    wire \Commands_frame_decoder.WDT8lto13_1_cascade_ ;
    wire \Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ;
    wire \Commands_frame_decoder.preinitZ0 ;
    wire \Commands_frame_decoder.WDT8lt14_0_cascade_ ;
    wire \Commands_frame_decoder.WDT8lt14_0 ;
    wire \Commands_frame_decoder.N_377_0 ;
    wire \Commands_frame_decoder.N_377_0_cascade_ ;
    wire \Commands_frame_decoder.N_384 ;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ;
    wire frame_decoder_OFF4data_7;
    wire \Commands_frame_decoder.source_CH4data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ;
    wire \dron_frame_decoder_1.WDT10lto13_1 ;
    wire \dron_frame_decoder_1.WDT10lt14_0_cascade_ ;
    wire \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa ;
    wire \Commands_frame_decoder.stateZ0Z_2 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ;
    wire \Commands_frame_decoder.stateZ0Z_3 ;
    wire \pid_alt.m7_e_4 ;
    wire \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_19 ;
    wire \pid_alt.un1_reset_i_a5_1_10_7_cascade_ ;
    wire \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_18 ;
    wire \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_17 ;
    wire \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_20 ;
    wire \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ;
    wire \pid_alt.error_i_acumm_preregZ0Z_16 ;
    wire \pid_alt.state_0_g_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0 ;
    wire \Commands_frame_decoder.un1_sink_data_valid_2_0_0 ;
    wire \pid_alt.pid_preregZ0Z_14 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ;
    wire \pid_alt.pid_preregZ0Z_16 ;
    wire \pid_alt.source_pid_1_sqmuxa_0_a2_2_5 ;
    wire \dron_frame_decoder_1.N_755_0 ;
    wire \dron_frame_decoder_1.drone_altitude_7 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa ;
    wire drone_H_disp_side_i_4;
    wire drone_H_disp_side_i_7;
    wire drone_H_disp_side_i_5;
    wire \pid_side.error_axbZ0Z_2 ;
    wire \pid_side.error_axbZ0Z_3 ;
    wire alt_kp_4;
    wire \Commands_frame_decoder.state_RNIF38SZ0Z_6 ;
    wire \pid_alt.state_RNIFCSD1Z0Z_0 ;
    wire \pid_alt.N_850_0 ;
    wire uart_input_drone_c;
    wire \uart_drone_sync.aux_0__0__0_0 ;
    wire \uart_drone_sync.aux_1__0__0_0 ;
    wire \Commands_frame_decoder.count_1_sqmuxa ;
    wire \Commands_frame_decoder.state_0_sqmuxa ;
    wire \Commands_frame_decoder.WDTZ0Z_0 ;
    wire bfn_8_7_0_;
    wire \Commands_frame_decoder.WDTZ0Z_1 ;
    wire \Commands_frame_decoder.un1_WDT_cry_0 ;
    wire \Commands_frame_decoder.WDTZ0Z_2 ;
    wire \Commands_frame_decoder.un1_WDT_cry_1 ;
    wire \Commands_frame_decoder.WDTZ0Z_3 ;
    wire \Commands_frame_decoder.un1_WDT_cry_2 ;
    wire \Commands_frame_decoder.WDTZ0Z_4 ;
    wire \Commands_frame_decoder.un1_WDT_cry_3 ;
    wire \Commands_frame_decoder.WDTZ0Z_5 ;
    wire \Commands_frame_decoder.un1_WDT_cry_4 ;
    wire \Commands_frame_decoder.WDTZ0Z_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_5 ;
    wire \Commands_frame_decoder.WDTZ0Z_7 ;
    wire \Commands_frame_decoder.un1_WDT_cry_6 ;
    wire \Commands_frame_decoder.un1_WDT_cry_7 ;
    wire \Commands_frame_decoder.WDTZ0Z_8 ;
    wire bfn_8_8_0_;
    wire \Commands_frame_decoder.WDTZ0Z_9 ;
    wire \Commands_frame_decoder.un1_WDT_cry_8 ;
    wire \Commands_frame_decoder.WDTZ0Z_10 ;
    wire \Commands_frame_decoder.un1_WDT_cry_9 ;
    wire \Commands_frame_decoder.WDTZ0Z_11 ;
    wire \Commands_frame_decoder.un1_WDT_cry_10 ;
    wire \Commands_frame_decoder.WDTZ0Z_12 ;
    wire \Commands_frame_decoder.un1_WDT_cry_11 ;
    wire \Commands_frame_decoder.WDTZ0Z_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_12 ;
    wire \Commands_frame_decoder.WDTZ0Z_14 ;
    wire \Commands_frame_decoder.un1_WDT_cry_13 ;
    wire \Commands_frame_decoder.un1_WDT_cry_14 ;
    wire \Commands_frame_decoder.WDTZ0Z_15 ;
    wire bfn_8_9_0_;
    wire frame_decoder_CH4data_1;
    wire frame_decoder_OFF4data_1;
    wire \scaler_4.un3_source_data_0_cry_0 ;
    wire frame_decoder_CH4data_2;
    wire frame_decoder_OFF4data_2;
    wire \scaler_4.un3_source_data_0_cry_1 ;
    wire frame_decoder_CH4data_3;
    wire frame_decoder_OFF4data_3;
    wire \scaler_4.un3_source_data_0_cry_2 ;
    wire frame_decoder_CH4data_4;
    wire frame_decoder_OFF4data_4;
    wire \scaler_4.un3_source_data_0_cry_3 ;
    wire frame_decoder_CH4data_5;
    wire frame_decoder_OFF4data_5;
    wire \scaler_4.un3_source_data_0_cry_4 ;
    wire frame_decoder_CH4data_6;
    wire frame_decoder_OFF4data_6;
    wire \scaler_4.un3_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_axb_7 ;
    wire \scaler_4.un3_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_7 ;
    wire \scaler_4.N_1684_i_l_ofxZ0 ;
    wire bfn_8_10_0_;
    wire \scaler_4.un3_source_data_0_cry_8 ;
    wire \Commands_frame_decoder.un1_state57_iZ0 ;
    wire \dron_frame_decoder_1.WDT10_0_i ;
    wire \dron_frame_decoder_1.WDTZ0Z_0 ;
    wire bfn_8_11_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_1 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_0 ;
    wire \dron_frame_decoder_1.WDTZ0Z_2 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_1 ;
    wire \dron_frame_decoder_1.WDTZ0Z_3 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_2 ;
    wire \dron_frame_decoder_1.WDTZ0Z_4 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_3 ;
    wire \dron_frame_decoder_1.WDTZ0Z_5 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_4 ;
    wire \dron_frame_decoder_1.WDTZ0Z_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_5 ;
    wire \dron_frame_decoder_1.WDTZ0Z_7 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_6 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_7 ;
    wire \dron_frame_decoder_1.WDTZ0Z_8 ;
    wire bfn_8_12_0_;
    wire \dron_frame_decoder_1.WDTZ0Z_9 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_8 ;
    wire \dron_frame_decoder_1.WDTZ0Z_10 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_9 ;
    wire \dron_frame_decoder_1.WDTZ0Z_11 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_10 ;
    wire \dron_frame_decoder_1.WDTZ0Z_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_11 ;
    wire \dron_frame_decoder_1.WDTZ0Z_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_12 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_13 ;
    wire \dron_frame_decoder_1.un1_WDT_cry_14 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ;
    wire \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ;
    wire \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ;
    wire \dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_ ;
    wire \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0 ;
    wire xy_kp_4;
    wire \Commands_frame_decoder.stateZ0Z_6 ;
    wire \Commands_frame_decoder.stateZ0Z_7 ;
    wire \Commands_frame_decoder.stateZ0Z_8 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ;
    wire \Commands_frame_decoder.stateZ0Z_9 ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa ;
    wire \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ;
    wire \Commands_frame_decoder.N_415 ;
    wire \Commands_frame_decoder.stateZ0Z_10 ;
    wire bfn_8_17_0_;
    wire \pid_side.un1_pid_prereg_cry_1 ;
    wire \pid_side.un1_pid_prereg_cry_2 ;
    wire \pid_side.un1_pid_prereg_cry_3 ;
    wire \pid_side.un1_pid_prereg_cry_4 ;
    wire \pid_side.un1_pid_prereg_cry_5 ;
    wire \pid_side.un1_pid_prereg_cry_6 ;
    wire \pid_side.un1_pid_prereg_cry_7 ;
    wire \pid_side.un1_pid_prereg_cry_8 ;
    wire bfn_8_18_0_;
    wire \pid_side.un1_pid_prereg_cry_9 ;
    wire \pid_side.un1_pid_prereg_cry_10 ;
    wire \pid_side.un1_pid_prereg_cry_11 ;
    wire \pid_side.un1_pid_prereg_cry_12 ;
    wire \pid_side.un1_pid_prereg_cry_13 ;
    wire \pid_side.un1_pid_prereg_cry_14 ;
    wire \pid_side.un1_pid_prereg_cry_15 ;
    wire \pid_side.un1_pid_prereg_cry_16 ;
    wire bfn_8_19_0_;
    wire \pid_side.un1_pid_prereg_cry_17 ;
    wire \pid_side.un1_pid_prereg_cry_18 ;
    wire \pid_side.un1_pid_prereg_cry_19 ;
    wire \pid_side.un1_pid_prereg_cry_20 ;
    wire \Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ;
    wire drone_H_disp_side_0;
    wire drone_H_disp_side_2;
    wire drone_H_disp_side_3;
    wire \dron_frame_decoder_1.drone_H_disp_side_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_5 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_6 ;
    wire \dron_frame_decoder_1.drone_H_disp_side_7 ;
    wire \dron_frame_decoder_1.N_747_0 ;
    wire alt_ki_7;
    wire uart_input_pc_c;
    wire \uart_pc_sync.aux_0__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_1__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_2__0_Z0Z_0 ;
    wire \uart_pc_sync.aux_3__0_Z0Z_0 ;
    wire \Commands_frame_decoder.stateZ0Z_14 ;
    wire \Commands_frame_decoder.countZ0Z_0 ;
    wire debug_CH3_20A_c;
    wire uart_pc_data_rdy;
    wire \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ;
    wire \Commands_frame_decoder.N_422 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2 ;
    wire \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ;
    wire \uart_pc.data_AuxZ0Z_4 ;
    wire \uart_pc.data_AuxZ1Z_0 ;
    wire \scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ;
    wire bfn_9_10_0_;
    wire \scaler_4.un2_source_data_0_cry_1 ;
    wire \scaler_4.un3_source_data_0_cry_1_c_RNI74CL ;
    wire \scaler_4.un2_source_data_0_cry_2 ;
    wire \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ;
    wire \scaler_4.un2_source_data_0_cry_3 ;
    wire \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ;
    wire \scaler_4.un2_source_data_0_cry_4 ;
    wire \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ;
    wire \scaler_4.un2_source_data_0_cry_5 ;
    wire \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ;
    wire \scaler_4.un2_source_data_0_cry_6 ;
    wire \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ;
    wire \scaler_4.un2_source_data_0_cry_7 ;
    wire \scaler_4.un2_source_data_0_cry_8 ;
    wire \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ;
    wire \scaler_4.un3_source_data_0_cry_8_c_RNIS918 ;
    wire bfn_9_11_0_;
    wire \scaler_4.un2_source_data_0_cry_9 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ;
    wire \dron_frame_decoder_1.N_412_4_cascade_ ;
    wire \dron_frame_decoder_1.WDTZ0Z_15 ;
    wire \dron_frame_decoder_1.WDTZ0Z_14 ;
    wire \dron_frame_decoder_1.WDT10lt14_0 ;
    wire \dron_frame_decoder_1.N_177_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_0 ;
    wire \dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3 ;
    wire \dron_frame_decoder_1.stateZ0Z_4 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ;
    wire \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ;
    wire \dron_frame_decoder_1.stateZ0Z_7 ;
    wire \dron_frame_decoder_1.stateZ0Z_6 ;
    wire \dron_frame_decoder_1.N_412_4 ;
    wire \dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0 ;
    wire \dron_frame_decoder_1.N_175 ;
    wire \dron_frame_decoder_1.stateZ0Z_5 ;
    wire \dron_frame_decoder_1.N_431 ;
    wire \dron_frame_decoder_1.N_435 ;
    wire \dron_frame_decoder_1.stateZ0Z_1 ;
    wire \pid_side.un1_pid_prereg_cry_8_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_9 ;
    wire \dron_frame_decoder_1.N_428 ;
    wire \dron_frame_decoder_1.stateZ0Z_3 ;
    wire \pid_side.un1_pid_prereg_cry_7_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_8 ;
    wire \pid_side.error_p_regZ0Z_11 ;
    wire \pid_side.un1_pid_prereg_cry_10_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_3_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_4 ;
    wire \pid_side.error_p_regZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_cry_5_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_18_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_19 ;
    wire \pid_side.error_p_regZ0Z_15 ;
    wire \pid_side.un1_pid_prereg_cry_14_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_14 ;
    wire \pid_side.un1_pid_prereg_cry_13_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_16_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_17 ;
    wire \pid_side.un1_pid_prereg_cry_19_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_20 ;
    wire \pid_side.error_p_regZ0Z_12 ;
    wire \pid_side.un1_pid_prereg_cry_11_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_17_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_18 ;
    wire \pid_alt.error_d_reg_prevZ0Z_15 ;
    wire \pid_alt.error_p_regZ0Z_15 ;
    wire \pid_alt.error_d_regZ0Z_15 ;
    wire \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ;
    wire \pid_side.error_axb_8_l_ofxZ0 ;
    wire side_command_7;
    wire \pid_side.error_axbZ0Z_7 ;
    wire drone_H_disp_front_2;
    wire drone_H_disp_side_1;
    wire \pid_side.error_axbZ0Z_1 ;
    wire \pid_alt.state_1_0_0 ;
    wire \uart_pc.state_srsts_0_0_0_cascade_ ;
    wire \uart_pc.N_143_cascade_ ;
    wire \uart_pc.data_rdyc_1 ;
    wire \uart_pc.data_rdyc_1_cascade_ ;
    wire \uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ;
    wire \uart_drone.stateZ0Z_1 ;
    wire \uart_drone.state_srsts_i_0_2_cascade_ ;
    wire \scaler_4.un2_source_data_0 ;
    wire frame_decoder_OFF4data_0;
    wire frame_decoder_CH4data_0;
    wire \scaler_4.debug_CH3_20A_c_0 ;
    wire \uart_pc.data_AuxZ1Z_2 ;
    wire \uart_pc.data_AuxZ1Z_1 ;
    wire \uart_pc.data_Auxce_0_3 ;
    wire \uart_pc.data_AuxZ0Z_3 ;
    wire \uart_pc.data_AuxZ0Z_5 ;
    wire \uart_pc.data_Auxce_0_0_4 ;
    wire \uart_pc.data_Auxce_0_5 ;
    wire \uart_pc.data_Auxce_0_0_2 ;
    wire \uart_drone.data_rdyc_1_0 ;
    wire \uart_drone.timer_Count_RNIES9Q1Z0Z_2 ;
    wire \dron_frame_decoder_1.stateZ0Z_2 ;
    wire uart_drone_data_rdy;
    wire \pid_alt.pid_preregZ0Z_10 ;
    wire \pid_alt.un1_reset_i_a2_3_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_8 ;
    wire \pid_alt.un1_reset_i_a5_1_10_5_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_6 ;
    wire \pid_side.un1_pid_prereg_cry_9_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_10 ;
    wire \pid_side.un1_reset_i_a2_3_cascade_ ;
    wire \pid_side.pid_preregZ0Z_18 ;
    wire \pid_side.pid_preregZ0Z_17 ;
    wire \pid_side.pid_preregZ0Z_19 ;
    wire \pid_side.pid_preregZ0Z_20 ;
    wire \dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ;
    wire drone_H_disp_side_11;
    wire drone_H_disp_side_13;
    wire drone_H_disp_side_14;
    wire \dron_frame_decoder_1.N_739_0 ;
    wire drone_H_disp_side_12;
    wire drone_H_disp_side_i_12;
    wire drone_H_disp_front_3;
    wire xy_kp_3;
    wire \uart_drone_sync.aux_2__0__0_0 ;
    wire bfn_11_7_0_;
    wire \uart_pc.timer_Count_RNO_0Z0Z_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_1 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_3 ;
    wire \uart_pc.un4_timer_Count_1_cry_2 ;
    wire \uart_pc.un4_timer_Count_1_cry_3 ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_4 ;
    wire \uart_pc.un1_state_2_0_a3_0 ;
    wire \uart_pc.timer_CountZ0Z_0 ;
    wire \uart_pc.timer_Count_0_sqmuxa ;
    wire \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_1 ;
    wire \uart_drone.data_rdyc_1 ;
    wire \uart_drone_sync.aux_3__0__0_0 ;
    wire \uart_drone.timer_Count_0_sqmuxa_cascade_ ;
    wire \uart_pc.N_145_cascade_ ;
    wire \uart_pc.N_144_1 ;
    wire \uart_pc.N_144_1_cascade_ ;
    wire \uart_pc.N_143 ;
    wire \uart_pc.stateZ0Z_4 ;
    wire \uart_pc.N_152_cascade_ ;
    wire \uart_pc.stateZ0Z_3 ;
    wire \uart_pc.CO0_cascade_ ;
    wire \uart_pc.un1_state_4_0 ;
    wire \uart_pc.un1_state_7_0 ;
    wire \uart_pc.data_Auxce_0_0_0 ;
    wire \uart_pc.bit_CountZ0Z_1 ;
    wire \uart_pc.bit_CountZ0Z_2 ;
    wire \uart_pc.bit_CountZ0Z_0 ;
    wire \uart_pc.data_Auxce_0_1 ;
    wire \uart_drone.data_AuxZ0Z_0 ;
    wire \uart_drone.data_AuxZ0Z_1 ;
    wire \uart_drone.data_AuxZ0Z_2 ;
    wire \uart_drone.data_AuxZ0Z_3 ;
    wire \uart_drone.data_AuxZ0Z_4 ;
    wire \uart_drone.data_AuxZ0Z_5 ;
    wire \uart_drone.data_AuxZ0Z_6 ;
    wire \uart_drone.data_AuxZ0Z_7 ;
    wire \pid_alt.pid_preregZ0Z_9 ;
    wire \uart_drone.data_Auxce_0_0_0 ;
    wire \uart_drone.data_Auxce_0_1 ;
    wire \uart_drone.data_Auxce_0_3 ;
    wire \uart_drone.data_Auxce_0_0_4 ;
    wire \pid_alt.un1_reset_i_a5_0_6_3 ;
    wire \pid_alt.N_306_5 ;
    wire \pid_alt.un1_reset_i_a5_0_6_2_cascade_ ;
    wire \pid_alt.un1_reset_i_a5_1_10_8 ;
    wire \pid_alt.un1_reset_i_a5_1_10_9 ;
    wire \pid_alt.un1_reset_i_a5_0_6_cascade_ ;
    wire \pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_ ;
    wire \uart_drone.data_Auxce_0_5 ;
    wire \pid_alt.N_530 ;
    wire \pid_alt.N_535 ;
    wire \pid_alt.pid_preregZ0Z_5 ;
    wire \pid_alt.N_535_cascade_ ;
    wire \pid_alt.pid_preregZ0Z_4 ;
    wire \uart_drone.data_Auxce_0_6 ;
    wire \pid_alt.pid_preregZ0Z_12 ;
    wire \pid_alt.pid_preregZ0Z_13 ;
    wire \pid_alt.pid_preregZ0Z_24 ;
    wire \pid_alt.N_551 ;
    wire \pid_side.un1_pid_prereg_cry_6_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_7 ;
    wire \pid_side.un1_pid_prereg_cry_2_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_16 ;
    wire \pid_side.un1_pid_prereg_cry_15_THRU_CO ;
    wire \pid_side.un1_pid_prereg_cry_4_THRU_CO ;
    wire \pid_side.error_p_regZ0Z_5 ;
    wire \pid_side.error_p_regZ0Z_13 ;
    wire \pid_side.un1_pid_prereg_cry_12_THRU_CO ;
    wire xy_kp_1;
    wire xy_kp_7;
    wire \pid_alt.stateZ0Z_0 ;
    wire \pid_alt.state_0_0 ;
    wire \uart_pc.timer_CountZ0Z_4 ;
    wire debug_CH0_16A_c;
    wire \uart_drone.state_srsts_0_0_0_cascade_ ;
    wire \uart_drone.stateZ0Z_0 ;
    wire \uart_drone.timer_Count_RNO_0_0_1_cascade_ ;
    wire \uart_pc.timer_CountZ1Z_2 ;
    wire \uart_pc.timer_CountZ1Z_3 ;
    wire \uart_pc.N_126_li ;
    wire \uart_drone.un1_state_2_0 ;
    wire scaler_4_data_6;
    wire bfn_12_10_0_;
    wire \ppm_encoder_1.un1_rudder_cry_6 ;
    wire \ppm_encoder_1.un1_rudder_cry_7 ;
    wire \ppm_encoder_1.un1_rudder_cry_8 ;
    wire \ppm_encoder_1.un1_rudder_cry_9 ;
    wire \ppm_encoder_1.un1_rudder_cry_10 ;
    wire \ppm_encoder_1.un1_rudder_cry_11 ;
    wire \ppm_encoder_1.un1_rudder_cry_12 ;
    wire \ppm_encoder_1.un1_rudder_cry_13 ;
    wire scaler_4_data_14;
    wire bfn_12_11_0_;
    wire bfn_12_12_0_;
    wire \ppm_encoder_1.un1_throttle_cry_0 ;
    wire \ppm_encoder_1.un1_throttle_cry_1 ;
    wire \ppm_encoder_1.un1_throttle_cry_2 ;
    wire \ppm_encoder_1.un1_throttle_cry_3 ;
    wire \ppm_encoder_1.un1_throttle_cry_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_5 ;
    wire \ppm_encoder_1.un1_throttle_cry_6 ;
    wire \ppm_encoder_1.un1_throttle_cry_7 ;
    wire bfn_12_13_0_;
    wire throttle_order_9;
    wire \ppm_encoder_1.un1_throttle_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_8 ;
    wire \ppm_encoder_1.un1_throttle_cry_9 ;
    wire \ppm_encoder_1.un1_throttle_cry_10 ;
    wire \ppm_encoder_1.un1_throttle_cry_11 ;
    wire \ppm_encoder_1.un1_throttle_cry_12 ;
    wire \ppm_encoder_1.un1_throttle_cry_13 ;
    wire \pid_alt.N_72_i_1 ;
    wire \uart_drone.data_Auxce_0_0_2 ;
    wire \pid_alt.pid_preregZ0Z_0 ;
    wire \pid_alt.pid_preregZ0Z_1 ;
    wire \pid_alt.pid_preregZ0Z_2 ;
    wire \pid_alt.pid_preregZ0Z_3 ;
    wire \pid_alt.N_472_1 ;
    wire \pid_alt.pid_preregZ0Z_11 ;
    wire \pid_alt.N_72_i ;
    wire \pid_alt.N_299 ;
    wire \pid_alt.pid_preregZ0Z_7 ;
    wire \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ;
    wire \ppm_encoder_1.N_292 ;
    wire \uart_drone.un1_state_7_0_cascade_ ;
    wire \uart_drone.N_152_cascade_ ;
    wire \uart_drone.bit_CountZ0Z_1 ;
    wire \uart_drone.un1_state_7_0 ;
    wire \uart_drone.bit_CountZ0Z_2 ;
    wire \uart_drone.N_152 ;
    wire \pid_front.N_533_cascade_ ;
    wire \pid_front.N_10_1 ;
    wire \pid_front.un1_reset_i_a5_0_2_cascade_ ;
    wire \pid_front.un1_reset_i_a5_0_3 ;
    wire \pid_front.pid_preregZ0Z_1 ;
    wire \uart_pc.stateZ0Z_2 ;
    wire \uart_pc.state_srsts_i_0_2 ;
    wire \uart_pc.stateZ0Z_0 ;
    wire \uart_pc.stateZ0Z_1 ;
    wire \uart_drone.timer_CountZ1Z_1 ;
    wire \uart_drone.un1_state_2_0_a3_0 ;
    wire bfn_13_8_0_;
    wire \uart_drone.timer_CountZ1Z_2 ;
    wire \uart_drone.timer_Count_RNO_0_0_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_1 ;
    wire \uart_drone.timer_Count_RNO_0_0_3 ;
    wire \uart_drone.un4_timer_Count_1_cry_2 ;
    wire \uart_drone.un4_timer_Count_1_cry_3 ;
    wire \uart_drone.timer_Count_RNO_0_0_4 ;
    wire \uart_drone.timer_Count_0_sqmuxa ;
    wire \uart_drone.timer_CountZ0Z_0 ;
    wire \uart_drone.N_126_li ;
    wire \uart_drone.N_143 ;
    wire scaler_4_data_12;
    wire \ppm_encoder_1.un1_rudder_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_rudder_cry_7_THRU_CO ;
    wire scaler_4_data_8;
    wire \ppm_encoder_1.un1_rudder_cry_6_THRU_CO ;
    wire scaler_4_data_7;
    wire scaler_4_data_11;
    wire \ppm_encoder_1.un1_rudder_cry_10_THRU_CO ;
    wire throttle_order_11;
    wire \ppm_encoder_1.un1_throttle_cry_10_THRU_CO ;
    wire scaler_4_data_13;
    wire \ppm_encoder_1.un1_rudder_cry_12_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_1_THRU_CO ;
    wire throttle_order_2;
    wire ppm_output_c;
    wire \ppm_encoder_1.un1_throttle_cry_9_THRU_CO ;
    wire throttle_order_10;
    wire \ppm_encoder_1.un1_throttle_cry_11_THRU_CO ;
    wire throttle_order_12;
    wire \ppm_encoder_1.un1_throttle_cry_2_THRU_CO ;
    wire throttle_order_3;
    wire \ppm_encoder_1.un1_throttle_cry_4_THRU_CO ;
    wire throttle_order_5;
    wire \ppm_encoder_1.un1_throttle_cry_5_THRU_CO ;
    wire throttle_order_6;
    wire \ppm_encoder_1.N_314_cascade_ ;
    wire \ppm_encoder_1.N_288_cascade_ ;
    wire \pid_alt.error_i_acumm_preregZ0Z_21 ;
    wire \pid_alt.N_557 ;
    wire \pid_alt.error_i_acumm7lto13 ;
    wire \pid_alt.error_i_acummZ0Z_13 ;
    wire \pid_alt.N_72_i_0 ;
    wire \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ;
    wire \uart_drone.stateZ0Z_4 ;
    wire \uart_drone.state_RNIOU0NZ0Z_4 ;
    wire \ppm_encoder_1.N_291 ;
    wire \uart_drone.timer_CountZ0Z_4 ;
    wire \uart_drone.timer_CountZ1Z_3 ;
    wire \uart_drone.stateZ0Z_2 ;
    wire \uart_drone.N_144_1 ;
    wire \uart_drone.N_145_cascade_ ;
    wire \uart_drone.stateZ0Z_3 ;
    wire debug_CH1_0A_c;
    wire \pid_side.state_ns_0_cascade_ ;
    wire \dron_frame_decoder_1.N_763_0 ;
    wire \pid_front.un1_reset_i_a5_0_5 ;
    wire \pid_front.un1_reset_i_1_cascade_ ;
    wire \pid_front.N_532 ;
    wire \pid_front.un1_reset_i_a2_3 ;
    wire \pid_front.stateZ0Z_1 ;
    wire \pid_front.N_287 ;
    wire \pid_front.N_533 ;
    wire \pid_front.state_0_1 ;
    wire \pid_front.pid_prereg_RNI2A6A6Z0Z_2 ;
    wire \pid_front.un1_reset_i_a5_1_6 ;
    wire \pid_front.N_315 ;
    wire drone_H_disp_front_1;
    wire \pid_front.un1_reset_i_a5_1_5_cascade_ ;
    wire \pid_front.un1_reset_i_a5_1_8 ;
    wire \pid_front.pid_preregZ0Z_10 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_8 ;
    wire \reset_module_System.reset6_15_cascade_ ;
    wire \reset_module_System.count_1_1 ;
    wire bfn_14_7_0_;
    wire \reset_module_System.count_1_cry_1 ;
    wire \reset_module_System.countZ0Z_3 ;
    wire \reset_module_System.count_1_cry_2 ;
    wire \reset_module_System.count_1_cry_3 ;
    wire \reset_module_System.count_1_cry_4 ;
    wire \reset_module_System.countZ0Z_6 ;
    wire \reset_module_System.count_1_cry_5 ;
    wire \reset_module_System.count_1_cry_6 ;
    wire \reset_module_System.count_1_cry_7 ;
    wire \reset_module_System.count_1_cry_8 ;
    wire bfn_14_8_0_;
    wire \reset_module_System.countZ0Z_10 ;
    wire \reset_module_System.count_1_cry_9 ;
    wire \reset_module_System.countZ0Z_11 ;
    wire \reset_module_System.count_1_cry_10 ;
    wire \reset_module_System.count_1_cry_11 ;
    wire \reset_module_System.count_1_cry_12 ;
    wire \reset_module_System.countZ0Z_14 ;
    wire \reset_module_System.count_1_cry_13 ;
    wire \reset_module_System.count_1_cry_14 ;
    wire \reset_module_System.count_1_cry_15 ;
    wire \reset_module_System.count_1_cry_16 ;
    wire \reset_module_System.countZ0Z_17 ;
    wire bfn_14_9_0_;
    wire \reset_module_System.count_1_cry_17 ;
    wire \reset_module_System.count_1_cry_18 ;
    wire \reset_module_System.countZ0Z_20 ;
    wire \reset_module_System.count_1_cry_19 ;
    wire \reset_module_System.count_1_cry_20 ;
    wire \reset_module_System.countZ0Z_19 ;
    wire \reset_module_System.countZ0Z_15 ;
    wire \reset_module_System.countZ0Z_21 ;
    wire \reset_module_System.countZ0Z_13 ;
    wire scaler_4_data_10;
    wire \ppm_encoder_1.un1_rudder_cry_9_THRU_CO ;
    wire \ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_11 ;
    wire \ppm_encoder_1.throttleZ0Z_11 ;
    wire \ppm_encoder_1.N_297_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_11 ;
    wire \ppm_encoder_1.elevatorZ0Z_11 ;
    wire \ppm_encoder_1.rudderZ0Z_12 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_1_12 ;
    wire \ppm_encoder_1.throttleZ0Z_12 ;
    wire \ppm_encoder_1.N_298_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_12 ;
    wire \ppm_encoder_1.elevatorZ0Z_12 ;
    wire bfn_14_14_0_;
    wire \ppm_encoder_1.un1_aileron_cry_0 ;
    wire \ppm_encoder_1.un1_aileron_cry_1 ;
    wire \ppm_encoder_1.un1_aileron_cry_2 ;
    wire \ppm_encoder_1.un1_aileron_cry_3 ;
    wire \ppm_encoder_1.un1_aileron_cry_4 ;
    wire \ppm_encoder_1.un1_aileron_cry_5 ;
    wire \ppm_encoder_1.un1_aileron_cry_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_7 ;
    wire bfn_14_15_0_;
    wire \ppm_encoder_1.un1_aileron_cry_8 ;
    wire \ppm_encoder_1.un1_aileron_cry_9 ;
    wire \ppm_encoder_1.un1_aileron_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_10 ;
    wire \ppm_encoder_1.un1_aileron_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_aileron_cry_11 ;
    wire \ppm_encoder_1.un1_aileron_cry_12 ;
    wire \ppm_encoder_1.un1_aileron_cry_13 ;
    wire drone_altitude_0;
    wire \pid_alt.drone_altitude_i_0 ;
    wire \pid_side.pid_preregZ0Z_10 ;
    wire side_order_11;
    wire \pid_side.pid_preregZ0Z_6 ;
    wire \pid_side.pid_preregZ0Z_8 ;
    wire \pid_side.pid_preregZ0Z_9 ;
    wire \uart_drone.bit_CountZ0Z_0 ;
    wire \uart_drone.un1_state_4_0 ;
    wire \uart_drone.CO0 ;
    wire \pid_side.pid_preregZ0Z_11 ;
    wire \pid_side.pid_preregZ0Z_7 ;
    wire \pid_side.un1_reset_i_a5_1_5 ;
    wire \pid_side.pid_preregZ0Z_15 ;
    wire \pid_side.pid_preregZ0Z_14 ;
    wire \pid_side.m7_e_4 ;
    wire \pid_side.pid_preregZ0Z_16 ;
    wire \pid_side.un1_reset_i_a5_1_7 ;
    wire \pid_side.N_563_cascade_ ;
    wire \pid_side.un1_reset_i_a5_1_8 ;
    wire \pid_side.N_311_cascade_ ;
    wire \pid_side.un1_reset_i_a5_1_6 ;
    wire \pid_side.error_p_regZ0Z_2 ;
    wire \pid_side.un1_pid_prereg_cry_1_THRU_CO ;
    wire \pid_side.un1_reset_i_a5_0_2 ;
    wire \pid_side.un1_reset_i_a5_0_3 ;
    wire \pid_front.N_569 ;
    wire \pid_front.pid_preregZ0Z_14 ;
    wire \pid_front.m7_e_4 ;
    wire \pid_front.pid_preregZ0Z_18 ;
    wire \pid_front.pid_preregZ0Z_19 ;
    wire \pid_front.pid_preregZ0Z_9 ;
    wire \pid_front.pid_preregZ0Z_11 ;
    wire \pid_front.pid_preregZ0Z_13 ;
    wire \reset_module_System.count_1_2 ;
    wire \reset_module_System.countZ0Z_2 ;
    wire \reset_module_System.reset6_15 ;
    wire \reset_module_System.reset6_14 ;
    wire \reset_module_System.countZ0Z_8 ;
    wire \reset_module_System.countZ0Z_7 ;
    wire \reset_module_System.countZ0Z_9 ;
    wire \reset_module_System.countZ0Z_5 ;
    wire \reset_module_System.countZ0Z_4 ;
    wire \reset_module_System.countZ0Z_1 ;
    wire \reset_module_System.countZ0Z_18 ;
    wire \reset_module_System.countZ0Z_16 ;
    wire \reset_module_System.reset6_3_cascade_ ;
    wire \reset_module_System.reset6_13 ;
    wire \reset_module_System.countZ0Z_12 ;
    wire \reset_module_System.countZ0Z_0 ;
    wire \reset_module_System.reset6_17_cascade_ ;
    wire \reset_module_System.reset6_11 ;
    wire \reset_module_System.reset6_19 ;
    wire \ppm_encoder_1.un1_rudder_cry_8_THRU_CO ;
    wire scaler_4_data_9;
    wire \ppm_encoder_1.init_pulsesZ0Z_11 ;
    wire \ppm_encoder_1.rudderZ0Z_11 ;
    wire \ppm_encoder_1.N_313_cascade_ ;
    wire bfn_15_11_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_10_7 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_10_8 ;
    wire bfn_15_12_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_11 ;
    wire \ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ;
    wire \ppm_encoder_1.un1_init_pulses_10_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_10 ;
    wire \ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_10_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_16 ;
    wire bfn_15_13_0_;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_17 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_0_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_10_18 ;
    wire \ppm_encoder_1.un1_init_pulses_0_12 ;
    wire \ppm_encoder_1.N_287 ;
    wire \ppm_encoder_1.un1_aileron_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_throttle_cry_0_THRU_CO ;
    wire throttle_order_1;
    wire \ppm_encoder_1.un1_aileron_cry_1_THRU_CO ;
    wire \ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ;
    wire \ppm_encoder_1.elevatorZ0Z_9 ;
    wire \ppm_encoder_1.N_295 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ;
    wire \ppm_encoder_1.rudderZ0Z_9 ;
    wire \ppm_encoder_1.throttleZ0Z_9 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_9 ;
    wire \ppm_encoder_1.throttleZ0Z_10 ;
    wire \ppm_encoder_1.un1_init_pulses_0_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ;
    wire \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_10 ;
    wire \ppm_encoder_1.N_296 ;
    wire \ppm_encoder_1.un1_aileron_cry_9_THRU_CO ;
    wire side_order_10;
    wire \ppm_encoder_1.aileronZ0Z_10 ;
    wire \pid_side.N_531 ;
    wire \pid_side.un1_reset_i_a5_0_5 ;
    wire \pid_side.un1_reset_i_1 ;
    wire side_order_1;
    wire \pid_side.pid_preregZ0Z_2 ;
    wire side_order_2;
    wire \pid_side.stateZ0Z_1 ;
    wire \pid_side.pid_preregZ0Z_3 ;
    wire \pid_side.N_291_cascade_ ;
    wire \pid_side.N_451_1 ;
    wire front_order_0;
    wire bfn_15_18_0_;
    wire front_order_1;
    wire \ppm_encoder_1.un1_elevator_cry_0_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_0 ;
    wire \ppm_encoder_1.un1_elevator_cry_1 ;
    wire front_order_3;
    wire \ppm_encoder_1.un1_elevator_cry_2_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_2 ;
    wire \ppm_encoder_1.un1_elevator_cry_3 ;
    wire \ppm_encoder_1.un1_elevator_cry_4 ;
    wire \ppm_encoder_1.un1_elevator_cry_5 ;
    wire \ppm_encoder_1.un1_elevator_cry_6 ;
    wire \ppm_encoder_1.un1_elevator_cry_7 ;
    wire bfn_15_19_0_;
    wire front_order_9;
    wire \ppm_encoder_1.un1_elevator_cry_8_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_8 ;
    wire \ppm_encoder_1.un1_elevator_cry_9 ;
    wire front_order_11;
    wire \ppm_encoder_1.un1_elevator_cry_10_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_10 ;
    wire front_order_12;
    wire \ppm_encoder_1.un1_elevator_cry_11_THRU_CO ;
    wire \ppm_encoder_1.un1_elevator_cry_11 ;
    wire \ppm_encoder_1.un1_elevator_cry_12 ;
    wire \ppm_encoder_1.un1_elevator_cry_13 ;
    wire \pid_front.pid_preregZ0Z_0 ;
    wire \pid_front.un1_reset_i_a5_1_7 ;
    wire uart_drone_data_7;
    wire \pid_front.pid_preregZ0Z_17 ;
    wire \pid_front.pid_preregZ0Z_20 ;
    wire \pid_front.pid_preregZ0Z_7 ;
    wire \pid_front.pid_preregZ0Z_6 ;
    wire \pid_front.pid_preregZ0Z_12 ;
    wire \pid_front.pid_preregZ0Z_16 ;
    wire \pid_front.pid_preregZ0Z_2 ;
    wire \pid_front.pid_preregZ0Z_15 ;
    wire uart_drone_data_2;
    wire uart_drone_data_3;
    wire uart_drone_data_4;
    wire uart_drone_data_5;
    wire uart_drone_data_1;
    wire scaler_4_data_4;
    wire scaler_4_data_5;
    wire \ppm_encoder_1.pid_altitude_dv_0 ;
    wire bfn_16_8_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_2 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_5 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_7 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_6 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_7 ;
    wire \ppm_encoder_1.un1_init_pulses_11_8 ;
    wire bfn_16_9_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_9 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_11 ;
    wire \ppm_encoder_1.un1_init_pulses_11_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_10 ;
    wire \ppm_encoder_1.un1_init_pulses_11_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_11 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_13 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_15 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_16 ;
    wire \ppm_encoder_1.un1_init_pulses_11_16 ;
    wire bfn_16_10_0_;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_17 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_16 ;
    wire \ppm_encoder_1.un1_init_pulses_3_cry_17 ;
    wire \ppm_encoder_1.un1_init_pulses_11_18 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_9 ;
    wire \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ;
    wire \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_13 ;
    wire \ppm_encoder_1.un1_init_pulses_10_13 ;
    wire \ppm_encoder_1.un1_init_pulses_11_14 ;
    wire \ppm_encoder_1.un1_init_pulses_10_14 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_14 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_11_15 ;
    wire \ppm_encoder_1.un1_init_pulses_10_15 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_11_1 ;
    wire \ppm_encoder_1.un1_init_pulses_10_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_10 ;
    wire \ppm_encoder_1.un1_init_pulses_10_10 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_10 ;
    wire \ppm_encoder_1.rudderZ0Z_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_8 ;
    wire \ppm_encoder_1.N_294_cascade_ ;
    wire side_order_8;
    wire \ppm_encoder_1.un1_aileron_cry_7_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_8 ;
    wire front_order_8;
    wire \ppm_encoder_1.un1_elevator_cry_7_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_8 ;
    wire throttle_order_8;
    wire \ppm_encoder_1.un1_throttle_cry_7_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_8 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ;
    wire \ppm_encoder_1.throttleZ0Z_2 ;
    wire \ppm_encoder_1.aileronZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0_2 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ;
    wire \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ;
    wire \ppm_encoder_1.aileronZ0Z_1 ;
    wire \ppm_encoder_1.elevatorZ0Z_1 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0_1 ;
    wire \ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ;
    wire \ppm_encoder_1.throttleZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ;
    wire \ppm_encoder_1.throttle_m_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ;
    wire \pid_side.pid_preregZ0Z_12 ;
    wire side_order_12;
    wire \pid_side.N_563 ;
    wire \pid_side.pid_preregZ0Z_21 ;
    wire \pid_side.pid_preregZ0Z_13 ;
    wire \pid_side.pid_preregZ0Z_4 ;
    wire \pid_side.N_534 ;
    wire \pid_side.N_291 ;
    wire \pid_side.pid_preregZ0Z_5 ;
    wire \pid_side.state_0_1 ;
    wire \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ;
    wire \ppm_encoder_1.throttleZ0Z_5 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_5 ;
    wire \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ;
    wire \ppm_encoder_1.throttleZ0Z_6 ;
    wire \ppm_encoder_1.rudderZ0Z_6 ;
    wire \ppm_encoder_1.un1_init_pulses_0_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ;
    wire \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_6 ;
    wire side_order_6;
    wire \ppm_encoder_1.un1_aileron_cry_5_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_6 ;
    wire \ppm_encoder_1.un1_aileron_cry_2_THRU_CO ;
    wire side_order_3;
    wire \ppm_encoder_1.un1_aileron_cry_4_THRU_CO ;
    wire side_order_5;
    wire \ppm_encoder_1.aileronZ0Z_5 ;
    wire side_order_9;
    wire \ppm_encoder_1.un1_aileron_cry_8_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_9 ;
    wire front_order_10;
    wire \ppm_encoder_1.un1_elevator_cry_9_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_10 ;
    wire front_order_2;
    wire \ppm_encoder_1.un1_elevator_cry_1_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_2 ;
    wire \ppm_encoder_1.un1_elevator_cry_5_THRU_CO ;
    wire front_order_6;
    wire \ppm_encoder_1.elevatorZ0Z_6 ;
    wire front_order_5;
    wire \ppm_encoder_1.un1_elevator_cry_4_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_5 ;
    wire xy_kp_5;
    wire \Commands_frame_decoder.state_RNIG48SZ0Z_7 ;
    wire \pid_front.pid_preregZ0Z_4 ;
    wire \pid_front.pid_preregZ0Z_5 ;
    wire \pid_front.pid_preregZ0Z_3 ;
    wire alt_ki_6;
    wire \Commands_frame_decoder.state_RNIQRI31Z0Z_10 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_4 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_5 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_6 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_7 ;
    wire uart_pc_data_0;
    wire uart_pc_data_1;
    wire uart_pc_data_2;
    wire uart_pc_data_3;
    wire uart_pc_data_4;
    wire uart_pc_data_5;
    wire uart_pc_data_6;
    wire uart_pc_data_7;
    wire \Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_10 ;
    wire \dron_frame_decoder_1.drone_H_disp_front_9 ;
    wire front_command_7;
    wire drone_H_disp_front_11;
    wire \uart_pc.data_Auxce_0_6 ;
    wire \uart_pc.data_AuxZ0Z_6 ;
    wire \uart_pc.un1_state_2_0 ;
    wire debug_CH2_18A_c;
    wire \uart_pc.N_152 ;
    wire \uart_pc.data_AuxZ0Z_7 ;
    wire \uart_pc.state_RNIEAGSZ0Z_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_13 ;
    wire \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ;
    wire \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_6 ;
    wire \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_12 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_12 ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_18 ;
    wire \ppm_encoder_1.un1_init_pulses_11_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_3 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_3 ;
    wire \ppm_encoder_1.un1_init_pulses_10_4 ;
    wire \ppm_encoder_1.un1_init_pulses_11_4 ;
    wire \ppm_encoder_1.un1_init_pulses_0_4 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_4 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_4 ;
    wire \ppm_encoder_1.rudderZ0Z_4 ;
    wire \ppm_encoder_1.un1_init_pulses_10_5 ;
    wire \ppm_encoder_1.un1_init_pulses_11_5 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_1 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ;
    wire \ppm_encoder_1.init_pulsesZ0Z_2 ;
    wire \ppm_encoder_1.un1_init_pulses_0Z0Z_1 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_0 ;
    wire \ppm_encoder_1.un1_init_pulses_11_0 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_6 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_10_mux ;
    wire \ppm_encoder_1.init_pulsesZ0Z_10 ;
    wire \ppm_encoder_1.rudderZ0Z_10 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ;
    wire \ppm_encoder_1.rudderZ0Z_13 ;
    wire \ppm_encoder_1.un1_init_pulses_0_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_13 ;
    wire \ppm_encoder_1.N_299_cascade_ ;
    wire side_order_13;
    wire \ppm_encoder_1.un1_aileron_cry_12_THRU_CO ;
    wire \ppm_encoder_1.aileronZ0Z_13 ;
    wire front_order_13;
    wire \ppm_encoder_1.un1_elevator_cry_12_THRU_CO ;
    wire \ppm_encoder_1.elevatorZ0Z_13 ;
    wire throttle_order_13;
    wire \ppm_encoder_1.un1_throttle_cry_12_THRU_CO ;
    wire \ppm_encoder_1.throttleZ0Z_13 ;
    wire \ppm_encoder_1.rudderZ0Z_14 ;
    wire \ppm_encoder_1.un1_init_pulses_0_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ;
    wire \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_14 ;
    wire \ppm_encoder_1.throttleZ0Z_14 ;
    wire \ppm_encoder_1.elevatorZ0Z_14 ;
    wire \ppm_encoder_1.N_300_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_14 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ;
    wire \ppm_encoder_1.pulses2countZ0Z_14 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ;
    wire \ppm_encoder_1.un1_init_pulses_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_0 ;
    wire \ppm_encoder_1.throttleZ0Z_3 ;
    wire \ppm_encoder_1.un1_init_pulses_0_3 ;
    wire \ppm_encoder_1.elevatorZ0Z_3 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ;
    wire \ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ;
    wire \pid_side.pid_preregZ0Z_0 ;
    wire \pid_side.state_0_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ;
    wire \ppm_encoder_1.PPM_STATE_53_d_cascade_ ;
    wire \ppm_encoder_1.N_134_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ;
    wire \ppm_encoder_1.N_221 ;
    wire \ppm_encoder_1.N_232_cascade_ ;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ;
    wire \ppm_encoder_1.N_139 ;
    wire \ppm_encoder_1.N_232 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_1 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ;
    wire \ppm_encoder_1.PPM_STATEZ0Z_0 ;
    wire \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ;
    wire \ppm_encoder_1.pulses2countZ0Z_2 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ;
    wire \ppm_encoder_1.pulses2countZ0Z_3 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_0 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ;
    wire \ppm_encoder_1.pulses2countZ0Z_1 ;
    wire \ppm_encoder_1.aileronZ0Z_3 ;
    wire \ppm_encoder_1.N_289 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ;
    wire \ppm_encoder_1.N_139_17 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ;
    wire \pid_front.stateZ0Z_0 ;
    wire \pid_front.pid_preregZ0Z_8 ;
    wire uart_drone_data_0;
    wire \dron_frame_decoder_1.N_731_0 ;
    wire drone_H_disp_front_0;
    wire \pid_front.error_axb_0 ;
    wire bfn_17_23_0_;
    wire \pid_front.error_axbZ0Z_1 ;
    wire \pid_front.error_1 ;
    wire \pid_front.error_cry_0 ;
    wire \pid_front.error_axbZ0Z_2 ;
    wire \pid_front.error_2 ;
    wire \pid_front.error_cry_1 ;
    wire \pid_front.error_axbZ0Z_3 ;
    wire \pid_front.error_3 ;
    wire \pid_front.error_cry_2 ;
    wire front_command_0;
    wire drone_H_disp_front_i_4;
    wire \pid_front.error_4 ;
    wire \pid_front.error_cry_3 ;
    wire drone_H_disp_front_i_5;
    wire front_command_1;
    wire \pid_front.error_5 ;
    wire \pid_front.error_cry_0_0 ;
    wire drone_H_disp_front_i_6;
    wire front_command_2;
    wire \pid_front.error_6 ;
    wire \pid_front.error_cry_1_0 ;
    wire drone_H_disp_front_i_7;
    wire front_command_3;
    wire \pid_front.error_7 ;
    wire \pid_front.error_cry_2_0 ;
    wire \pid_front.error_cry_3_0 ;
    wire front_command_4;
    wire drone_H_disp_front_i_8;
    wire \pid_front.error_8 ;
    wire bfn_17_24_0_;
    wire drone_H_disp_front_i_9;
    wire front_command_5;
    wire \pid_front.error_9 ;
    wire \pid_front.error_cry_4 ;
    wire front_command_6;
    wire drone_H_disp_front_i_10;
    wire \pid_front.error_10 ;
    wire \pid_front.error_cry_5 ;
    wire \pid_front.error_axbZ0Z_7 ;
    wire \pid_front.error_11 ;
    wire \pid_front.error_cry_6 ;
    wire \pid_front.error_axb_8_l_ofx_0 ;
    wire drone_H_disp_front_12;
    wire \pid_front.error_12 ;
    wire \pid_front.error_cry_7 ;
    wire drone_H_disp_front_i_12;
    wire drone_H_disp_front_13;
    wire \pid_front.error_13 ;
    wire \pid_front.error_cry_8 ;
    wire drone_H_disp_front_i_13;
    wire \pid_front.error_14 ;
    wire \pid_front.error_cry_9 ;
    wire drone_H_disp_front_15;
    wire \pid_front.error_cry_10 ;
    wire \pid_front.error_15 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_1 ;
    wire \ppm_encoder_1.un1_init_pulses_11_9 ;
    wire \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_10_9 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_9 ;
    wire \ppm_encoder_1.un1_init_pulses_0_5 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_8 ;
    wire \ppm_encoder_1.un1_init_pulses_0_8 ;
    wire \ppm_encoder_1.un1_init_pulses_3_axb_15 ;
    wire throttle_order_0;
    wire \ppm_encoder_1.elevatorZ0Z_0 ;
    wire \ppm_encoder_1.throttleZ0Z_0 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ;
    wire \ppm_encoder_1.N_286_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_7 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ;
    wire \ppm_encoder_1.rudderZ0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_16 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_17 ;
    wire \ppm_encoder_1.pulses2countZ0Z_17 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_15 ;
    wire \ppm_encoder_1.pulses2countZ0Z_15 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_18 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_153_d ;
    wire \ppm_encoder_1.pulses2countZ0Z_18 ;
    wire \ppm_encoder_1.init_pulsesZ0Z_16 ;
    wire \ppm_encoder_1.CHOOSE_CHANNEL_d_12 ;
    wire \ppm_encoder_1.PPM_STATE_53_d ;
    wire \ppm_encoder_1.un1_init_pulses_0_axb_16 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ;
    wire \ppm_encoder_1.pulses2countZ0Z_6 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ;
    wire \ppm_encoder_1.pulses2countZ0Z_7 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ;
    wire \ppm_encoder_1.pulses2count_9_sn_N_11_mux ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ;
    wire \ppm_encoder_1.N_1818_0 ;
    wire \ppm_encoder_1.rudderZ0Z_7 ;
    wire \ppm_encoder_1.init_pulses_3_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_0_sqmuxa_0 ;
    wire \ppm_encoder_1.un1_init_pulses_0_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ;
    wire \ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_7 ;
    wire \ppm_encoder_1.N_293_cascade_ ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ;
    wire \ppm_encoder_1.un1_aileron_cry_6_THRU_CO ;
    wire side_order_7;
    wire \ppm_encoder_1.aileronZ0Z_7 ;
    wire \ppm_encoder_1.un1_elevator_cry_6_THRU_CO ;
    wire front_order_7;
    wire \ppm_encoder_1.elevatorZ0Z_7 ;
    wire \ppm_encoder_1.un1_throttle_cry_6_THRU_CO ;
    wire throttle_order_7;
    wire \ppm_encoder_1.throttleZ0Z_7 ;
    wire \ppm_encoder_1.init_pulses_2_sqmuxa_0 ;
    wire \ppm_encoder_1.init_pulses_1_sqmuxa_0 ;
    wire \ppm_encoder_1.un2_throttle_iv_1_4 ;
    wire \ppm_encoder_1.un1_aileron_cry_3_THRU_CO ;
    wire side_order_4;
    wire \ppm_encoder_1.un1_elevator_cry_3_THRU_CO ;
    wire front_order_4;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ;
    wire \ppm_encoder_1.elevatorZ0Z_4 ;
    wire \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ;
    wire \ppm_encoder_1.N_290_cascade_ ;
    wire \ppm_encoder_1.aileronZ0Z_4 ;
    wire \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ;
    wire \ppm_encoder_1.un1_throttle_cry_3_THRU_CO ;
    wire throttle_order_4;
    wire \ppm_encoder_1.throttleZ0Z_4 ;
    wire pid_altitude_dv;
    wire side_order_0;
    wire \ppm_encoder_1.aileronZ0Z_0 ;
    wire \ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ;
    wire bfn_18_17_0_;
    wire \ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_1 ;
    wire \ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_2 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_3 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_4 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_5 ;
    wire \ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_6 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_7 ;
    wire \ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ;
    wire bfn_18_18_0_;
    wire \ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ;
    wire \ppm_encoder_1.counter24_0_data_tmp_8 ;
    wire \ppm_encoder_1.counter24_0_N_2 ;
    wire \ppm_encoder_1.counter24_0_N_2_THRU_CO ;
    wire \ppm_encoder_1.pulses2countZ0Z_4 ;
    wire \ppm_encoder_1.pulses2countZ0Z_5 ;
    wire \ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_10 ;
    wire \ppm_encoder_1.pulses2countZ0Z_11 ;
    wire \ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ;
    wire \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_8 ;
    wire \ppm_encoder_1.pulses2countZ0Z_9 ;
    wire \ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ;
    wire \ppm_encoder_1.pulses2countZ0Z_12 ;
    wire \ppm_encoder_1.pulses2countZ0Z_13 ;
    wire \ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ;
    wire \ppm_encoder_1.N_1818_i ;
    wire \ppm_encoder_1.counterZ0Z_0 ;
    wire bfn_18_19_0_;
    wire \ppm_encoder_1.counterZ0Z_1 ;
    wire \ppm_encoder_1.un1_counter_13_cry_0 ;
    wire \ppm_encoder_1.counterZ0Z_2 ;
    wire \ppm_encoder_1.un1_counter_13_cry_1 ;
    wire \ppm_encoder_1.counterZ0Z_3 ;
    wire \ppm_encoder_1.un1_counter_13_cry_2 ;
    wire \ppm_encoder_1.counterZ0Z_4 ;
    wire \ppm_encoder_1.un1_counter_13_cry_3 ;
    wire \ppm_encoder_1.counterZ0Z_5 ;
    wire \ppm_encoder_1.un1_counter_13_cry_4 ;
    wire \ppm_encoder_1.counterZ0Z_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_5 ;
    wire \ppm_encoder_1.counterZ0Z_7 ;
    wire \ppm_encoder_1.un1_counter_13_cry_6 ;
    wire \ppm_encoder_1.un1_counter_13_cry_7 ;
    wire \ppm_encoder_1.counterZ0Z_8 ;
    wire bfn_18_20_0_;
    wire \ppm_encoder_1.counterZ0Z_9 ;
    wire \ppm_encoder_1.un1_counter_13_cry_8 ;
    wire \ppm_encoder_1.counterZ0Z_10 ;
    wire \ppm_encoder_1.un1_counter_13_cry_9 ;
    wire \ppm_encoder_1.counterZ0Z_11 ;
    wire \ppm_encoder_1.un1_counter_13_cry_10 ;
    wire \ppm_encoder_1.counterZ0Z_12 ;
    wire \ppm_encoder_1.un1_counter_13_cry_11 ;
    wire \ppm_encoder_1.counterZ0Z_13 ;
    wire \ppm_encoder_1.un1_counter_13_cry_12 ;
    wire \ppm_encoder_1.counterZ0Z_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_13 ;
    wire \ppm_encoder_1.counterZ0Z_15 ;
    wire \ppm_encoder_1.un1_counter_13_cry_14 ;
    wire \ppm_encoder_1.un1_counter_13_cry_15 ;
    wire \ppm_encoder_1.counterZ0Z_16 ;
    wire bfn_18_21_0_;
    wire \ppm_encoder_1.counterZ0Z_17 ;
    wire \ppm_encoder_1.un1_counter_13_cry_16 ;
    wire \ppm_encoder_1.un1_counter_13_cry_17 ;
    wire \ppm_encoder_1.counterZ0Z_18 ;
    wire \ppm_encoder_1.N_661_g ;
    wire bfn_18_22_0_;
    wire \pid_front.un1_pid_prereg_cry_1_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_1 ;
    wire \pid_front.un1_pid_prereg_cry_2_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_2 ;
    wire \pid_front.un1_pid_prereg_cry_3_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_3 ;
    wire \pid_front.un1_pid_prereg_cry_4_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_4 ;
    wire \pid_front.un1_pid_prereg_cry_5_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_5 ;
    wire \pid_front.un1_pid_prereg_cry_6_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_6 ;
    wire \pid_front.un1_pid_prereg_cry_7_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_7 ;
    wire \pid_front.un1_pid_prereg_cry_8 ;
    wire \pid_front.un1_pid_prereg_cry_8_THRU_CO ;
    wire bfn_18_23_0_;
    wire \pid_front.un1_pid_prereg_cry_9_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_9 ;
    wire \pid_front.un1_pid_prereg_cry_10_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_10 ;
    wire CONSTANT_ONE_NET;
    wire \pid_front.un1_pid_prereg_cry_11_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_11 ;
    wire \pid_front.un1_pid_prereg_cry_12_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_12 ;
    wire \pid_front.un1_pid_prereg_cry_13_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_13 ;
    wire \pid_front.un1_pid_prereg_cry_14_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_14 ;
    wire \pid_front.un1_pid_prereg_cry_15_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_15 ;
    wire \pid_front.un1_pid_prereg_cry_16 ;
    wire \pid_front.un1_pid_prereg_cry_16_THRU_CO ;
    wire bfn_18_24_0_;
    wire \pid_front.un1_pid_prereg_cry_17_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_17 ;
    wire \pid_front.un1_pid_prereg_cry_18_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_18 ;
    wire \pid_front.un1_pid_prereg_cry_19_THRU_CO ;
    wire \pid_front.un1_pid_prereg_cry_19 ;
    wire \pid_front.un1_pid_prereg_cry_20 ;
    wire \pid_front.pid_preregZ0Z_21 ;
    wire \pid_front.state_0_0 ;
    wire uart_drone_data_6;
    wire drone_H_disp_front_14;
    wire \dron_frame_decoder_1.N_723_0 ;
    wire GB_BUFFER_reset_system_g_THRU_CO;
    wire \pid_side.O_0_4 ;
    wire \pid_side.error_p_regZ0Z_0 ;
    wire \pid_side.O_0_5 ;
    wire \pid_side.state_RNINK4UZ0Z_1 ;
    wire \pid_side.O_0_7 ;
    wire \pid_side.error_p_regZ0Z_3 ;
    wire \pid_front.O_4 ;
    wire \pid_front.error_p_regZ0Z_0 ;
    wire \pid_side.stateZ0Z_0 ;
    wire \pid_side.error_p_regZ0Z_1 ;
    wire \pid_side.pid_preregZ0Z_1 ;
    wire reset_system_g;
    wire \pid_front.state_ns_0 ;
    wire reset_system;
    wire \pid_front.O_5 ;
    wire \pid_front.error_p_regZ0Z_1 ;
    wire \pid_front.O_13 ;
    wire \pid_front.error_p_regZ0Z_9 ;
    wire \pid_front.O_6 ;
    wire \pid_front.error_p_regZ0Z_2 ;
    wire \pid_front.O_9 ;
    wire \pid_front.error_p_regZ0Z_5 ;
    wire \pid_front.O_8 ;
    wire \pid_front.error_p_regZ0Z_4 ;
    wire \pid_front.O_18 ;
    wire \pid_front.error_p_regZ0Z_14 ;
    wire \pid_front.O_12 ;
    wire \pid_front.error_p_regZ0Z_8 ;
    wire \pid_front.O_14 ;
    wire \pid_front.error_p_regZ0Z_10 ;
    wire \pid_front.O_11 ;
    wire \pid_front.error_p_regZ0Z_7 ;
    wire \pid_front.O_7 ;
    wire \pid_front.error_p_regZ0Z_3 ;
    wire \pid_front.O_20 ;
    wire \pid_front.error_p_regZ0Z_16 ;
    wire \pid_front.O_10 ;
    wire \pid_front.error_p_regZ0Z_6 ;
    wire \pid_front.O_22 ;
    wire \pid_front.error_p_regZ0Z_18 ;
    wire \pid_front.O_23 ;
    wire \pid_front.error_p_regZ0Z_19 ;
    wire \pid_front.O_17 ;
    wire \pid_front.error_p_regZ0Z_13 ;
    wire \pid_front.O_19 ;
    wire \pid_front.error_p_regZ0Z_15 ;
    wire \pid_front.O_15 ;
    wire \pid_front.error_p_regZ0Z_11 ;
    wire \pid_front.O_16 ;
    wire \pid_front.error_p_regZ0Z_12 ;
    wire \pid_front.O_24 ;
    wire \pid_front.error_p_regZ0Z_20 ;
    wire \pid_front.state_RNIVIRQZ0Z_1 ;
    wire \pid_front.O_21 ;
    wire \pid_front.error_p_regZ0Z_17 ;
    wire _gnd_net_;
    wire clk_system_c_g;
    wire N_851_g;

    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48236),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48235),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__22032,N__22089,N__21468,N__21520,N__21573,N__21630,N__21696,N__21759,N__21810,N__21873,N__21169,N__21225,N__21303,N__21342,N__21396,N__34334}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__21944,N__20234,N__20246,N__25973,N__20261,N__20273,N__21956,N__23333}),
            .OHOLDTOP(),
            .O({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,\pid_alt.O_3_24 ,\pid_alt.O_3_23 ,\pid_alt.O_3_22 ,\pid_alt.O_3_21 ,\pid_alt.O_3_20 ,\pid_alt.O_3_19 ,\pid_alt.O_3_18 ,\pid_alt.O_3_17 ,\pid_alt.O_3_16 ,\pid_alt.O_3_15 ,\pid_alt.O_3_14 ,\pid_alt.O_3_13 ,\pid_alt.O_3_12 ,\pid_alt.O_3_11 ,\pid_alt.O_3_10 ,\pid_alt.O_3_9 ,\pid_alt.O_3_8 ,\pid_alt.O_3_7 ,\pid_alt.O_3_6 ,\pid_alt.O_3_5 ,\pid_alt.O_3_4 ,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50}));
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_1_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_1_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48206),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48199),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66}),
            .ADDSUBBOT(),
            .A({N__22033,N__22090,N__21475,N__21519,N__21574,N__21631,N__21697,N__21763,N__21811,N__21883,N__21165,N__21232,N__21304,N__21343,N__21397,N__34327}),
            .C({dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82}),
            .B({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,N__27089,N__38870,N__19781,N__19697,N__19661,N__19673,N__19685,N__19709}),
            .OHOLDTOP(),
            .O({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,\pid_alt.O_2_24 ,\pid_alt.O_2_23 ,\pid_alt.O_2_22 ,\pid_alt.O_2_21 ,\pid_alt.O_2_20 ,\pid_alt.O_2_19 ,\pid_alt.O_2_18 ,\pid_alt.O_2_17 ,\pid_alt.O_2_16 ,\pid_alt.O_2_15 ,\pid_alt.O_2_14 ,\pid_alt.O_2_13 ,\pid_alt.O_2_12 ,\pid_alt.O_2_11 ,\pid_alt.O_2_10 ,\pid_alt.O_2_9 ,\pid_alt.O_2_8 ,\pid_alt.O_2_7 ,\pid_alt.O_2_6 ,\pid_alt.O_2_5 ,\pid_alt.O_2_4 ,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101}));
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_alt.un2_error_2_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_alt.un2_error_2_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48230),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48229),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117}),
            .ADDSUBBOT(),
            .A({N__22037,N__22097,N__21479,N__21527,N__21575,N__21635,N__21701,N__21767,N__21815,N__21884,N__21170,N__21239,N__21308,N__21350,N__21398,N__34326}),
            .C({dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133}),
            .B({dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,N__19583,N__19601,N__19745,N__20198,N__20222,N__19592,N__19733,N__20210}),
            .OHOLDTOP(),
            .O({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,\pid_alt.O_1_24 ,\pid_alt.O_1_23 ,\pid_alt.O_1_22 ,\pid_alt.O_1_21 ,\pid_alt.O_1_20 ,\pid_alt.O_1_19 ,\pid_alt.O_1_18 ,\pid_alt.O_1_17 ,\pid_alt.O_1_16 ,\pid_alt.O_1_15 ,\pid_alt.O_1_14 ,\pid_alt.O_1_13 ,\pid_alt.O_1_12 ,\pid_alt.O_1_11 ,\pid_alt.O_1_10 ,\pid_alt.O_1_9 ,\pid_alt.O_1_8 ,\pid_alt.O_1_7 ,\pid_alt.O_1_6 ,\pid_alt.O_1_5 ,\pid_alt.O_1_4 ,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}));
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_front.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_front.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_front.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48234),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48233),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168}),
            .ADDSUBBOT(),
            .A({N__43391,N__43424,N__43451,N__43499,N__43553,N__43577,N__43610,N__42875,N__42914,N__42947,N__42980,N__43013,N__43046,N__43076,N__42443,N__42482}),
            .C({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .B({dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__30757,N__25076,N__39067,N__26756,N__29504,N__25112,N__30796,N__25142}),
            .OHOLDTOP(),
            .O({dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,\pid_front.O_24 ,\pid_front.O_23 ,\pid_front.O_22 ,\pid_front.O_21 ,\pid_front.O_20 ,\pid_front.O_19 ,\pid_front.O_18 ,\pid_front.O_17 ,\pid_front.O_16 ,\pid_front.O_15 ,\pid_front.O_14 ,\pid_front.O_13 ,\pid_front.O_12 ,\pid_front.O_11 ,\pid_front.O_10 ,\pid_front.O_9 ,\pid_front.O_8 ,\pid_front.O_7 ,\pid_front.O_6 ,\pid_front.O_5 ,\pid_front.O_4 ,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203}));
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .NEG_TRIGGER=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .MODE_8x8=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .D_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .C_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_SIGNED=1'b1;
    defparam \pid_side.un2_error_mulonly_0_24_0 .B_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pid_side.un2_error_mulonly_0_24_0 .A_SIGNED=1'b1;
    SB_MAC16 \pid_side.un2_error_mulonly_0_24_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__48193),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__48192),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219}),
            .ADDSUBBOT(),
            .A({N__23345,N__23366,N__23384,N__23402,N__23420,N__23438,N__23468,N__23495,N__23216,N__23234,N__23249,N__23264,N__23282,N__23297,N__23315,N__27158}),
            .C({dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235}),
            .B({dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,N__30758,N__25069,N__39071,N__26755,N__29503,N__25105,N__30797,N__25141}),
            .OHOLDTOP(),
            .O({dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,\pid_side.O_0_24 ,\pid_side.O_0_23 ,\pid_side.O_0_22 ,\pid_side.O_0_21 ,\pid_side.O_0_20 ,\pid_side.O_0_19 ,\pid_side.O_0_18 ,\pid_side.O_0_17 ,\pid_side.O_0_16 ,\pid_side.O_0_15 ,\pid_side.O_0_14 ,\pid_side.O_0_13 ,\pid_side.O_0_12 ,\pid_side.O_0_11 ,\pid_side.O_0_10 ,\pid_side.O_0_9 ,\pid_side.O_0_8 ,\pid_side.O_0_7 ,\pid_side.O_0_6 ,\pid_side.O_0_5 ,\pid_side.O_0_4 ,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254}));
    PRE_IO_GBUF clk_system_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__52029),
            .GLOBALBUFFEROUTPUT(clk_system_c_g));
    defparam clk_system_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_system_ibuf_gb_io_iopad (
            .OE(N__52031),
            .DIN(N__52030),
            .DOUT(N__52029),
            .PACKAGEPIN(clk_system));
    defparam clk_system_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_system_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_system_ibuf_gb_io_preio (
            .PADOEN(N__52031),
            .PADOUT(N__52030),
            .PADIN(N__52029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_drone_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_drone_ibuf_iopad (
            .OE(N__52020),
            .DIN(N__52019),
            .DOUT(N__52018),
            .PACKAGEPIN(uart_input_drone));
    defparam uart_input_drone_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_drone_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_drone_ibuf_preio (
            .PADOEN(N__52020),
            .PADOUT(N__52019),
            .PADIN(N__52018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_drone_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam uart_input_pc_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD uart_input_pc_ibuf_iopad (
            .OE(N__52011),
            .DIN(N__52010),
            .DOUT(N__52009),
            .PACKAGEPIN(uart_input_pc));
    defparam uart_input_pc_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam uart_input_pc_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO uart_input_pc_ibuf_preio (
            .PADOEN(N__52011),
            .PADOUT(N__52010),
            .PADIN(N__52009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(uart_input_pc_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH2_18A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH2_18A_obuf_iopad (
            .OE(N__52002),
            .DIN(N__52001),
            .DOUT(N__52000),
            .PACKAGEPIN(debug_CH2_18A));
    defparam debug_CH2_18A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH2_18A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH2_18A_obuf_preio (
            .PADOEN(N__52002),
            .PADOUT(N__52001),
            .PADIN(N__52000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__40706),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH0_16A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH0_16A_obuf_iopad (
            .OE(N__51993),
            .DIN(N__51992),
            .DOUT(N__51991),
            .PACKAGEPIN(debug_CH0_16A));
    defparam debug_CH0_16A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH0_16A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH0_16A_obuf_preio (
            .PADOEN(N__51993),
            .PADOUT(N__51992),
            .PADIN(N__51991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH1_0A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH1_0A_obuf_iopad (
            .OE(N__51984),
            .DIN(N__51983),
            .DOUT(N__51982),
            .PACKAGEPIN(debug_CH1_0A));
    defparam debug_CH1_0A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH1_0A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH1_0A_obuf_preio (
            .PADOEN(N__51984),
            .PADOUT(N__51983),
            .PADIN(N__51982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH5_31B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH5_31B_obuf_iopad (
            .OE(N__51975),
            .DIN(N__51974),
            .DOUT(N__51973),
            .PACKAGEPIN(debug_CH5_31B));
    defparam debug_CH5_31B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH5_31B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH5_31B_obuf_preio (
            .PADOEN(N__51975),
            .PADOUT(N__51974),
            .PADIN(N__51973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH4_2A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH4_2A_obuf_iopad (
            .OE(N__51966),
            .DIN(N__51965),
            .DOUT(N__51964),
            .PACKAGEPIN(debug_CH4_2A));
    defparam debug_CH4_2A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH4_2A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH4_2A_obuf_preio (
            .PADOEN(N__51966),
            .PADOUT(N__51965),
            .PADIN(N__51964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ppm_output_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD ppm_output_obuf_iopad (
            .OE(N__51957),
            .DIN(N__51956),
            .DOUT(N__51955),
            .PACKAGEPIN(ppm_output));
    defparam ppm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ppm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ppm_output_obuf_preio (
            .PADOEN(N__51957),
            .PADOUT(N__51956),
            .PADIN(N__51955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32519),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH3_20A_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH3_20A_obuf_iopad (
            .OE(N__51948),
            .DIN(N__51947),
            .DOUT(N__51946),
            .PACKAGEPIN(debug_CH3_20A));
    defparam debug_CH3_20A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH3_20A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH3_20A_obuf_preio (
            .PADOEN(N__51948),
            .PADOUT(N__51947),
            .PADIN(N__51946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27203),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam debug_CH6_5B_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD debug_CH6_5B_obuf_iopad (
            .OE(N__51939),
            .DIN(N__51938),
            .DOUT(N__51937),
            .PACKAGEPIN(debug_CH6_5B));
    defparam debug_CH6_5B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam debug_CH6_5B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_CH6_5B_obuf_preio (
            .PADOEN(N__51939),
            .PADOUT(N__51938),
            .PADIN(N__51937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12609 (
            .O(N__51920),
            .I(N__51917));
    LocalMux I__12608 (
            .O(N__51917),
            .I(N__51914));
    Odrv4 I__12607 (
            .O(N__51914),
            .I(\pid_front.O_23 ));
    CascadeMux I__12606 (
            .O(N__51911),
            .I(N__51908));
    InMux I__12605 (
            .O(N__51908),
            .I(N__51904));
    InMux I__12604 (
            .O(N__51907),
            .I(N__51901));
    LocalMux I__12603 (
            .O(N__51904),
            .I(N__51898));
    LocalMux I__12602 (
            .O(N__51901),
            .I(N__51895));
    Sp12to4 I__12601 (
            .O(N__51898),
            .I(N__51892));
    Span4Mux_h I__12600 (
            .O(N__51895),
            .I(N__51888));
    Span12Mux_h I__12599 (
            .O(N__51892),
            .I(N__51885));
    InMux I__12598 (
            .O(N__51891),
            .I(N__51882));
    Span4Mux_h I__12597 (
            .O(N__51888),
            .I(N__51879));
    Odrv12 I__12596 (
            .O(N__51885),
            .I(\pid_front.error_p_regZ0Z_19 ));
    LocalMux I__12595 (
            .O(N__51882),
            .I(\pid_front.error_p_regZ0Z_19 ));
    Odrv4 I__12594 (
            .O(N__51879),
            .I(\pid_front.error_p_regZ0Z_19 ));
    InMux I__12593 (
            .O(N__51872),
            .I(N__51869));
    LocalMux I__12592 (
            .O(N__51869),
            .I(N__51866));
    Odrv4 I__12591 (
            .O(N__51866),
            .I(\pid_front.O_17 ));
    InMux I__12590 (
            .O(N__51863),
            .I(N__51860));
    LocalMux I__12589 (
            .O(N__51860),
            .I(N__51857));
    Span4Mux_h I__12588 (
            .O(N__51857),
            .I(N__51852));
    InMux I__12587 (
            .O(N__51856),
            .I(N__51849));
    InMux I__12586 (
            .O(N__51855),
            .I(N__51846));
    Sp12to4 I__12585 (
            .O(N__51852),
            .I(N__51841));
    LocalMux I__12584 (
            .O(N__51849),
            .I(N__51841));
    LocalMux I__12583 (
            .O(N__51846),
            .I(\pid_front.error_p_regZ0Z_13 ));
    Odrv12 I__12582 (
            .O(N__51841),
            .I(\pid_front.error_p_regZ0Z_13 ));
    InMux I__12581 (
            .O(N__51836),
            .I(N__51833));
    LocalMux I__12580 (
            .O(N__51833),
            .I(N__51830));
    Odrv4 I__12579 (
            .O(N__51830),
            .I(\pid_front.O_19 ));
    InMux I__12578 (
            .O(N__51827),
            .I(N__51824));
    LocalMux I__12577 (
            .O(N__51824),
            .I(N__51819));
    InMux I__12576 (
            .O(N__51823),
            .I(N__51816));
    InMux I__12575 (
            .O(N__51822),
            .I(N__51813));
    Sp12to4 I__12574 (
            .O(N__51819),
            .I(N__51808));
    LocalMux I__12573 (
            .O(N__51816),
            .I(N__51808));
    LocalMux I__12572 (
            .O(N__51813),
            .I(\pid_front.error_p_regZ0Z_15 ));
    Odrv12 I__12571 (
            .O(N__51808),
            .I(\pid_front.error_p_regZ0Z_15 ));
    InMux I__12570 (
            .O(N__51803),
            .I(N__51800));
    LocalMux I__12569 (
            .O(N__51800),
            .I(\pid_front.O_15 ));
    InMux I__12568 (
            .O(N__51797),
            .I(N__51792));
    InMux I__12567 (
            .O(N__51796),
            .I(N__51789));
    InMux I__12566 (
            .O(N__51795),
            .I(N__51786));
    LocalMux I__12565 (
            .O(N__51792),
            .I(N__51781));
    LocalMux I__12564 (
            .O(N__51789),
            .I(N__51781));
    LocalMux I__12563 (
            .O(N__51786),
            .I(\pid_front.error_p_regZ0Z_11 ));
    Odrv12 I__12562 (
            .O(N__51781),
            .I(\pid_front.error_p_regZ0Z_11 ));
    InMux I__12561 (
            .O(N__51776),
            .I(N__51773));
    LocalMux I__12560 (
            .O(N__51773),
            .I(N__51770));
    Odrv4 I__12559 (
            .O(N__51770),
            .I(\pid_front.O_16 ));
    InMux I__12558 (
            .O(N__51767),
            .I(N__51764));
    LocalMux I__12557 (
            .O(N__51764),
            .I(N__51761));
    Span4Mux_h I__12556 (
            .O(N__51761),
            .I(N__51757));
    InMux I__12555 (
            .O(N__51760),
            .I(N__51754));
    Span4Mux_h I__12554 (
            .O(N__51757),
            .I(N__51751));
    LocalMux I__12553 (
            .O(N__51754),
            .I(N__51747));
    Span4Mux_h I__12552 (
            .O(N__51751),
            .I(N__51744));
    InMux I__12551 (
            .O(N__51750),
            .I(N__51741));
    Span4Mux_h I__12550 (
            .O(N__51747),
            .I(N__51738));
    Odrv4 I__12549 (
            .O(N__51744),
            .I(\pid_front.error_p_regZ0Z_12 ));
    LocalMux I__12548 (
            .O(N__51741),
            .I(\pid_front.error_p_regZ0Z_12 ));
    Odrv4 I__12547 (
            .O(N__51738),
            .I(\pid_front.error_p_regZ0Z_12 ));
    InMux I__12546 (
            .O(N__51731),
            .I(N__51728));
    LocalMux I__12545 (
            .O(N__51728),
            .I(N__51725));
    Odrv4 I__12544 (
            .O(N__51725),
            .I(\pid_front.O_24 ));
    CascadeMux I__12543 (
            .O(N__51722),
            .I(N__51719));
    InMux I__12542 (
            .O(N__51719),
            .I(N__51716));
    LocalMux I__12541 (
            .O(N__51716),
            .I(N__51713));
    Span4Mux_h I__12540 (
            .O(N__51713),
            .I(N__51708));
    InMux I__12539 (
            .O(N__51712),
            .I(N__51703));
    InMux I__12538 (
            .O(N__51711),
            .I(N__51703));
    Span4Mux_h I__12537 (
            .O(N__51708),
            .I(N__51700));
    LocalMux I__12536 (
            .O(N__51703),
            .I(N__51696));
    Span4Mux_h I__12535 (
            .O(N__51700),
            .I(N__51693));
    InMux I__12534 (
            .O(N__51699),
            .I(N__51690));
    Span4Mux_h I__12533 (
            .O(N__51696),
            .I(N__51687));
    Odrv4 I__12532 (
            .O(N__51693),
            .I(\pid_front.error_p_regZ0Z_20 ));
    LocalMux I__12531 (
            .O(N__51690),
            .I(\pid_front.error_p_regZ0Z_20 ));
    Odrv4 I__12530 (
            .O(N__51687),
            .I(\pid_front.error_p_regZ0Z_20 ));
    CascadeMux I__12529 (
            .O(N__51680),
            .I(N__51672));
    InMux I__12528 (
            .O(N__51679),
            .I(N__51652));
    InMux I__12527 (
            .O(N__51678),
            .I(N__51652));
    InMux I__12526 (
            .O(N__51677),
            .I(N__51645));
    InMux I__12525 (
            .O(N__51676),
            .I(N__51645));
    InMux I__12524 (
            .O(N__51675),
            .I(N__51645));
    InMux I__12523 (
            .O(N__51672),
            .I(N__51640));
    InMux I__12522 (
            .O(N__51671),
            .I(N__51640));
    InMux I__12521 (
            .O(N__51670),
            .I(N__51629));
    InMux I__12520 (
            .O(N__51669),
            .I(N__51629));
    InMux I__12519 (
            .O(N__51668),
            .I(N__51629));
    InMux I__12518 (
            .O(N__51667),
            .I(N__51629));
    InMux I__12517 (
            .O(N__51666),
            .I(N__51629));
    InMux I__12516 (
            .O(N__51665),
            .I(N__51618));
    InMux I__12515 (
            .O(N__51664),
            .I(N__51618));
    InMux I__12514 (
            .O(N__51663),
            .I(N__51618));
    InMux I__12513 (
            .O(N__51662),
            .I(N__51618));
    InMux I__12512 (
            .O(N__51661),
            .I(N__51618));
    InMux I__12511 (
            .O(N__51660),
            .I(N__51613));
    InMux I__12510 (
            .O(N__51659),
            .I(N__51613));
    InMux I__12509 (
            .O(N__51658),
            .I(N__51610));
    InMux I__12508 (
            .O(N__51657),
            .I(N__51607));
    LocalMux I__12507 (
            .O(N__51652),
            .I(N__51602));
    LocalMux I__12506 (
            .O(N__51645),
            .I(N__51602));
    LocalMux I__12505 (
            .O(N__51640),
            .I(N__51595));
    LocalMux I__12504 (
            .O(N__51629),
            .I(N__51595));
    LocalMux I__12503 (
            .O(N__51618),
            .I(N__51595));
    LocalMux I__12502 (
            .O(N__51613),
            .I(N__51592));
    LocalMux I__12501 (
            .O(N__51610),
            .I(N__51587));
    LocalMux I__12500 (
            .O(N__51607),
            .I(N__51587));
    Span4Mux_v I__12499 (
            .O(N__51602),
            .I(N__51582));
    Span4Mux_v I__12498 (
            .O(N__51595),
            .I(N__51582));
    Odrv4 I__12497 (
            .O(N__51592),
            .I(\pid_front.state_RNIVIRQZ0Z_1 ));
    Odrv4 I__12496 (
            .O(N__51587),
            .I(\pid_front.state_RNIVIRQZ0Z_1 ));
    Odrv4 I__12495 (
            .O(N__51582),
            .I(\pid_front.state_RNIVIRQZ0Z_1 ));
    InMux I__12494 (
            .O(N__51575),
            .I(N__51572));
    LocalMux I__12493 (
            .O(N__51572),
            .I(\pid_front.O_21 ));
    InMux I__12492 (
            .O(N__51569),
            .I(N__51566));
    LocalMux I__12491 (
            .O(N__51566),
            .I(N__51563));
    Span4Mux_v I__12490 (
            .O(N__51563),
            .I(N__51558));
    InMux I__12489 (
            .O(N__51562),
            .I(N__51555));
    InMux I__12488 (
            .O(N__51561),
            .I(N__51552));
    Sp12to4 I__12487 (
            .O(N__51558),
            .I(N__51547));
    LocalMux I__12486 (
            .O(N__51555),
            .I(N__51547));
    LocalMux I__12485 (
            .O(N__51552),
            .I(\pid_front.error_p_regZ0Z_17 ));
    Odrv12 I__12484 (
            .O(N__51547),
            .I(\pid_front.error_p_regZ0Z_17 ));
    ClkMux I__12483 (
            .O(N__51542),
            .I(N__50831));
    ClkMux I__12482 (
            .O(N__51541),
            .I(N__50831));
    ClkMux I__12481 (
            .O(N__51540),
            .I(N__50831));
    ClkMux I__12480 (
            .O(N__51539),
            .I(N__50831));
    ClkMux I__12479 (
            .O(N__51538),
            .I(N__50831));
    ClkMux I__12478 (
            .O(N__51537),
            .I(N__50831));
    ClkMux I__12477 (
            .O(N__51536),
            .I(N__50831));
    ClkMux I__12476 (
            .O(N__51535),
            .I(N__50831));
    ClkMux I__12475 (
            .O(N__51534),
            .I(N__50831));
    ClkMux I__12474 (
            .O(N__51533),
            .I(N__50831));
    ClkMux I__12473 (
            .O(N__51532),
            .I(N__50831));
    ClkMux I__12472 (
            .O(N__51531),
            .I(N__50831));
    ClkMux I__12471 (
            .O(N__51530),
            .I(N__50831));
    ClkMux I__12470 (
            .O(N__51529),
            .I(N__50831));
    ClkMux I__12469 (
            .O(N__51528),
            .I(N__50831));
    ClkMux I__12468 (
            .O(N__51527),
            .I(N__50831));
    ClkMux I__12467 (
            .O(N__51526),
            .I(N__50831));
    ClkMux I__12466 (
            .O(N__51525),
            .I(N__50831));
    ClkMux I__12465 (
            .O(N__51524),
            .I(N__50831));
    ClkMux I__12464 (
            .O(N__51523),
            .I(N__50831));
    ClkMux I__12463 (
            .O(N__51522),
            .I(N__50831));
    ClkMux I__12462 (
            .O(N__51521),
            .I(N__50831));
    ClkMux I__12461 (
            .O(N__51520),
            .I(N__50831));
    ClkMux I__12460 (
            .O(N__51519),
            .I(N__50831));
    ClkMux I__12459 (
            .O(N__51518),
            .I(N__50831));
    ClkMux I__12458 (
            .O(N__51517),
            .I(N__50831));
    ClkMux I__12457 (
            .O(N__51516),
            .I(N__50831));
    ClkMux I__12456 (
            .O(N__51515),
            .I(N__50831));
    ClkMux I__12455 (
            .O(N__51514),
            .I(N__50831));
    ClkMux I__12454 (
            .O(N__51513),
            .I(N__50831));
    ClkMux I__12453 (
            .O(N__51512),
            .I(N__50831));
    ClkMux I__12452 (
            .O(N__51511),
            .I(N__50831));
    ClkMux I__12451 (
            .O(N__51510),
            .I(N__50831));
    ClkMux I__12450 (
            .O(N__51509),
            .I(N__50831));
    ClkMux I__12449 (
            .O(N__51508),
            .I(N__50831));
    ClkMux I__12448 (
            .O(N__51507),
            .I(N__50831));
    ClkMux I__12447 (
            .O(N__51506),
            .I(N__50831));
    ClkMux I__12446 (
            .O(N__51505),
            .I(N__50831));
    ClkMux I__12445 (
            .O(N__51504),
            .I(N__50831));
    ClkMux I__12444 (
            .O(N__51503),
            .I(N__50831));
    ClkMux I__12443 (
            .O(N__51502),
            .I(N__50831));
    ClkMux I__12442 (
            .O(N__51501),
            .I(N__50831));
    ClkMux I__12441 (
            .O(N__51500),
            .I(N__50831));
    ClkMux I__12440 (
            .O(N__51499),
            .I(N__50831));
    ClkMux I__12439 (
            .O(N__51498),
            .I(N__50831));
    ClkMux I__12438 (
            .O(N__51497),
            .I(N__50831));
    ClkMux I__12437 (
            .O(N__51496),
            .I(N__50831));
    ClkMux I__12436 (
            .O(N__51495),
            .I(N__50831));
    ClkMux I__12435 (
            .O(N__51494),
            .I(N__50831));
    ClkMux I__12434 (
            .O(N__51493),
            .I(N__50831));
    ClkMux I__12433 (
            .O(N__51492),
            .I(N__50831));
    ClkMux I__12432 (
            .O(N__51491),
            .I(N__50831));
    ClkMux I__12431 (
            .O(N__51490),
            .I(N__50831));
    ClkMux I__12430 (
            .O(N__51489),
            .I(N__50831));
    ClkMux I__12429 (
            .O(N__51488),
            .I(N__50831));
    ClkMux I__12428 (
            .O(N__51487),
            .I(N__50831));
    ClkMux I__12427 (
            .O(N__51486),
            .I(N__50831));
    ClkMux I__12426 (
            .O(N__51485),
            .I(N__50831));
    ClkMux I__12425 (
            .O(N__51484),
            .I(N__50831));
    ClkMux I__12424 (
            .O(N__51483),
            .I(N__50831));
    ClkMux I__12423 (
            .O(N__51482),
            .I(N__50831));
    ClkMux I__12422 (
            .O(N__51481),
            .I(N__50831));
    ClkMux I__12421 (
            .O(N__51480),
            .I(N__50831));
    ClkMux I__12420 (
            .O(N__51479),
            .I(N__50831));
    ClkMux I__12419 (
            .O(N__51478),
            .I(N__50831));
    ClkMux I__12418 (
            .O(N__51477),
            .I(N__50831));
    ClkMux I__12417 (
            .O(N__51476),
            .I(N__50831));
    ClkMux I__12416 (
            .O(N__51475),
            .I(N__50831));
    ClkMux I__12415 (
            .O(N__51474),
            .I(N__50831));
    ClkMux I__12414 (
            .O(N__51473),
            .I(N__50831));
    ClkMux I__12413 (
            .O(N__51472),
            .I(N__50831));
    ClkMux I__12412 (
            .O(N__51471),
            .I(N__50831));
    ClkMux I__12411 (
            .O(N__51470),
            .I(N__50831));
    ClkMux I__12410 (
            .O(N__51469),
            .I(N__50831));
    ClkMux I__12409 (
            .O(N__51468),
            .I(N__50831));
    ClkMux I__12408 (
            .O(N__51467),
            .I(N__50831));
    ClkMux I__12407 (
            .O(N__51466),
            .I(N__50831));
    ClkMux I__12406 (
            .O(N__51465),
            .I(N__50831));
    ClkMux I__12405 (
            .O(N__51464),
            .I(N__50831));
    ClkMux I__12404 (
            .O(N__51463),
            .I(N__50831));
    ClkMux I__12403 (
            .O(N__51462),
            .I(N__50831));
    ClkMux I__12402 (
            .O(N__51461),
            .I(N__50831));
    ClkMux I__12401 (
            .O(N__51460),
            .I(N__50831));
    ClkMux I__12400 (
            .O(N__51459),
            .I(N__50831));
    ClkMux I__12399 (
            .O(N__51458),
            .I(N__50831));
    ClkMux I__12398 (
            .O(N__51457),
            .I(N__50831));
    ClkMux I__12397 (
            .O(N__51456),
            .I(N__50831));
    ClkMux I__12396 (
            .O(N__51455),
            .I(N__50831));
    ClkMux I__12395 (
            .O(N__51454),
            .I(N__50831));
    ClkMux I__12394 (
            .O(N__51453),
            .I(N__50831));
    ClkMux I__12393 (
            .O(N__51452),
            .I(N__50831));
    ClkMux I__12392 (
            .O(N__51451),
            .I(N__50831));
    ClkMux I__12391 (
            .O(N__51450),
            .I(N__50831));
    ClkMux I__12390 (
            .O(N__51449),
            .I(N__50831));
    ClkMux I__12389 (
            .O(N__51448),
            .I(N__50831));
    ClkMux I__12388 (
            .O(N__51447),
            .I(N__50831));
    ClkMux I__12387 (
            .O(N__51446),
            .I(N__50831));
    ClkMux I__12386 (
            .O(N__51445),
            .I(N__50831));
    ClkMux I__12385 (
            .O(N__51444),
            .I(N__50831));
    ClkMux I__12384 (
            .O(N__51443),
            .I(N__50831));
    ClkMux I__12383 (
            .O(N__51442),
            .I(N__50831));
    ClkMux I__12382 (
            .O(N__51441),
            .I(N__50831));
    ClkMux I__12381 (
            .O(N__51440),
            .I(N__50831));
    ClkMux I__12380 (
            .O(N__51439),
            .I(N__50831));
    ClkMux I__12379 (
            .O(N__51438),
            .I(N__50831));
    ClkMux I__12378 (
            .O(N__51437),
            .I(N__50831));
    ClkMux I__12377 (
            .O(N__51436),
            .I(N__50831));
    ClkMux I__12376 (
            .O(N__51435),
            .I(N__50831));
    ClkMux I__12375 (
            .O(N__51434),
            .I(N__50831));
    ClkMux I__12374 (
            .O(N__51433),
            .I(N__50831));
    ClkMux I__12373 (
            .O(N__51432),
            .I(N__50831));
    ClkMux I__12372 (
            .O(N__51431),
            .I(N__50831));
    ClkMux I__12371 (
            .O(N__51430),
            .I(N__50831));
    ClkMux I__12370 (
            .O(N__51429),
            .I(N__50831));
    ClkMux I__12369 (
            .O(N__51428),
            .I(N__50831));
    ClkMux I__12368 (
            .O(N__51427),
            .I(N__50831));
    ClkMux I__12367 (
            .O(N__51426),
            .I(N__50831));
    ClkMux I__12366 (
            .O(N__51425),
            .I(N__50831));
    ClkMux I__12365 (
            .O(N__51424),
            .I(N__50831));
    ClkMux I__12364 (
            .O(N__51423),
            .I(N__50831));
    ClkMux I__12363 (
            .O(N__51422),
            .I(N__50831));
    ClkMux I__12362 (
            .O(N__51421),
            .I(N__50831));
    ClkMux I__12361 (
            .O(N__51420),
            .I(N__50831));
    ClkMux I__12360 (
            .O(N__51419),
            .I(N__50831));
    ClkMux I__12359 (
            .O(N__51418),
            .I(N__50831));
    ClkMux I__12358 (
            .O(N__51417),
            .I(N__50831));
    ClkMux I__12357 (
            .O(N__51416),
            .I(N__50831));
    ClkMux I__12356 (
            .O(N__51415),
            .I(N__50831));
    ClkMux I__12355 (
            .O(N__51414),
            .I(N__50831));
    ClkMux I__12354 (
            .O(N__51413),
            .I(N__50831));
    ClkMux I__12353 (
            .O(N__51412),
            .I(N__50831));
    ClkMux I__12352 (
            .O(N__51411),
            .I(N__50831));
    ClkMux I__12351 (
            .O(N__51410),
            .I(N__50831));
    ClkMux I__12350 (
            .O(N__51409),
            .I(N__50831));
    ClkMux I__12349 (
            .O(N__51408),
            .I(N__50831));
    ClkMux I__12348 (
            .O(N__51407),
            .I(N__50831));
    ClkMux I__12347 (
            .O(N__51406),
            .I(N__50831));
    ClkMux I__12346 (
            .O(N__51405),
            .I(N__50831));
    ClkMux I__12345 (
            .O(N__51404),
            .I(N__50831));
    ClkMux I__12344 (
            .O(N__51403),
            .I(N__50831));
    ClkMux I__12343 (
            .O(N__51402),
            .I(N__50831));
    ClkMux I__12342 (
            .O(N__51401),
            .I(N__50831));
    ClkMux I__12341 (
            .O(N__51400),
            .I(N__50831));
    ClkMux I__12340 (
            .O(N__51399),
            .I(N__50831));
    ClkMux I__12339 (
            .O(N__51398),
            .I(N__50831));
    ClkMux I__12338 (
            .O(N__51397),
            .I(N__50831));
    ClkMux I__12337 (
            .O(N__51396),
            .I(N__50831));
    ClkMux I__12336 (
            .O(N__51395),
            .I(N__50831));
    ClkMux I__12335 (
            .O(N__51394),
            .I(N__50831));
    ClkMux I__12334 (
            .O(N__51393),
            .I(N__50831));
    ClkMux I__12333 (
            .O(N__51392),
            .I(N__50831));
    ClkMux I__12332 (
            .O(N__51391),
            .I(N__50831));
    ClkMux I__12331 (
            .O(N__51390),
            .I(N__50831));
    ClkMux I__12330 (
            .O(N__51389),
            .I(N__50831));
    ClkMux I__12329 (
            .O(N__51388),
            .I(N__50831));
    ClkMux I__12328 (
            .O(N__51387),
            .I(N__50831));
    ClkMux I__12327 (
            .O(N__51386),
            .I(N__50831));
    ClkMux I__12326 (
            .O(N__51385),
            .I(N__50831));
    ClkMux I__12325 (
            .O(N__51384),
            .I(N__50831));
    ClkMux I__12324 (
            .O(N__51383),
            .I(N__50831));
    ClkMux I__12323 (
            .O(N__51382),
            .I(N__50831));
    ClkMux I__12322 (
            .O(N__51381),
            .I(N__50831));
    ClkMux I__12321 (
            .O(N__51380),
            .I(N__50831));
    ClkMux I__12320 (
            .O(N__51379),
            .I(N__50831));
    ClkMux I__12319 (
            .O(N__51378),
            .I(N__50831));
    ClkMux I__12318 (
            .O(N__51377),
            .I(N__50831));
    ClkMux I__12317 (
            .O(N__51376),
            .I(N__50831));
    ClkMux I__12316 (
            .O(N__51375),
            .I(N__50831));
    ClkMux I__12315 (
            .O(N__51374),
            .I(N__50831));
    ClkMux I__12314 (
            .O(N__51373),
            .I(N__50831));
    ClkMux I__12313 (
            .O(N__51372),
            .I(N__50831));
    ClkMux I__12312 (
            .O(N__51371),
            .I(N__50831));
    ClkMux I__12311 (
            .O(N__51370),
            .I(N__50831));
    ClkMux I__12310 (
            .O(N__51369),
            .I(N__50831));
    ClkMux I__12309 (
            .O(N__51368),
            .I(N__50831));
    ClkMux I__12308 (
            .O(N__51367),
            .I(N__50831));
    ClkMux I__12307 (
            .O(N__51366),
            .I(N__50831));
    ClkMux I__12306 (
            .O(N__51365),
            .I(N__50831));
    ClkMux I__12305 (
            .O(N__51364),
            .I(N__50831));
    ClkMux I__12304 (
            .O(N__51363),
            .I(N__50831));
    ClkMux I__12303 (
            .O(N__51362),
            .I(N__50831));
    ClkMux I__12302 (
            .O(N__51361),
            .I(N__50831));
    ClkMux I__12301 (
            .O(N__51360),
            .I(N__50831));
    ClkMux I__12300 (
            .O(N__51359),
            .I(N__50831));
    ClkMux I__12299 (
            .O(N__51358),
            .I(N__50831));
    ClkMux I__12298 (
            .O(N__51357),
            .I(N__50831));
    ClkMux I__12297 (
            .O(N__51356),
            .I(N__50831));
    ClkMux I__12296 (
            .O(N__51355),
            .I(N__50831));
    ClkMux I__12295 (
            .O(N__51354),
            .I(N__50831));
    ClkMux I__12294 (
            .O(N__51353),
            .I(N__50831));
    ClkMux I__12293 (
            .O(N__51352),
            .I(N__50831));
    ClkMux I__12292 (
            .O(N__51351),
            .I(N__50831));
    ClkMux I__12291 (
            .O(N__51350),
            .I(N__50831));
    ClkMux I__12290 (
            .O(N__51349),
            .I(N__50831));
    ClkMux I__12289 (
            .O(N__51348),
            .I(N__50831));
    ClkMux I__12288 (
            .O(N__51347),
            .I(N__50831));
    ClkMux I__12287 (
            .O(N__51346),
            .I(N__50831));
    ClkMux I__12286 (
            .O(N__51345),
            .I(N__50831));
    ClkMux I__12285 (
            .O(N__51344),
            .I(N__50831));
    ClkMux I__12284 (
            .O(N__51343),
            .I(N__50831));
    ClkMux I__12283 (
            .O(N__51342),
            .I(N__50831));
    ClkMux I__12282 (
            .O(N__51341),
            .I(N__50831));
    ClkMux I__12281 (
            .O(N__51340),
            .I(N__50831));
    ClkMux I__12280 (
            .O(N__51339),
            .I(N__50831));
    ClkMux I__12279 (
            .O(N__51338),
            .I(N__50831));
    ClkMux I__12278 (
            .O(N__51337),
            .I(N__50831));
    ClkMux I__12277 (
            .O(N__51336),
            .I(N__50831));
    ClkMux I__12276 (
            .O(N__51335),
            .I(N__50831));
    ClkMux I__12275 (
            .O(N__51334),
            .I(N__50831));
    ClkMux I__12274 (
            .O(N__51333),
            .I(N__50831));
    ClkMux I__12273 (
            .O(N__51332),
            .I(N__50831));
    ClkMux I__12272 (
            .O(N__51331),
            .I(N__50831));
    ClkMux I__12271 (
            .O(N__51330),
            .I(N__50831));
    ClkMux I__12270 (
            .O(N__51329),
            .I(N__50831));
    ClkMux I__12269 (
            .O(N__51328),
            .I(N__50831));
    ClkMux I__12268 (
            .O(N__51327),
            .I(N__50831));
    ClkMux I__12267 (
            .O(N__51326),
            .I(N__50831));
    ClkMux I__12266 (
            .O(N__51325),
            .I(N__50831));
    ClkMux I__12265 (
            .O(N__51324),
            .I(N__50831));
    ClkMux I__12264 (
            .O(N__51323),
            .I(N__50831));
    ClkMux I__12263 (
            .O(N__51322),
            .I(N__50831));
    ClkMux I__12262 (
            .O(N__51321),
            .I(N__50831));
    ClkMux I__12261 (
            .O(N__51320),
            .I(N__50831));
    ClkMux I__12260 (
            .O(N__51319),
            .I(N__50831));
    ClkMux I__12259 (
            .O(N__51318),
            .I(N__50831));
    ClkMux I__12258 (
            .O(N__51317),
            .I(N__50831));
    ClkMux I__12257 (
            .O(N__51316),
            .I(N__50831));
    ClkMux I__12256 (
            .O(N__51315),
            .I(N__50831));
    ClkMux I__12255 (
            .O(N__51314),
            .I(N__50831));
    ClkMux I__12254 (
            .O(N__51313),
            .I(N__50831));
    ClkMux I__12253 (
            .O(N__51312),
            .I(N__50831));
    ClkMux I__12252 (
            .O(N__51311),
            .I(N__50831));
    ClkMux I__12251 (
            .O(N__51310),
            .I(N__50831));
    ClkMux I__12250 (
            .O(N__51309),
            .I(N__50831));
    ClkMux I__12249 (
            .O(N__51308),
            .I(N__50831));
    ClkMux I__12248 (
            .O(N__51307),
            .I(N__50831));
    ClkMux I__12247 (
            .O(N__51306),
            .I(N__50831));
    GlobalMux I__12246 (
            .O(N__50831),
            .I(N__50828));
    gio2CtrlBuf I__12245 (
            .O(N__50828),
            .I(clk_system_c_g));
    InMux I__12244 (
            .O(N__50825),
            .I(N__50788));
    InMux I__12243 (
            .O(N__50824),
            .I(N__50788));
    InMux I__12242 (
            .O(N__50823),
            .I(N__50788));
    InMux I__12241 (
            .O(N__50822),
            .I(N__50781));
    InMux I__12240 (
            .O(N__50821),
            .I(N__50781));
    InMux I__12239 (
            .O(N__50820),
            .I(N__50781));
    InMux I__12238 (
            .O(N__50819),
            .I(N__50776));
    InMux I__12237 (
            .O(N__50818),
            .I(N__50776));
    InMux I__12236 (
            .O(N__50817),
            .I(N__50773));
    InMux I__12235 (
            .O(N__50816),
            .I(N__50762));
    InMux I__12234 (
            .O(N__50815),
            .I(N__50762));
    InMux I__12233 (
            .O(N__50814),
            .I(N__50762));
    InMux I__12232 (
            .O(N__50813),
            .I(N__50762));
    InMux I__12231 (
            .O(N__50812),
            .I(N__50762));
    InMux I__12230 (
            .O(N__50811),
            .I(N__50755));
    InMux I__12229 (
            .O(N__50810),
            .I(N__50755));
    InMux I__12228 (
            .O(N__50809),
            .I(N__50755));
    InMux I__12227 (
            .O(N__50808),
            .I(N__50746));
    InMux I__12226 (
            .O(N__50807),
            .I(N__50746));
    InMux I__12225 (
            .O(N__50806),
            .I(N__50746));
    InMux I__12224 (
            .O(N__50805),
            .I(N__50746));
    InMux I__12223 (
            .O(N__50804),
            .I(N__50741));
    InMux I__12222 (
            .O(N__50803),
            .I(N__50741));
    InMux I__12221 (
            .O(N__50802),
            .I(N__50738));
    InMux I__12220 (
            .O(N__50801),
            .I(N__50735));
    InMux I__12219 (
            .O(N__50800),
            .I(N__50730));
    InMux I__12218 (
            .O(N__50799),
            .I(N__50730));
    InMux I__12217 (
            .O(N__50798),
            .I(N__50727));
    InMux I__12216 (
            .O(N__50797),
            .I(N__50724));
    InMux I__12215 (
            .O(N__50796),
            .I(N__50721));
    InMux I__12214 (
            .O(N__50795),
            .I(N__50718));
    LocalMux I__12213 (
            .O(N__50788),
            .I(N__50687));
    LocalMux I__12212 (
            .O(N__50781),
            .I(N__50684));
    LocalMux I__12211 (
            .O(N__50776),
            .I(N__50681));
    LocalMux I__12210 (
            .O(N__50773),
            .I(N__50678));
    LocalMux I__12209 (
            .O(N__50762),
            .I(N__50675));
    LocalMux I__12208 (
            .O(N__50755),
            .I(N__50672));
    LocalMux I__12207 (
            .O(N__50746),
            .I(N__50669));
    LocalMux I__12206 (
            .O(N__50741),
            .I(N__50666));
    LocalMux I__12205 (
            .O(N__50738),
            .I(N__50663));
    LocalMux I__12204 (
            .O(N__50735),
            .I(N__50660));
    LocalMux I__12203 (
            .O(N__50730),
            .I(N__50657));
    LocalMux I__12202 (
            .O(N__50727),
            .I(N__50654));
    LocalMux I__12201 (
            .O(N__50724),
            .I(N__50651));
    LocalMux I__12200 (
            .O(N__50721),
            .I(N__50648));
    LocalMux I__12199 (
            .O(N__50718),
            .I(N__50645));
    SRMux I__12198 (
            .O(N__50717),
            .I(N__50558));
    SRMux I__12197 (
            .O(N__50716),
            .I(N__50558));
    SRMux I__12196 (
            .O(N__50715),
            .I(N__50558));
    SRMux I__12195 (
            .O(N__50714),
            .I(N__50558));
    SRMux I__12194 (
            .O(N__50713),
            .I(N__50558));
    SRMux I__12193 (
            .O(N__50712),
            .I(N__50558));
    SRMux I__12192 (
            .O(N__50711),
            .I(N__50558));
    SRMux I__12191 (
            .O(N__50710),
            .I(N__50558));
    SRMux I__12190 (
            .O(N__50709),
            .I(N__50558));
    SRMux I__12189 (
            .O(N__50708),
            .I(N__50558));
    SRMux I__12188 (
            .O(N__50707),
            .I(N__50558));
    SRMux I__12187 (
            .O(N__50706),
            .I(N__50558));
    SRMux I__12186 (
            .O(N__50705),
            .I(N__50558));
    SRMux I__12185 (
            .O(N__50704),
            .I(N__50558));
    SRMux I__12184 (
            .O(N__50703),
            .I(N__50558));
    SRMux I__12183 (
            .O(N__50702),
            .I(N__50558));
    SRMux I__12182 (
            .O(N__50701),
            .I(N__50558));
    SRMux I__12181 (
            .O(N__50700),
            .I(N__50558));
    SRMux I__12180 (
            .O(N__50699),
            .I(N__50558));
    SRMux I__12179 (
            .O(N__50698),
            .I(N__50558));
    SRMux I__12178 (
            .O(N__50697),
            .I(N__50558));
    SRMux I__12177 (
            .O(N__50696),
            .I(N__50558));
    SRMux I__12176 (
            .O(N__50695),
            .I(N__50558));
    SRMux I__12175 (
            .O(N__50694),
            .I(N__50558));
    SRMux I__12174 (
            .O(N__50693),
            .I(N__50558));
    SRMux I__12173 (
            .O(N__50692),
            .I(N__50558));
    SRMux I__12172 (
            .O(N__50691),
            .I(N__50558));
    SRMux I__12171 (
            .O(N__50690),
            .I(N__50558));
    Glb2LocalMux I__12170 (
            .O(N__50687),
            .I(N__50558));
    Glb2LocalMux I__12169 (
            .O(N__50684),
            .I(N__50558));
    Glb2LocalMux I__12168 (
            .O(N__50681),
            .I(N__50558));
    Glb2LocalMux I__12167 (
            .O(N__50678),
            .I(N__50558));
    Glb2LocalMux I__12166 (
            .O(N__50675),
            .I(N__50558));
    Glb2LocalMux I__12165 (
            .O(N__50672),
            .I(N__50558));
    Glb2LocalMux I__12164 (
            .O(N__50669),
            .I(N__50558));
    Glb2LocalMux I__12163 (
            .O(N__50666),
            .I(N__50558));
    Glb2LocalMux I__12162 (
            .O(N__50663),
            .I(N__50558));
    Glb2LocalMux I__12161 (
            .O(N__50660),
            .I(N__50558));
    Glb2LocalMux I__12160 (
            .O(N__50657),
            .I(N__50558));
    Glb2LocalMux I__12159 (
            .O(N__50654),
            .I(N__50558));
    Glb2LocalMux I__12158 (
            .O(N__50651),
            .I(N__50558));
    Glb2LocalMux I__12157 (
            .O(N__50648),
            .I(N__50558));
    Glb2LocalMux I__12156 (
            .O(N__50645),
            .I(N__50558));
    GlobalMux I__12155 (
            .O(N__50558),
            .I(N__50555));
    gio2CtrlBuf I__12154 (
            .O(N__50555),
            .I(N_851_g));
    InMux I__12153 (
            .O(N__50552),
            .I(N__50549));
    LocalMux I__12152 (
            .O(N__50549),
            .I(N__50546));
    Odrv4 I__12151 (
            .O(N__50546),
            .I(\pid_front.O_18 ));
    InMux I__12150 (
            .O(N__50543),
            .I(N__50540));
    LocalMux I__12149 (
            .O(N__50540),
            .I(N__50536));
    InMux I__12148 (
            .O(N__50539),
            .I(N__50533));
    Span4Mux_h I__12147 (
            .O(N__50536),
            .I(N__50530));
    LocalMux I__12146 (
            .O(N__50533),
            .I(N__50527));
    Span4Mux_h I__12145 (
            .O(N__50530),
            .I(N__50524));
    Span4Mux_h I__12144 (
            .O(N__50527),
            .I(N__50520));
    Span4Mux_h I__12143 (
            .O(N__50524),
            .I(N__50517));
    InMux I__12142 (
            .O(N__50523),
            .I(N__50514));
    Span4Mux_h I__12141 (
            .O(N__50520),
            .I(N__50511));
    Odrv4 I__12140 (
            .O(N__50517),
            .I(\pid_front.error_p_regZ0Z_14 ));
    LocalMux I__12139 (
            .O(N__50514),
            .I(\pid_front.error_p_regZ0Z_14 ));
    Odrv4 I__12138 (
            .O(N__50511),
            .I(\pid_front.error_p_regZ0Z_14 ));
    InMux I__12137 (
            .O(N__50504),
            .I(N__50501));
    LocalMux I__12136 (
            .O(N__50501),
            .I(N__50498));
    Odrv4 I__12135 (
            .O(N__50498),
            .I(\pid_front.O_12 ));
    InMux I__12134 (
            .O(N__50495),
            .I(N__50492));
    LocalMux I__12133 (
            .O(N__50492),
            .I(N__50488));
    InMux I__12132 (
            .O(N__50491),
            .I(N__50485));
    Span4Mux_v I__12131 (
            .O(N__50488),
            .I(N__50479));
    LocalMux I__12130 (
            .O(N__50485),
            .I(N__50479));
    InMux I__12129 (
            .O(N__50484),
            .I(N__50476));
    Span4Mux_h I__12128 (
            .O(N__50479),
            .I(N__50473));
    LocalMux I__12127 (
            .O(N__50476),
            .I(\pid_front.error_p_regZ0Z_8 ));
    Odrv4 I__12126 (
            .O(N__50473),
            .I(\pid_front.error_p_regZ0Z_8 ));
    InMux I__12125 (
            .O(N__50468),
            .I(N__50465));
    LocalMux I__12124 (
            .O(N__50465),
            .I(N__50462));
    Odrv4 I__12123 (
            .O(N__50462),
            .I(\pid_front.O_14 ));
    InMux I__12122 (
            .O(N__50459),
            .I(N__50456));
    LocalMux I__12121 (
            .O(N__50456),
            .I(N__50453));
    Span4Mux_v I__12120 (
            .O(N__50453),
            .I(N__50449));
    InMux I__12119 (
            .O(N__50452),
            .I(N__50446));
    Span4Mux_h I__12118 (
            .O(N__50449),
            .I(N__50442));
    LocalMux I__12117 (
            .O(N__50446),
            .I(N__50439));
    InMux I__12116 (
            .O(N__50445),
            .I(N__50436));
    Sp12to4 I__12115 (
            .O(N__50442),
            .I(N__50431));
    Span12Mux_s8_v I__12114 (
            .O(N__50439),
            .I(N__50431));
    LocalMux I__12113 (
            .O(N__50436),
            .I(\pid_front.error_p_regZ0Z_10 ));
    Odrv12 I__12112 (
            .O(N__50431),
            .I(\pid_front.error_p_regZ0Z_10 ));
    InMux I__12111 (
            .O(N__50426),
            .I(N__50423));
    LocalMux I__12110 (
            .O(N__50423),
            .I(N__50420));
    Odrv4 I__12109 (
            .O(N__50420),
            .I(\pid_front.O_11 ));
    InMux I__12108 (
            .O(N__50417),
            .I(N__50413));
    CascadeMux I__12107 (
            .O(N__50416),
            .I(N__50410));
    LocalMux I__12106 (
            .O(N__50413),
            .I(N__50406));
    InMux I__12105 (
            .O(N__50410),
            .I(N__50403));
    InMux I__12104 (
            .O(N__50409),
            .I(N__50400));
    Span12Mux_h I__12103 (
            .O(N__50406),
            .I(N__50395));
    LocalMux I__12102 (
            .O(N__50403),
            .I(N__50395));
    LocalMux I__12101 (
            .O(N__50400),
            .I(\pid_front.error_p_regZ0Z_7 ));
    Odrv12 I__12100 (
            .O(N__50395),
            .I(\pid_front.error_p_regZ0Z_7 ));
    InMux I__12099 (
            .O(N__50390),
            .I(N__50387));
    LocalMux I__12098 (
            .O(N__50387),
            .I(\pid_front.O_7 ));
    InMux I__12097 (
            .O(N__50384),
            .I(N__50381));
    LocalMux I__12096 (
            .O(N__50381),
            .I(N__50378));
    Span4Mux_h I__12095 (
            .O(N__50378),
            .I(N__50374));
    InMux I__12094 (
            .O(N__50377),
            .I(N__50370));
    Span4Mux_h I__12093 (
            .O(N__50374),
            .I(N__50367));
    InMux I__12092 (
            .O(N__50373),
            .I(N__50364));
    LocalMux I__12091 (
            .O(N__50370),
            .I(N__50361));
    Odrv4 I__12090 (
            .O(N__50367),
            .I(\pid_front.error_p_regZ0Z_3 ));
    LocalMux I__12089 (
            .O(N__50364),
            .I(\pid_front.error_p_regZ0Z_3 ));
    Odrv12 I__12088 (
            .O(N__50361),
            .I(\pid_front.error_p_regZ0Z_3 ));
    InMux I__12087 (
            .O(N__50354),
            .I(N__50351));
    LocalMux I__12086 (
            .O(N__50351),
            .I(N__50348));
    Odrv4 I__12085 (
            .O(N__50348),
            .I(\pid_front.O_20 ));
    InMux I__12084 (
            .O(N__50345),
            .I(N__50342));
    LocalMux I__12083 (
            .O(N__50342),
            .I(N__50338));
    InMux I__12082 (
            .O(N__50341),
            .I(N__50335));
    Span4Mux_h I__12081 (
            .O(N__50338),
            .I(N__50329));
    LocalMux I__12080 (
            .O(N__50335),
            .I(N__50329));
    InMux I__12079 (
            .O(N__50334),
            .I(N__50326));
    Span4Mux_h I__12078 (
            .O(N__50329),
            .I(N__50323));
    LocalMux I__12077 (
            .O(N__50326),
            .I(\pid_front.error_p_regZ0Z_16 ));
    Odrv4 I__12076 (
            .O(N__50323),
            .I(\pid_front.error_p_regZ0Z_16 ));
    InMux I__12075 (
            .O(N__50318),
            .I(N__50315));
    LocalMux I__12074 (
            .O(N__50315),
            .I(\pid_front.O_10 ));
    InMux I__12073 (
            .O(N__50312),
            .I(N__50308));
    CascadeMux I__12072 (
            .O(N__50311),
            .I(N__50305));
    LocalMux I__12071 (
            .O(N__50308),
            .I(N__50302));
    InMux I__12070 (
            .O(N__50305),
            .I(N__50299));
    Span4Mux_v I__12069 (
            .O(N__50302),
            .I(N__50296));
    LocalMux I__12068 (
            .O(N__50299),
            .I(N__50293));
    Span4Mux_h I__12067 (
            .O(N__50296),
            .I(N__50289));
    Span4Mux_v I__12066 (
            .O(N__50293),
            .I(N__50286));
    InMux I__12065 (
            .O(N__50292),
            .I(N__50283));
    Span4Mux_h I__12064 (
            .O(N__50289),
            .I(N__50278));
    Span4Mux_h I__12063 (
            .O(N__50286),
            .I(N__50278));
    LocalMux I__12062 (
            .O(N__50283),
            .I(\pid_front.error_p_regZ0Z_6 ));
    Odrv4 I__12061 (
            .O(N__50278),
            .I(\pid_front.error_p_regZ0Z_6 ));
    InMux I__12060 (
            .O(N__50273),
            .I(N__50270));
    LocalMux I__12059 (
            .O(N__50270),
            .I(N__50267));
    Odrv4 I__12058 (
            .O(N__50267),
            .I(\pid_front.O_22 ));
    CascadeMux I__12057 (
            .O(N__50264),
            .I(N__50261));
    InMux I__12056 (
            .O(N__50261),
            .I(N__50258));
    LocalMux I__12055 (
            .O(N__50258),
            .I(N__50255));
    Span4Mux_v I__12054 (
            .O(N__50255),
            .I(N__50252));
    Span4Mux_h I__12053 (
            .O(N__50252),
            .I(N__50248));
    InMux I__12052 (
            .O(N__50251),
            .I(N__50245));
    Sp12to4 I__12051 (
            .O(N__50248),
            .I(N__50239));
    LocalMux I__12050 (
            .O(N__50245),
            .I(N__50239));
    InMux I__12049 (
            .O(N__50244),
            .I(N__50236));
    Span12Mux_s7_v I__12048 (
            .O(N__50239),
            .I(N__50233));
    LocalMux I__12047 (
            .O(N__50236),
            .I(\pid_front.error_p_regZ0Z_18 ));
    Odrv12 I__12046 (
            .O(N__50233),
            .I(\pid_front.error_p_regZ0Z_18 ));
    CascadeMux I__12045 (
            .O(N__50228),
            .I(N__50223));
    CascadeMux I__12044 (
            .O(N__50227),
            .I(N__50219));
    CascadeMux I__12043 (
            .O(N__50226),
            .I(N__50209));
    InMux I__12042 (
            .O(N__50223),
            .I(N__50197));
    InMux I__12041 (
            .O(N__50222),
            .I(N__50197));
    InMux I__12040 (
            .O(N__50219),
            .I(N__50180));
    InMux I__12039 (
            .O(N__50218),
            .I(N__50180));
    InMux I__12038 (
            .O(N__50217),
            .I(N__50180));
    InMux I__12037 (
            .O(N__50216),
            .I(N__50180));
    InMux I__12036 (
            .O(N__50215),
            .I(N__50180));
    InMux I__12035 (
            .O(N__50214),
            .I(N__50180));
    InMux I__12034 (
            .O(N__50213),
            .I(N__50180));
    InMux I__12033 (
            .O(N__50212),
            .I(N__50180));
    InMux I__12032 (
            .O(N__50209),
            .I(N__50160));
    InMux I__12031 (
            .O(N__50208),
            .I(N__50160));
    InMux I__12030 (
            .O(N__50207),
            .I(N__50160));
    InMux I__12029 (
            .O(N__50206),
            .I(N__50160));
    InMux I__12028 (
            .O(N__50205),
            .I(N__50160));
    InMux I__12027 (
            .O(N__50204),
            .I(N__50160));
    InMux I__12026 (
            .O(N__50203),
            .I(N__50160));
    InMux I__12025 (
            .O(N__50202),
            .I(N__50160));
    LocalMux I__12024 (
            .O(N__50197),
            .I(N__50155));
    LocalMux I__12023 (
            .O(N__50180),
            .I(N__50155));
    InMux I__12022 (
            .O(N__50179),
            .I(N__50152));
    InMux I__12021 (
            .O(N__50178),
            .I(N__50147));
    InMux I__12020 (
            .O(N__50177),
            .I(N__50147));
    LocalMux I__12019 (
            .O(N__50160),
            .I(N__50144));
    Span4Mux_v I__12018 (
            .O(N__50155),
            .I(N__50141));
    LocalMux I__12017 (
            .O(N__50152),
            .I(N__50136));
    LocalMux I__12016 (
            .O(N__50147),
            .I(N__50136));
    Span12Mux_s3_h I__12015 (
            .O(N__50144),
            .I(N__50131));
    Sp12to4 I__12014 (
            .O(N__50141),
            .I(N__50131));
    Odrv12 I__12013 (
            .O(N__50136),
            .I(\pid_side.state_RNINK4UZ0Z_1 ));
    Odrv12 I__12012 (
            .O(N__50131),
            .I(\pid_side.state_RNINK4UZ0Z_1 ));
    InMux I__12011 (
            .O(N__50126),
            .I(N__50123));
    LocalMux I__12010 (
            .O(N__50123),
            .I(N__50120));
    Span12Mux_h I__12009 (
            .O(N__50120),
            .I(N__50117));
    Odrv12 I__12008 (
            .O(N__50117),
            .I(\pid_side.O_0_7 ));
    InMux I__12007 (
            .O(N__50114),
            .I(N__50111));
    LocalMux I__12006 (
            .O(N__50111),
            .I(N__50108));
    Span4Mux_h I__12005 (
            .O(N__50108),
            .I(N__50104));
    InMux I__12004 (
            .O(N__50107),
            .I(N__50101));
    Sp12to4 I__12003 (
            .O(N__50104),
            .I(N__50096));
    LocalMux I__12002 (
            .O(N__50101),
            .I(N__50096));
    Span12Mux_v I__12001 (
            .O(N__50096),
            .I(N__50092));
    InMux I__12000 (
            .O(N__50095),
            .I(N__50089));
    Span12Mux_h I__11999 (
            .O(N__50092),
            .I(N__50086));
    LocalMux I__11998 (
            .O(N__50089),
            .I(\pid_side.error_p_regZ0Z_3 ));
    Odrv12 I__11997 (
            .O(N__50086),
            .I(\pid_side.error_p_regZ0Z_3 ));
    InMux I__11996 (
            .O(N__50081),
            .I(N__50078));
    LocalMux I__11995 (
            .O(N__50078),
            .I(N__50075));
    Odrv12 I__11994 (
            .O(N__50075),
            .I(\pid_front.O_4 ));
    InMux I__11993 (
            .O(N__50072),
            .I(N__50069));
    LocalMux I__11992 (
            .O(N__50069),
            .I(N__50066));
    Span4Mux_v I__11991 (
            .O(N__50066),
            .I(N__50063));
    Span4Mux_v I__11990 (
            .O(N__50063),
            .I(N__50060));
    Span4Mux_h I__11989 (
            .O(N__50060),
            .I(N__50056));
    InMux I__11988 (
            .O(N__50059),
            .I(N__50053));
    Odrv4 I__11987 (
            .O(N__50056),
            .I(\pid_front.error_p_regZ0Z_0 ));
    LocalMux I__11986 (
            .O(N__50053),
            .I(\pid_front.error_p_regZ0Z_0 ));
    InMux I__11985 (
            .O(N__50048),
            .I(N__50041));
    CascadeMux I__11984 (
            .O(N__50047),
            .I(N__50036));
    CascadeMux I__11983 (
            .O(N__50046),
            .I(N__50031));
    CascadeMux I__11982 (
            .O(N__50045),
            .I(N__50028));
    CascadeMux I__11981 (
            .O(N__50044),
            .I(N__50024));
    LocalMux I__11980 (
            .O(N__50041),
            .I(N__50016));
    CascadeMux I__11979 (
            .O(N__50040),
            .I(N__50013));
    CascadeMux I__11978 (
            .O(N__50039),
            .I(N__50009));
    InMux I__11977 (
            .O(N__50036),
            .I(N__50006));
    InMux I__11976 (
            .O(N__50035),
            .I(N__50003));
    InMux I__11975 (
            .O(N__50034),
            .I(N__49996));
    InMux I__11974 (
            .O(N__50031),
            .I(N__49996));
    InMux I__11973 (
            .O(N__50028),
            .I(N__49996));
    InMux I__11972 (
            .O(N__50027),
            .I(N__49989));
    InMux I__11971 (
            .O(N__50024),
            .I(N__49989));
    InMux I__11970 (
            .O(N__50023),
            .I(N__49989));
    CascadeMux I__11969 (
            .O(N__50022),
            .I(N__49986));
    CascadeMux I__11968 (
            .O(N__50021),
            .I(N__49982));
    CascadeMux I__11967 (
            .O(N__50020),
            .I(N__49979));
    InMux I__11966 (
            .O(N__50019),
            .I(N__49971));
    Span4Mux_h I__11965 (
            .O(N__50016),
            .I(N__49968));
    InMux I__11964 (
            .O(N__50013),
            .I(N__49963));
    InMux I__11963 (
            .O(N__50012),
            .I(N__49963));
    InMux I__11962 (
            .O(N__50009),
            .I(N__49960));
    LocalMux I__11961 (
            .O(N__50006),
            .I(N__49957));
    LocalMux I__11960 (
            .O(N__50003),
            .I(N__49950));
    LocalMux I__11959 (
            .O(N__49996),
            .I(N__49950));
    LocalMux I__11958 (
            .O(N__49989),
            .I(N__49950));
    InMux I__11957 (
            .O(N__49986),
            .I(N__49945));
    InMux I__11956 (
            .O(N__49985),
            .I(N__49945));
    InMux I__11955 (
            .O(N__49982),
            .I(N__49940));
    InMux I__11954 (
            .O(N__49979),
            .I(N__49940));
    CascadeMux I__11953 (
            .O(N__49978),
            .I(N__49937));
    CascadeMux I__11952 (
            .O(N__49977),
            .I(N__49934));
    CascadeMux I__11951 (
            .O(N__49976),
            .I(N__49931));
    CascadeMux I__11950 (
            .O(N__49975),
            .I(N__49927));
    InMux I__11949 (
            .O(N__49974),
            .I(N__49923));
    LocalMux I__11948 (
            .O(N__49971),
            .I(N__49918));
    Span4Mux_h I__11947 (
            .O(N__49968),
            .I(N__49918));
    LocalMux I__11946 (
            .O(N__49963),
            .I(N__49915));
    LocalMux I__11945 (
            .O(N__49960),
            .I(N__49912));
    Span4Mux_v I__11944 (
            .O(N__49957),
            .I(N__49903));
    Span4Mux_v I__11943 (
            .O(N__49950),
            .I(N__49903));
    LocalMux I__11942 (
            .O(N__49945),
            .I(N__49903));
    LocalMux I__11941 (
            .O(N__49940),
            .I(N__49903));
    InMux I__11940 (
            .O(N__49937),
            .I(N__49900));
    InMux I__11939 (
            .O(N__49934),
            .I(N__49891));
    InMux I__11938 (
            .O(N__49931),
            .I(N__49891));
    InMux I__11937 (
            .O(N__49930),
            .I(N__49891));
    InMux I__11936 (
            .O(N__49927),
            .I(N__49891));
    InMux I__11935 (
            .O(N__49926),
            .I(N__49888));
    LocalMux I__11934 (
            .O(N__49923),
            .I(N__49881));
    Span4Mux_h I__11933 (
            .O(N__49918),
            .I(N__49881));
    Span4Mux_h I__11932 (
            .O(N__49915),
            .I(N__49881));
    Odrv12 I__11931 (
            .O(N__49912),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__11930 (
            .O(N__49903),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__11929 (
            .O(N__49900),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__11928 (
            .O(N__49891),
            .I(\pid_side.stateZ0Z_0 ));
    LocalMux I__11927 (
            .O(N__49888),
            .I(\pid_side.stateZ0Z_0 ));
    Odrv4 I__11926 (
            .O(N__49881),
            .I(\pid_side.stateZ0Z_0 ));
    InMux I__11925 (
            .O(N__49868),
            .I(N__49864));
    InMux I__11924 (
            .O(N__49867),
            .I(N__49861));
    LocalMux I__11923 (
            .O(N__49864),
            .I(N__49858));
    LocalMux I__11922 (
            .O(N__49861),
            .I(N__49855));
    Span4Mux_v I__11921 (
            .O(N__49858),
            .I(N__49851));
    Span4Mux_v I__11920 (
            .O(N__49855),
            .I(N__49848));
    InMux I__11919 (
            .O(N__49854),
            .I(N__49845));
    Sp12to4 I__11918 (
            .O(N__49851),
            .I(N__49842));
    Odrv4 I__11917 (
            .O(N__49848),
            .I(\pid_side.error_p_regZ0Z_1 ));
    LocalMux I__11916 (
            .O(N__49845),
            .I(\pid_side.error_p_regZ0Z_1 ));
    Odrv12 I__11915 (
            .O(N__49842),
            .I(\pid_side.error_p_regZ0Z_1 ));
    CascadeMux I__11914 (
            .O(N__49835),
            .I(N__49832));
    InMux I__11913 (
            .O(N__49832),
            .I(N__49827));
    InMux I__11912 (
            .O(N__49831),
            .I(N__49822));
    InMux I__11911 (
            .O(N__49830),
            .I(N__49822));
    LocalMux I__11910 (
            .O(N__49827),
            .I(N__49818));
    LocalMux I__11909 (
            .O(N__49822),
            .I(N__49815));
    InMux I__11908 (
            .O(N__49821),
            .I(N__49812));
    Span4Mux_v I__11907 (
            .O(N__49818),
            .I(N__49807));
    Span4Mux_h I__11906 (
            .O(N__49815),
            .I(N__49807));
    LocalMux I__11905 (
            .O(N__49812),
            .I(N__49802));
    Span4Mux_h I__11904 (
            .O(N__49807),
            .I(N__49802));
    Odrv4 I__11903 (
            .O(N__49802),
            .I(\pid_side.pid_preregZ0Z_1 ));
    CascadeMux I__11902 (
            .O(N__49799),
            .I(N__49792));
    CascadeMux I__11901 (
            .O(N__49798),
            .I(N__49789));
    CascadeMux I__11900 (
            .O(N__49797),
            .I(N__49786));
    CascadeMux I__11899 (
            .O(N__49796),
            .I(N__49761));
    InMux I__11898 (
            .O(N__49795),
            .I(N__49743));
    InMux I__11897 (
            .O(N__49792),
            .I(N__49738));
    InMux I__11896 (
            .O(N__49789),
            .I(N__49738));
    InMux I__11895 (
            .O(N__49786),
            .I(N__49729));
    InMux I__11894 (
            .O(N__49785),
            .I(N__49729));
    InMux I__11893 (
            .O(N__49784),
            .I(N__49729));
    InMux I__11892 (
            .O(N__49783),
            .I(N__49729));
    InMux I__11891 (
            .O(N__49782),
            .I(N__49726));
    InMux I__11890 (
            .O(N__49781),
            .I(N__49723));
    InMux I__11889 (
            .O(N__49780),
            .I(N__49718));
    InMux I__11888 (
            .O(N__49779),
            .I(N__49718));
    InMux I__11887 (
            .O(N__49778),
            .I(N__49715));
    InMux I__11886 (
            .O(N__49777),
            .I(N__49712));
    InMux I__11885 (
            .O(N__49776),
            .I(N__49709));
    InMux I__11884 (
            .O(N__49775),
            .I(N__49704));
    InMux I__11883 (
            .O(N__49774),
            .I(N__49704));
    InMux I__11882 (
            .O(N__49773),
            .I(N__49701));
    InMux I__11881 (
            .O(N__49772),
            .I(N__49698));
    InMux I__11880 (
            .O(N__49771),
            .I(N__49695));
    InMux I__11879 (
            .O(N__49770),
            .I(N__49692));
    InMux I__11878 (
            .O(N__49769),
            .I(N__49689));
    InMux I__11877 (
            .O(N__49768),
            .I(N__49686));
    InMux I__11876 (
            .O(N__49767),
            .I(N__49683));
    InMux I__11875 (
            .O(N__49766),
            .I(N__49678));
    InMux I__11874 (
            .O(N__49765),
            .I(N__49678));
    InMux I__11873 (
            .O(N__49764),
            .I(N__49675));
    InMux I__11872 (
            .O(N__49761),
            .I(N__49672));
    InMux I__11871 (
            .O(N__49760),
            .I(N__49669));
    InMux I__11870 (
            .O(N__49759),
            .I(N__49666));
    InMux I__11869 (
            .O(N__49758),
            .I(N__49663));
    InMux I__11868 (
            .O(N__49757),
            .I(N__49658));
    InMux I__11867 (
            .O(N__49756),
            .I(N__49658));
    InMux I__11866 (
            .O(N__49755),
            .I(N__49655));
    InMux I__11865 (
            .O(N__49754),
            .I(N__49652));
    InMux I__11864 (
            .O(N__49753),
            .I(N__49649));
    InMux I__11863 (
            .O(N__49752),
            .I(N__49646));
    InMux I__11862 (
            .O(N__49751),
            .I(N__49643));
    InMux I__11861 (
            .O(N__49750),
            .I(N__49638));
    InMux I__11860 (
            .O(N__49749),
            .I(N__49638));
    InMux I__11859 (
            .O(N__49748),
            .I(N__49635));
    InMux I__11858 (
            .O(N__49747),
            .I(N__49632));
    InMux I__11857 (
            .O(N__49746),
            .I(N__49629));
    LocalMux I__11856 (
            .O(N__49743),
            .I(N__49495));
    LocalMux I__11855 (
            .O(N__49738),
            .I(N__49492));
    LocalMux I__11854 (
            .O(N__49729),
            .I(N__49489));
    LocalMux I__11853 (
            .O(N__49726),
            .I(N__49486));
    LocalMux I__11852 (
            .O(N__49723),
            .I(N__49483));
    LocalMux I__11851 (
            .O(N__49718),
            .I(N__49480));
    LocalMux I__11850 (
            .O(N__49715),
            .I(N__49477));
    LocalMux I__11849 (
            .O(N__49712),
            .I(N__49474));
    LocalMux I__11848 (
            .O(N__49709),
            .I(N__49471));
    LocalMux I__11847 (
            .O(N__49704),
            .I(N__49468));
    LocalMux I__11846 (
            .O(N__49701),
            .I(N__49465));
    LocalMux I__11845 (
            .O(N__49698),
            .I(N__49462));
    LocalMux I__11844 (
            .O(N__49695),
            .I(N__49459));
    LocalMux I__11843 (
            .O(N__49692),
            .I(N__49456));
    LocalMux I__11842 (
            .O(N__49689),
            .I(N__49453));
    LocalMux I__11841 (
            .O(N__49686),
            .I(N__49450));
    LocalMux I__11840 (
            .O(N__49683),
            .I(N__49447));
    LocalMux I__11839 (
            .O(N__49678),
            .I(N__49444));
    LocalMux I__11838 (
            .O(N__49675),
            .I(N__49441));
    LocalMux I__11837 (
            .O(N__49672),
            .I(N__49438));
    LocalMux I__11836 (
            .O(N__49669),
            .I(N__49435));
    LocalMux I__11835 (
            .O(N__49666),
            .I(N__49432));
    LocalMux I__11834 (
            .O(N__49663),
            .I(N__49429));
    LocalMux I__11833 (
            .O(N__49658),
            .I(N__49426));
    LocalMux I__11832 (
            .O(N__49655),
            .I(N__49423));
    LocalMux I__11831 (
            .O(N__49652),
            .I(N__49420));
    LocalMux I__11830 (
            .O(N__49649),
            .I(N__49417));
    LocalMux I__11829 (
            .O(N__49646),
            .I(N__49414));
    LocalMux I__11828 (
            .O(N__49643),
            .I(N__49411));
    LocalMux I__11827 (
            .O(N__49638),
            .I(N__49408));
    LocalMux I__11826 (
            .O(N__49635),
            .I(N__49405));
    LocalMux I__11825 (
            .O(N__49632),
            .I(N__49402));
    LocalMux I__11824 (
            .O(N__49629),
            .I(N__49399));
    SRMux I__11823 (
            .O(N__49628),
            .I(N__49070));
    SRMux I__11822 (
            .O(N__49627),
            .I(N__49070));
    SRMux I__11821 (
            .O(N__49626),
            .I(N__49070));
    SRMux I__11820 (
            .O(N__49625),
            .I(N__49070));
    SRMux I__11819 (
            .O(N__49624),
            .I(N__49070));
    SRMux I__11818 (
            .O(N__49623),
            .I(N__49070));
    SRMux I__11817 (
            .O(N__49622),
            .I(N__49070));
    SRMux I__11816 (
            .O(N__49621),
            .I(N__49070));
    SRMux I__11815 (
            .O(N__49620),
            .I(N__49070));
    SRMux I__11814 (
            .O(N__49619),
            .I(N__49070));
    SRMux I__11813 (
            .O(N__49618),
            .I(N__49070));
    SRMux I__11812 (
            .O(N__49617),
            .I(N__49070));
    SRMux I__11811 (
            .O(N__49616),
            .I(N__49070));
    SRMux I__11810 (
            .O(N__49615),
            .I(N__49070));
    SRMux I__11809 (
            .O(N__49614),
            .I(N__49070));
    SRMux I__11808 (
            .O(N__49613),
            .I(N__49070));
    SRMux I__11807 (
            .O(N__49612),
            .I(N__49070));
    SRMux I__11806 (
            .O(N__49611),
            .I(N__49070));
    SRMux I__11805 (
            .O(N__49610),
            .I(N__49070));
    SRMux I__11804 (
            .O(N__49609),
            .I(N__49070));
    SRMux I__11803 (
            .O(N__49608),
            .I(N__49070));
    SRMux I__11802 (
            .O(N__49607),
            .I(N__49070));
    SRMux I__11801 (
            .O(N__49606),
            .I(N__49070));
    SRMux I__11800 (
            .O(N__49605),
            .I(N__49070));
    SRMux I__11799 (
            .O(N__49604),
            .I(N__49070));
    SRMux I__11798 (
            .O(N__49603),
            .I(N__49070));
    SRMux I__11797 (
            .O(N__49602),
            .I(N__49070));
    SRMux I__11796 (
            .O(N__49601),
            .I(N__49070));
    SRMux I__11795 (
            .O(N__49600),
            .I(N__49070));
    SRMux I__11794 (
            .O(N__49599),
            .I(N__49070));
    SRMux I__11793 (
            .O(N__49598),
            .I(N__49070));
    SRMux I__11792 (
            .O(N__49597),
            .I(N__49070));
    SRMux I__11791 (
            .O(N__49596),
            .I(N__49070));
    SRMux I__11790 (
            .O(N__49595),
            .I(N__49070));
    SRMux I__11789 (
            .O(N__49594),
            .I(N__49070));
    SRMux I__11788 (
            .O(N__49593),
            .I(N__49070));
    SRMux I__11787 (
            .O(N__49592),
            .I(N__49070));
    SRMux I__11786 (
            .O(N__49591),
            .I(N__49070));
    SRMux I__11785 (
            .O(N__49590),
            .I(N__49070));
    SRMux I__11784 (
            .O(N__49589),
            .I(N__49070));
    SRMux I__11783 (
            .O(N__49588),
            .I(N__49070));
    SRMux I__11782 (
            .O(N__49587),
            .I(N__49070));
    SRMux I__11781 (
            .O(N__49586),
            .I(N__49070));
    SRMux I__11780 (
            .O(N__49585),
            .I(N__49070));
    SRMux I__11779 (
            .O(N__49584),
            .I(N__49070));
    SRMux I__11778 (
            .O(N__49583),
            .I(N__49070));
    SRMux I__11777 (
            .O(N__49582),
            .I(N__49070));
    SRMux I__11776 (
            .O(N__49581),
            .I(N__49070));
    SRMux I__11775 (
            .O(N__49580),
            .I(N__49070));
    SRMux I__11774 (
            .O(N__49579),
            .I(N__49070));
    SRMux I__11773 (
            .O(N__49578),
            .I(N__49070));
    SRMux I__11772 (
            .O(N__49577),
            .I(N__49070));
    SRMux I__11771 (
            .O(N__49576),
            .I(N__49070));
    SRMux I__11770 (
            .O(N__49575),
            .I(N__49070));
    SRMux I__11769 (
            .O(N__49574),
            .I(N__49070));
    SRMux I__11768 (
            .O(N__49573),
            .I(N__49070));
    SRMux I__11767 (
            .O(N__49572),
            .I(N__49070));
    SRMux I__11766 (
            .O(N__49571),
            .I(N__49070));
    SRMux I__11765 (
            .O(N__49570),
            .I(N__49070));
    SRMux I__11764 (
            .O(N__49569),
            .I(N__49070));
    SRMux I__11763 (
            .O(N__49568),
            .I(N__49070));
    SRMux I__11762 (
            .O(N__49567),
            .I(N__49070));
    SRMux I__11761 (
            .O(N__49566),
            .I(N__49070));
    SRMux I__11760 (
            .O(N__49565),
            .I(N__49070));
    SRMux I__11759 (
            .O(N__49564),
            .I(N__49070));
    SRMux I__11758 (
            .O(N__49563),
            .I(N__49070));
    SRMux I__11757 (
            .O(N__49562),
            .I(N__49070));
    SRMux I__11756 (
            .O(N__49561),
            .I(N__49070));
    SRMux I__11755 (
            .O(N__49560),
            .I(N__49070));
    SRMux I__11754 (
            .O(N__49559),
            .I(N__49070));
    SRMux I__11753 (
            .O(N__49558),
            .I(N__49070));
    SRMux I__11752 (
            .O(N__49557),
            .I(N__49070));
    SRMux I__11751 (
            .O(N__49556),
            .I(N__49070));
    SRMux I__11750 (
            .O(N__49555),
            .I(N__49070));
    SRMux I__11749 (
            .O(N__49554),
            .I(N__49070));
    SRMux I__11748 (
            .O(N__49553),
            .I(N__49070));
    SRMux I__11747 (
            .O(N__49552),
            .I(N__49070));
    SRMux I__11746 (
            .O(N__49551),
            .I(N__49070));
    SRMux I__11745 (
            .O(N__49550),
            .I(N__49070));
    SRMux I__11744 (
            .O(N__49549),
            .I(N__49070));
    SRMux I__11743 (
            .O(N__49548),
            .I(N__49070));
    SRMux I__11742 (
            .O(N__49547),
            .I(N__49070));
    SRMux I__11741 (
            .O(N__49546),
            .I(N__49070));
    SRMux I__11740 (
            .O(N__49545),
            .I(N__49070));
    SRMux I__11739 (
            .O(N__49544),
            .I(N__49070));
    SRMux I__11738 (
            .O(N__49543),
            .I(N__49070));
    SRMux I__11737 (
            .O(N__49542),
            .I(N__49070));
    SRMux I__11736 (
            .O(N__49541),
            .I(N__49070));
    SRMux I__11735 (
            .O(N__49540),
            .I(N__49070));
    SRMux I__11734 (
            .O(N__49539),
            .I(N__49070));
    SRMux I__11733 (
            .O(N__49538),
            .I(N__49070));
    SRMux I__11732 (
            .O(N__49537),
            .I(N__49070));
    SRMux I__11731 (
            .O(N__49536),
            .I(N__49070));
    SRMux I__11730 (
            .O(N__49535),
            .I(N__49070));
    SRMux I__11729 (
            .O(N__49534),
            .I(N__49070));
    SRMux I__11728 (
            .O(N__49533),
            .I(N__49070));
    SRMux I__11727 (
            .O(N__49532),
            .I(N__49070));
    SRMux I__11726 (
            .O(N__49531),
            .I(N__49070));
    SRMux I__11725 (
            .O(N__49530),
            .I(N__49070));
    SRMux I__11724 (
            .O(N__49529),
            .I(N__49070));
    SRMux I__11723 (
            .O(N__49528),
            .I(N__49070));
    SRMux I__11722 (
            .O(N__49527),
            .I(N__49070));
    SRMux I__11721 (
            .O(N__49526),
            .I(N__49070));
    SRMux I__11720 (
            .O(N__49525),
            .I(N__49070));
    SRMux I__11719 (
            .O(N__49524),
            .I(N__49070));
    SRMux I__11718 (
            .O(N__49523),
            .I(N__49070));
    SRMux I__11717 (
            .O(N__49522),
            .I(N__49070));
    SRMux I__11716 (
            .O(N__49521),
            .I(N__49070));
    SRMux I__11715 (
            .O(N__49520),
            .I(N__49070));
    SRMux I__11714 (
            .O(N__49519),
            .I(N__49070));
    SRMux I__11713 (
            .O(N__49518),
            .I(N__49070));
    SRMux I__11712 (
            .O(N__49517),
            .I(N__49070));
    SRMux I__11711 (
            .O(N__49516),
            .I(N__49070));
    SRMux I__11710 (
            .O(N__49515),
            .I(N__49070));
    SRMux I__11709 (
            .O(N__49514),
            .I(N__49070));
    SRMux I__11708 (
            .O(N__49513),
            .I(N__49070));
    SRMux I__11707 (
            .O(N__49512),
            .I(N__49070));
    SRMux I__11706 (
            .O(N__49511),
            .I(N__49070));
    SRMux I__11705 (
            .O(N__49510),
            .I(N__49070));
    SRMux I__11704 (
            .O(N__49509),
            .I(N__49070));
    SRMux I__11703 (
            .O(N__49508),
            .I(N__49070));
    SRMux I__11702 (
            .O(N__49507),
            .I(N__49070));
    SRMux I__11701 (
            .O(N__49506),
            .I(N__49070));
    SRMux I__11700 (
            .O(N__49505),
            .I(N__49070));
    SRMux I__11699 (
            .O(N__49504),
            .I(N__49070));
    SRMux I__11698 (
            .O(N__49503),
            .I(N__49070));
    SRMux I__11697 (
            .O(N__49502),
            .I(N__49070));
    SRMux I__11696 (
            .O(N__49501),
            .I(N__49070));
    SRMux I__11695 (
            .O(N__49500),
            .I(N__49070));
    SRMux I__11694 (
            .O(N__49499),
            .I(N__49070));
    SRMux I__11693 (
            .O(N__49498),
            .I(N__49070));
    Glb2LocalMux I__11692 (
            .O(N__49495),
            .I(N__49070));
    Glb2LocalMux I__11691 (
            .O(N__49492),
            .I(N__49070));
    Glb2LocalMux I__11690 (
            .O(N__49489),
            .I(N__49070));
    Glb2LocalMux I__11689 (
            .O(N__49486),
            .I(N__49070));
    Glb2LocalMux I__11688 (
            .O(N__49483),
            .I(N__49070));
    Glb2LocalMux I__11687 (
            .O(N__49480),
            .I(N__49070));
    Glb2LocalMux I__11686 (
            .O(N__49477),
            .I(N__49070));
    Glb2LocalMux I__11685 (
            .O(N__49474),
            .I(N__49070));
    Glb2LocalMux I__11684 (
            .O(N__49471),
            .I(N__49070));
    Glb2LocalMux I__11683 (
            .O(N__49468),
            .I(N__49070));
    Glb2LocalMux I__11682 (
            .O(N__49465),
            .I(N__49070));
    Glb2LocalMux I__11681 (
            .O(N__49462),
            .I(N__49070));
    Glb2LocalMux I__11680 (
            .O(N__49459),
            .I(N__49070));
    Glb2LocalMux I__11679 (
            .O(N__49456),
            .I(N__49070));
    Glb2LocalMux I__11678 (
            .O(N__49453),
            .I(N__49070));
    Glb2LocalMux I__11677 (
            .O(N__49450),
            .I(N__49070));
    Glb2LocalMux I__11676 (
            .O(N__49447),
            .I(N__49070));
    Glb2LocalMux I__11675 (
            .O(N__49444),
            .I(N__49070));
    Glb2LocalMux I__11674 (
            .O(N__49441),
            .I(N__49070));
    Glb2LocalMux I__11673 (
            .O(N__49438),
            .I(N__49070));
    Glb2LocalMux I__11672 (
            .O(N__49435),
            .I(N__49070));
    Glb2LocalMux I__11671 (
            .O(N__49432),
            .I(N__49070));
    Glb2LocalMux I__11670 (
            .O(N__49429),
            .I(N__49070));
    Glb2LocalMux I__11669 (
            .O(N__49426),
            .I(N__49070));
    Glb2LocalMux I__11668 (
            .O(N__49423),
            .I(N__49070));
    Glb2LocalMux I__11667 (
            .O(N__49420),
            .I(N__49070));
    Glb2LocalMux I__11666 (
            .O(N__49417),
            .I(N__49070));
    Glb2LocalMux I__11665 (
            .O(N__49414),
            .I(N__49070));
    Glb2LocalMux I__11664 (
            .O(N__49411),
            .I(N__49070));
    Glb2LocalMux I__11663 (
            .O(N__49408),
            .I(N__49070));
    Glb2LocalMux I__11662 (
            .O(N__49405),
            .I(N__49070));
    Glb2LocalMux I__11661 (
            .O(N__49402),
            .I(N__49070));
    Glb2LocalMux I__11660 (
            .O(N__49399),
            .I(N__49070));
    GlobalMux I__11659 (
            .O(N__49070),
            .I(N__49067));
    gio2CtrlBuf I__11658 (
            .O(N__49067),
            .I(reset_system_g));
    InMux I__11657 (
            .O(N__49064),
            .I(N__49061));
    LocalMux I__11656 (
            .O(N__49061),
            .I(N__49058));
    Span4Mux_v I__11655 (
            .O(N__49058),
            .I(N__49055));
    Span4Mux_h I__11654 (
            .O(N__49055),
            .I(N__49052));
    Span4Mux_h I__11653 (
            .O(N__49052),
            .I(N__49049));
    Odrv4 I__11652 (
            .O(N__49049),
            .I(\pid_front.state_ns_0 ));
    InMux I__11651 (
            .O(N__49046),
            .I(N__49043));
    LocalMux I__11650 (
            .O(N__49043),
            .I(N__49039));
    InMux I__11649 (
            .O(N__49042),
            .I(N__49035));
    Span4Mux_v I__11648 (
            .O(N__49039),
            .I(N__49030));
    InMux I__11647 (
            .O(N__49038),
            .I(N__49027));
    LocalMux I__11646 (
            .O(N__49035),
            .I(N__49019));
    IoInMux I__11645 (
            .O(N__49034),
            .I(N__49016));
    InMux I__11644 (
            .O(N__49033),
            .I(N__49011));
    Span4Mux_h I__11643 (
            .O(N__49030),
            .I(N__49005));
    LocalMux I__11642 (
            .O(N__49027),
            .I(N__49005));
    InMux I__11641 (
            .O(N__49026),
            .I(N__49000));
    InMux I__11640 (
            .O(N__49025),
            .I(N__49000));
    InMux I__11639 (
            .O(N__49024),
            .I(N__48997));
    InMux I__11638 (
            .O(N__49023),
            .I(N__48994));
    InMux I__11637 (
            .O(N__49022),
            .I(N__48990));
    Span4Mux_v I__11636 (
            .O(N__49019),
            .I(N__48984));
    LocalMux I__11635 (
            .O(N__49016),
            .I(N__48981));
    InMux I__11634 (
            .O(N__49015),
            .I(N__48974));
    InMux I__11633 (
            .O(N__49014),
            .I(N__48971));
    LocalMux I__11632 (
            .O(N__49011),
            .I(N__48962));
    InMux I__11631 (
            .O(N__49010),
            .I(N__48958));
    Span4Mux_v I__11630 (
            .O(N__49005),
            .I(N__48953));
    LocalMux I__11629 (
            .O(N__49000),
            .I(N__48946));
    LocalMux I__11628 (
            .O(N__48997),
            .I(N__48946));
    LocalMux I__11627 (
            .O(N__48994),
            .I(N__48946));
    InMux I__11626 (
            .O(N__48993),
            .I(N__48943));
    LocalMux I__11625 (
            .O(N__48990),
            .I(N__48940));
    InMux I__11624 (
            .O(N__48989),
            .I(N__48933));
    InMux I__11623 (
            .O(N__48988),
            .I(N__48933));
    InMux I__11622 (
            .O(N__48987),
            .I(N__48933));
    Span4Mux_v I__11621 (
            .O(N__48984),
            .I(N__48930));
    Span4Mux_s1_v I__11620 (
            .O(N__48981),
            .I(N__48927));
    InMux I__11619 (
            .O(N__48980),
            .I(N__48922));
    InMux I__11618 (
            .O(N__48979),
            .I(N__48922));
    InMux I__11617 (
            .O(N__48978),
            .I(N__48919));
    InMux I__11616 (
            .O(N__48977),
            .I(N__48916));
    LocalMux I__11615 (
            .O(N__48974),
            .I(N__48911));
    LocalMux I__11614 (
            .O(N__48971),
            .I(N__48911));
    InMux I__11613 (
            .O(N__48970),
            .I(N__48905));
    InMux I__11612 (
            .O(N__48969),
            .I(N__48905));
    InMux I__11611 (
            .O(N__48968),
            .I(N__48900));
    InMux I__11610 (
            .O(N__48967),
            .I(N__48900));
    InMux I__11609 (
            .O(N__48966),
            .I(N__48895));
    InMux I__11608 (
            .O(N__48965),
            .I(N__48895));
    Span4Mux_h I__11607 (
            .O(N__48962),
            .I(N__48892));
    InMux I__11606 (
            .O(N__48961),
            .I(N__48889));
    LocalMux I__11605 (
            .O(N__48958),
            .I(N__48886));
    InMux I__11604 (
            .O(N__48957),
            .I(N__48881));
    InMux I__11603 (
            .O(N__48956),
            .I(N__48881));
    Span4Mux_h I__11602 (
            .O(N__48953),
            .I(N__48876));
    Span4Mux_v I__11601 (
            .O(N__48946),
            .I(N__48876));
    LocalMux I__11600 (
            .O(N__48943),
            .I(N__48869));
    Span4Mux_v I__11599 (
            .O(N__48940),
            .I(N__48869));
    LocalMux I__11598 (
            .O(N__48933),
            .I(N__48869));
    Span4Mux_v I__11597 (
            .O(N__48930),
            .I(N__48864));
    Span4Mux_v I__11596 (
            .O(N__48927),
            .I(N__48864));
    LocalMux I__11595 (
            .O(N__48922),
            .I(N__48859));
    LocalMux I__11594 (
            .O(N__48919),
            .I(N__48859));
    LocalMux I__11593 (
            .O(N__48916),
            .I(N__48856));
    Span4Mux_v I__11592 (
            .O(N__48911),
            .I(N__48853));
    InMux I__11591 (
            .O(N__48910),
            .I(N__48850));
    LocalMux I__11590 (
            .O(N__48905),
            .I(N__48839));
    LocalMux I__11589 (
            .O(N__48900),
            .I(N__48839));
    LocalMux I__11588 (
            .O(N__48895),
            .I(N__48839));
    Sp12to4 I__11587 (
            .O(N__48892),
            .I(N__48839));
    LocalMux I__11586 (
            .O(N__48889),
            .I(N__48839));
    Span4Mux_v I__11585 (
            .O(N__48886),
            .I(N__48836));
    LocalMux I__11584 (
            .O(N__48881),
            .I(N__48831));
    Span4Mux_v I__11583 (
            .O(N__48876),
            .I(N__48831));
    Span4Mux_v I__11582 (
            .O(N__48869),
            .I(N__48826));
    Span4Mux_h I__11581 (
            .O(N__48864),
            .I(N__48826));
    Span4Mux_v I__11580 (
            .O(N__48859),
            .I(N__48823));
    Span4Mux_h I__11579 (
            .O(N__48856),
            .I(N__48820));
    Span4Mux_v I__11578 (
            .O(N__48853),
            .I(N__48817));
    LocalMux I__11577 (
            .O(N__48850),
            .I(N__48812));
    Span12Mux_v I__11576 (
            .O(N__48839),
            .I(N__48812));
    Span4Mux_v I__11575 (
            .O(N__48836),
            .I(N__48805));
    Span4Mux_v I__11574 (
            .O(N__48831),
            .I(N__48805));
    Span4Mux_h I__11573 (
            .O(N__48826),
            .I(N__48805));
    Odrv4 I__11572 (
            .O(N__48823),
            .I(reset_system));
    Odrv4 I__11571 (
            .O(N__48820),
            .I(reset_system));
    Odrv4 I__11570 (
            .O(N__48817),
            .I(reset_system));
    Odrv12 I__11569 (
            .O(N__48812),
            .I(reset_system));
    Odrv4 I__11568 (
            .O(N__48805),
            .I(reset_system));
    InMux I__11567 (
            .O(N__48794),
            .I(N__48791));
    LocalMux I__11566 (
            .O(N__48791),
            .I(N__48788));
    Odrv12 I__11565 (
            .O(N__48788),
            .I(\pid_front.O_5 ));
    InMux I__11564 (
            .O(N__48785),
            .I(N__48781));
    InMux I__11563 (
            .O(N__48784),
            .I(N__48778));
    LocalMux I__11562 (
            .O(N__48781),
            .I(N__48775));
    LocalMux I__11561 (
            .O(N__48778),
            .I(N__48771));
    Span12Mux_v I__11560 (
            .O(N__48775),
            .I(N__48768));
    InMux I__11559 (
            .O(N__48774),
            .I(N__48765));
    Span4Mux_h I__11558 (
            .O(N__48771),
            .I(N__48762));
    Odrv12 I__11557 (
            .O(N__48768),
            .I(\pid_front.error_p_regZ0Z_1 ));
    LocalMux I__11556 (
            .O(N__48765),
            .I(\pid_front.error_p_regZ0Z_1 ));
    Odrv4 I__11555 (
            .O(N__48762),
            .I(\pid_front.error_p_regZ0Z_1 ));
    InMux I__11554 (
            .O(N__48755),
            .I(N__48752));
    LocalMux I__11553 (
            .O(N__48752),
            .I(N__48749));
    Span4Mux_h I__11552 (
            .O(N__48749),
            .I(N__48746));
    Odrv4 I__11551 (
            .O(N__48746),
            .I(\pid_front.O_13 ));
    InMux I__11550 (
            .O(N__48743),
            .I(N__48740));
    LocalMux I__11549 (
            .O(N__48740),
            .I(N__48735));
    InMux I__11548 (
            .O(N__48739),
            .I(N__48732));
    InMux I__11547 (
            .O(N__48738),
            .I(N__48729));
    Span12Mux_h I__11546 (
            .O(N__48735),
            .I(N__48724));
    LocalMux I__11545 (
            .O(N__48732),
            .I(N__48724));
    LocalMux I__11544 (
            .O(N__48729),
            .I(\pid_front.error_p_regZ0Z_9 ));
    Odrv12 I__11543 (
            .O(N__48724),
            .I(\pid_front.error_p_regZ0Z_9 ));
    InMux I__11542 (
            .O(N__48719),
            .I(N__48716));
    LocalMux I__11541 (
            .O(N__48716),
            .I(N__48713));
    Odrv4 I__11540 (
            .O(N__48713),
            .I(\pid_front.O_6 ));
    InMux I__11539 (
            .O(N__48710),
            .I(N__48706));
    InMux I__11538 (
            .O(N__48709),
            .I(N__48703));
    LocalMux I__11537 (
            .O(N__48706),
            .I(N__48699));
    LocalMux I__11536 (
            .O(N__48703),
            .I(N__48696));
    InMux I__11535 (
            .O(N__48702),
            .I(N__48693));
    Span4Mux_h I__11534 (
            .O(N__48699),
            .I(N__48690));
    Odrv12 I__11533 (
            .O(N__48696),
            .I(\pid_front.error_p_regZ0Z_2 ));
    LocalMux I__11532 (
            .O(N__48693),
            .I(\pid_front.error_p_regZ0Z_2 ));
    Odrv4 I__11531 (
            .O(N__48690),
            .I(\pid_front.error_p_regZ0Z_2 ));
    InMux I__11530 (
            .O(N__48683),
            .I(N__48680));
    LocalMux I__11529 (
            .O(N__48680),
            .I(N__48677));
    Span4Mux_v I__11528 (
            .O(N__48677),
            .I(N__48674));
    Odrv4 I__11527 (
            .O(N__48674),
            .I(\pid_front.O_9 ));
    InMux I__11526 (
            .O(N__48671),
            .I(N__48668));
    LocalMux I__11525 (
            .O(N__48668),
            .I(N__48664));
    InMux I__11524 (
            .O(N__48667),
            .I(N__48661));
    Span4Mux_v I__11523 (
            .O(N__48664),
            .I(N__48657));
    LocalMux I__11522 (
            .O(N__48661),
            .I(N__48654));
    InMux I__11521 (
            .O(N__48660),
            .I(N__48651));
    Span4Mux_h I__11520 (
            .O(N__48657),
            .I(N__48648));
    Span12Mux_h I__11519 (
            .O(N__48654),
            .I(N__48645));
    LocalMux I__11518 (
            .O(N__48651),
            .I(\pid_front.error_p_regZ0Z_5 ));
    Odrv4 I__11517 (
            .O(N__48648),
            .I(\pid_front.error_p_regZ0Z_5 ));
    Odrv12 I__11516 (
            .O(N__48645),
            .I(\pid_front.error_p_regZ0Z_5 ));
    InMux I__11515 (
            .O(N__48638),
            .I(N__48635));
    LocalMux I__11514 (
            .O(N__48635),
            .I(N__48632));
    Span4Mux_v I__11513 (
            .O(N__48632),
            .I(N__48629));
    Odrv4 I__11512 (
            .O(N__48629),
            .I(\pid_front.O_8 ));
    InMux I__11511 (
            .O(N__48626),
            .I(N__48622));
    InMux I__11510 (
            .O(N__48625),
            .I(N__48619));
    LocalMux I__11509 (
            .O(N__48622),
            .I(N__48616));
    LocalMux I__11508 (
            .O(N__48619),
            .I(N__48613));
    Span4Mux_v I__11507 (
            .O(N__48616),
            .I(N__48609));
    Span4Mux_h I__11506 (
            .O(N__48613),
            .I(N__48606));
    InMux I__11505 (
            .O(N__48612),
            .I(N__48603));
    Span4Mux_h I__11504 (
            .O(N__48609),
            .I(N__48600));
    Span4Mux_h I__11503 (
            .O(N__48606),
            .I(N__48597));
    LocalMux I__11502 (
            .O(N__48603),
            .I(\pid_front.error_p_regZ0Z_4 ));
    Odrv4 I__11501 (
            .O(N__48600),
            .I(\pid_front.error_p_regZ0Z_4 ));
    Odrv4 I__11500 (
            .O(N__48597),
            .I(\pid_front.error_p_regZ0Z_4 ));
    InMux I__11499 (
            .O(N__48590),
            .I(N__48587));
    LocalMux I__11498 (
            .O(N__48587),
            .I(N__48584));
    Span4Mux_h I__11497 (
            .O(N__48584),
            .I(N__48581));
    Odrv4 I__11496 (
            .O(N__48581),
            .I(\pid_front.un1_pid_prereg_cry_17_THRU_CO ));
    InMux I__11495 (
            .O(N__48578),
            .I(\pid_front.un1_pid_prereg_cry_17 ));
    InMux I__11494 (
            .O(N__48575),
            .I(N__48572));
    LocalMux I__11493 (
            .O(N__48572),
            .I(N__48569));
    Span4Mux_v I__11492 (
            .O(N__48569),
            .I(N__48566));
    Odrv4 I__11491 (
            .O(N__48566),
            .I(\pid_front.un1_pid_prereg_cry_18_THRU_CO ));
    InMux I__11490 (
            .O(N__48563),
            .I(\pid_front.un1_pid_prereg_cry_18 ));
    InMux I__11489 (
            .O(N__48560),
            .I(N__48557));
    LocalMux I__11488 (
            .O(N__48557),
            .I(N__48554));
    Span4Mux_v I__11487 (
            .O(N__48554),
            .I(N__48551));
    Odrv4 I__11486 (
            .O(N__48551),
            .I(\pid_front.un1_pid_prereg_cry_19_THRU_CO ));
    InMux I__11485 (
            .O(N__48548),
            .I(\pid_front.un1_pid_prereg_cry_19 ));
    InMux I__11484 (
            .O(N__48545),
            .I(\pid_front.un1_pid_prereg_cry_20 ));
    CascadeMux I__11483 (
            .O(N__48542),
            .I(N__48539));
    InMux I__11482 (
            .O(N__48539),
            .I(N__48530));
    InMux I__11481 (
            .O(N__48538),
            .I(N__48530));
    InMux I__11480 (
            .O(N__48537),
            .I(N__48527));
    CascadeMux I__11479 (
            .O(N__48536),
            .I(N__48524));
    CascadeMux I__11478 (
            .O(N__48535),
            .I(N__48521));
    LocalMux I__11477 (
            .O(N__48530),
            .I(N__48516));
    LocalMux I__11476 (
            .O(N__48527),
            .I(N__48516));
    InMux I__11475 (
            .O(N__48524),
            .I(N__48513));
    InMux I__11474 (
            .O(N__48521),
            .I(N__48510));
    Span4Mux_h I__11473 (
            .O(N__48516),
            .I(N__48507));
    LocalMux I__11472 (
            .O(N__48513),
            .I(N__48504));
    LocalMux I__11471 (
            .O(N__48510),
            .I(N__48501));
    Span4Mux_v I__11470 (
            .O(N__48507),
            .I(N__48498));
    Span4Mux_h I__11469 (
            .O(N__48504),
            .I(N__48493));
    Span4Mux_v I__11468 (
            .O(N__48501),
            .I(N__48493));
    Span4Mux_h I__11467 (
            .O(N__48498),
            .I(N__48490));
    Span4Mux_h I__11466 (
            .O(N__48493),
            .I(N__48487));
    Odrv4 I__11465 (
            .O(N__48490),
            .I(\pid_front.pid_preregZ0Z_21 ));
    Odrv4 I__11464 (
            .O(N__48487),
            .I(\pid_front.pid_preregZ0Z_21 ));
    CEMux I__11463 (
            .O(N__48482),
            .I(N__48478));
    CEMux I__11462 (
            .O(N__48481),
            .I(N__48475));
    LocalMux I__11461 (
            .O(N__48478),
            .I(N__48472));
    LocalMux I__11460 (
            .O(N__48475),
            .I(N__48469));
    Span4Mux_h I__11459 (
            .O(N__48472),
            .I(N__48466));
    Span4Mux_v I__11458 (
            .O(N__48469),
            .I(N__48463));
    Span4Mux_h I__11457 (
            .O(N__48466),
            .I(N__48458));
    Span4Mux_h I__11456 (
            .O(N__48463),
            .I(N__48458));
    Odrv4 I__11455 (
            .O(N__48458),
            .I(\pid_front.state_0_0 ));
    InMux I__11454 (
            .O(N__48455),
            .I(N__48452));
    LocalMux I__11453 (
            .O(N__48452),
            .I(N__48449));
    Span4Mux_h I__11452 (
            .O(N__48449),
            .I(N__48445));
    InMux I__11451 (
            .O(N__48448),
            .I(N__48442));
    Span4Mux_v I__11450 (
            .O(N__48445),
            .I(N__48437));
    LocalMux I__11449 (
            .O(N__48442),
            .I(N__48437));
    Span4Mux_h I__11448 (
            .O(N__48437),
            .I(N__48430));
    InMux I__11447 (
            .O(N__48436),
            .I(N__48427));
    InMux I__11446 (
            .O(N__48435),
            .I(N__48423));
    InMux I__11445 (
            .O(N__48434),
            .I(N__48420));
    InMux I__11444 (
            .O(N__48433),
            .I(N__48417));
    Span4Mux_h I__11443 (
            .O(N__48430),
            .I(N__48412));
    LocalMux I__11442 (
            .O(N__48427),
            .I(N__48412));
    InMux I__11441 (
            .O(N__48426),
            .I(N__48409));
    LocalMux I__11440 (
            .O(N__48423),
            .I(N__48403));
    LocalMux I__11439 (
            .O(N__48420),
            .I(N__48403));
    LocalMux I__11438 (
            .O(N__48417),
            .I(N__48400));
    Span4Mux_v I__11437 (
            .O(N__48412),
            .I(N__48397));
    LocalMux I__11436 (
            .O(N__48409),
            .I(N__48394));
    CascadeMux I__11435 (
            .O(N__48408),
            .I(N__48391));
    Span12Mux_s10_h I__11434 (
            .O(N__48403),
            .I(N__48386));
    Span12Mux_s11_v I__11433 (
            .O(N__48400),
            .I(N__48386));
    Span4Mux_v I__11432 (
            .O(N__48397),
            .I(N__48381));
    Span4Mux_v I__11431 (
            .O(N__48394),
            .I(N__48381));
    InMux I__11430 (
            .O(N__48391),
            .I(N__48378));
    Odrv12 I__11429 (
            .O(N__48386),
            .I(uart_drone_data_6));
    Odrv4 I__11428 (
            .O(N__48381),
            .I(uart_drone_data_6));
    LocalMux I__11427 (
            .O(N__48378),
            .I(uart_drone_data_6));
    CascadeMux I__11426 (
            .O(N__48371),
            .I(N__48367));
    InMux I__11425 (
            .O(N__48370),
            .I(N__48362));
    InMux I__11424 (
            .O(N__48367),
            .I(N__48362));
    LocalMux I__11423 (
            .O(N__48362),
            .I(drone_H_disp_front_14));
    CEMux I__11422 (
            .O(N__48359),
            .I(N__48356));
    LocalMux I__11421 (
            .O(N__48356),
            .I(N__48351));
    CEMux I__11420 (
            .O(N__48355),
            .I(N__48348));
    CEMux I__11419 (
            .O(N__48354),
            .I(N__48345));
    Span4Mux_v I__11418 (
            .O(N__48351),
            .I(N__48341));
    LocalMux I__11417 (
            .O(N__48348),
            .I(N__48336));
    LocalMux I__11416 (
            .O(N__48345),
            .I(N__48336));
    CEMux I__11415 (
            .O(N__48344),
            .I(N__48333));
    Span4Mux_h I__11414 (
            .O(N__48341),
            .I(N__48326));
    Span4Mux_v I__11413 (
            .O(N__48336),
            .I(N__48326));
    LocalMux I__11412 (
            .O(N__48333),
            .I(N__48326));
    Span4Mux_h I__11411 (
            .O(N__48326),
            .I(N__48323));
    Span4Mux_v I__11410 (
            .O(N__48323),
            .I(N__48320));
    Span4Mux_v I__11409 (
            .O(N__48320),
            .I(N__48317));
    Odrv4 I__11408 (
            .O(N__48317),
            .I(\dron_frame_decoder_1.N_723_0 ));
    IoInMux I__11407 (
            .O(N__48314),
            .I(N__48311));
    LocalMux I__11406 (
            .O(N__48311),
            .I(GB_BUFFER_reset_system_g_THRU_CO));
    InMux I__11405 (
            .O(N__48308),
            .I(N__48305));
    LocalMux I__11404 (
            .O(N__48305),
            .I(N__48302));
    Span12Mux_h I__11403 (
            .O(N__48302),
            .I(N__48299));
    Odrv12 I__11402 (
            .O(N__48299),
            .I(\pid_side.O_0_4 ));
    InMux I__11401 (
            .O(N__48296),
            .I(N__48293));
    LocalMux I__11400 (
            .O(N__48293),
            .I(N__48290));
    Span4Mux_v I__11399 (
            .O(N__48290),
            .I(N__48286));
    InMux I__11398 (
            .O(N__48289),
            .I(N__48283));
    Odrv4 I__11397 (
            .O(N__48286),
            .I(\pid_side.error_p_regZ0Z_0 ));
    LocalMux I__11396 (
            .O(N__48283),
            .I(\pid_side.error_p_regZ0Z_0 ));
    InMux I__11395 (
            .O(N__48278),
            .I(N__48275));
    LocalMux I__11394 (
            .O(N__48275),
            .I(N__48272));
    Span12Mux_h I__11393 (
            .O(N__48272),
            .I(N__48269));
    Odrv12 I__11392 (
            .O(N__48269),
            .I(\pid_side.O_0_5 ));
    InMux I__11391 (
            .O(N__48266),
            .I(N__48263));
    LocalMux I__11390 (
            .O(N__48263),
            .I(N__48260));
    Span4Mux_h I__11389 (
            .O(N__48260),
            .I(N__48257));
    Odrv4 I__11388 (
            .O(N__48257),
            .I(\pid_front.un1_pid_prereg_cry_9_THRU_CO ));
    InMux I__11387 (
            .O(N__48254),
            .I(\pid_front.un1_pid_prereg_cry_9 ));
    InMux I__11386 (
            .O(N__48251),
            .I(N__48248));
    LocalMux I__11385 (
            .O(N__48248),
            .I(N__48245));
    Span4Mux_h I__11384 (
            .O(N__48245),
            .I(N__48242));
    Odrv4 I__11383 (
            .O(N__48242),
            .I(\pid_front.un1_pid_prereg_cry_10_THRU_CO ));
    InMux I__11382 (
            .O(N__48239),
            .I(\pid_front.un1_pid_prereg_cry_10 ));
    InMux I__11381 (
            .O(N__48236),
            .I(N__48226));
    InMux I__11380 (
            .O(N__48235),
            .I(N__48223));
    InMux I__11379 (
            .O(N__48234),
            .I(N__48220));
    InMux I__11378 (
            .O(N__48233),
            .I(N__48217));
    CascadeMux I__11377 (
            .O(N__48232),
            .I(N__48214));
    CascadeMux I__11376 (
            .O(N__48231),
            .I(N__48211));
    InMux I__11375 (
            .O(N__48230),
            .I(N__48203));
    InMux I__11374 (
            .O(N__48229),
            .I(N__48200));
    LocalMux I__11373 (
            .O(N__48226),
            .I(N__48194));
    LocalMux I__11372 (
            .O(N__48223),
            .I(N__48194));
    LocalMux I__11371 (
            .O(N__48220),
            .I(N__48185));
    LocalMux I__11370 (
            .O(N__48217),
            .I(N__48185));
    InMux I__11369 (
            .O(N__48214),
            .I(N__48180));
    InMux I__11368 (
            .O(N__48211),
            .I(N__48180));
    CascadeMux I__11367 (
            .O(N__48210),
            .I(N__48177));
    CascadeMux I__11366 (
            .O(N__48209),
            .I(N__48170));
    CascadeMux I__11365 (
            .O(N__48208),
            .I(N__48166));
    CascadeMux I__11364 (
            .O(N__48207),
            .I(N__48162));
    InMux I__11363 (
            .O(N__48206),
            .I(N__48158));
    LocalMux I__11362 (
            .O(N__48203),
            .I(N__48155));
    LocalMux I__11361 (
            .O(N__48200),
            .I(N__48152));
    InMux I__11360 (
            .O(N__48199),
            .I(N__48149));
    Span4Mux_v I__11359 (
            .O(N__48194),
            .I(N__48146));
    InMux I__11358 (
            .O(N__48193),
            .I(N__48143));
    InMux I__11357 (
            .O(N__48192),
            .I(N__48140));
    CascadeMux I__11356 (
            .O(N__48191),
            .I(N__48137));
    CascadeMux I__11355 (
            .O(N__48190),
            .I(N__48133));
    Span4Mux_v I__11354 (
            .O(N__48185),
            .I(N__48125));
    LocalMux I__11353 (
            .O(N__48180),
            .I(N__48122));
    InMux I__11352 (
            .O(N__48177),
            .I(N__48119));
    CascadeMux I__11351 (
            .O(N__48176),
            .I(N__48116));
    CascadeMux I__11350 (
            .O(N__48175),
            .I(N__48113));
    CascadeMux I__11349 (
            .O(N__48174),
            .I(N__48110));
    CascadeMux I__11348 (
            .O(N__48173),
            .I(N__48107));
    InMux I__11347 (
            .O(N__48170),
            .I(N__48099));
    InMux I__11346 (
            .O(N__48169),
            .I(N__48099));
    InMux I__11345 (
            .O(N__48166),
            .I(N__48096));
    InMux I__11344 (
            .O(N__48165),
            .I(N__48091));
    InMux I__11343 (
            .O(N__48162),
            .I(N__48091));
    CascadeMux I__11342 (
            .O(N__48161),
            .I(N__48088));
    LocalMux I__11341 (
            .O(N__48158),
            .I(N__48081));
    Span4Mux_v I__11340 (
            .O(N__48155),
            .I(N__48074));
    Span4Mux_v I__11339 (
            .O(N__48152),
            .I(N__48074));
    LocalMux I__11338 (
            .O(N__48149),
            .I(N__48074));
    Span4Mux_v I__11337 (
            .O(N__48146),
            .I(N__48069));
    LocalMux I__11336 (
            .O(N__48143),
            .I(N__48069));
    LocalMux I__11335 (
            .O(N__48140),
            .I(N__48066));
    InMux I__11334 (
            .O(N__48137),
            .I(N__48059));
    InMux I__11333 (
            .O(N__48136),
            .I(N__48059));
    InMux I__11332 (
            .O(N__48133),
            .I(N__48059));
    CascadeMux I__11331 (
            .O(N__48132),
            .I(N__48056));
    CascadeMux I__11330 (
            .O(N__48131),
            .I(N__48053));
    CascadeMux I__11329 (
            .O(N__48130),
            .I(N__48050));
    CascadeMux I__11328 (
            .O(N__48129),
            .I(N__48047));
    CascadeMux I__11327 (
            .O(N__48128),
            .I(N__48044));
    Span4Mux_h I__11326 (
            .O(N__48125),
            .I(N__48037));
    Span4Mux_v I__11325 (
            .O(N__48122),
            .I(N__48032));
    LocalMux I__11324 (
            .O(N__48119),
            .I(N__48032));
    InMux I__11323 (
            .O(N__48116),
            .I(N__48023));
    InMux I__11322 (
            .O(N__48113),
            .I(N__48023));
    InMux I__11321 (
            .O(N__48110),
            .I(N__48023));
    InMux I__11320 (
            .O(N__48107),
            .I(N__48023));
    CascadeMux I__11319 (
            .O(N__48106),
            .I(N__48020));
    CascadeMux I__11318 (
            .O(N__48105),
            .I(N__48017));
    CascadeMux I__11317 (
            .O(N__48104),
            .I(N__48014));
    LocalMux I__11316 (
            .O(N__48099),
            .I(N__48011));
    LocalMux I__11315 (
            .O(N__48096),
            .I(N__48006));
    LocalMux I__11314 (
            .O(N__48091),
            .I(N__48006));
    InMux I__11313 (
            .O(N__48088),
            .I(N__48003));
    CascadeMux I__11312 (
            .O(N__48087),
            .I(N__48000));
    CascadeMux I__11311 (
            .O(N__48086),
            .I(N__47997));
    CascadeMux I__11310 (
            .O(N__48085),
            .I(N__47994));
    CascadeMux I__11309 (
            .O(N__48084),
            .I(N__47991));
    Span4Mux_v I__11308 (
            .O(N__48081),
            .I(N__47982));
    Span4Mux_v I__11307 (
            .O(N__48074),
            .I(N__47982));
    Span4Mux_v I__11306 (
            .O(N__48069),
            .I(N__47982));
    Span4Mux_v I__11305 (
            .O(N__48066),
            .I(N__47979));
    LocalMux I__11304 (
            .O(N__48059),
            .I(N__47976));
    InMux I__11303 (
            .O(N__48056),
            .I(N__47971));
    InMux I__11302 (
            .O(N__48053),
            .I(N__47971));
    InMux I__11301 (
            .O(N__48050),
            .I(N__47966));
    InMux I__11300 (
            .O(N__48047),
            .I(N__47966));
    InMux I__11299 (
            .O(N__48044),
            .I(N__47963));
    CascadeMux I__11298 (
            .O(N__48043),
            .I(N__47960));
    CascadeMux I__11297 (
            .O(N__48042),
            .I(N__47957));
    CascadeMux I__11296 (
            .O(N__48041),
            .I(N__47954));
    CascadeMux I__11295 (
            .O(N__48040),
            .I(N__47951));
    Span4Mux_h I__11294 (
            .O(N__48037),
            .I(N__47948));
    Span4Mux_v I__11293 (
            .O(N__48032),
            .I(N__47943));
    LocalMux I__11292 (
            .O(N__48023),
            .I(N__47943));
    InMux I__11291 (
            .O(N__48020),
            .I(N__47936));
    InMux I__11290 (
            .O(N__48017),
            .I(N__47936));
    InMux I__11289 (
            .O(N__48014),
            .I(N__47936));
    Span4Mux_v I__11288 (
            .O(N__48011),
            .I(N__47929));
    Span4Mux_v I__11287 (
            .O(N__48006),
            .I(N__47929));
    LocalMux I__11286 (
            .O(N__48003),
            .I(N__47929));
    InMux I__11285 (
            .O(N__48000),
            .I(N__47926));
    InMux I__11284 (
            .O(N__47997),
            .I(N__47923));
    InMux I__11283 (
            .O(N__47994),
            .I(N__47918));
    InMux I__11282 (
            .O(N__47991),
            .I(N__47918));
    InMux I__11281 (
            .O(N__47990),
            .I(N__47915));
    InMux I__11280 (
            .O(N__47989),
            .I(N__47912));
    Span4Mux_h I__11279 (
            .O(N__47982),
            .I(N__47907));
    Span4Mux_h I__11278 (
            .O(N__47979),
            .I(N__47907));
    Span4Mux_v I__11277 (
            .O(N__47976),
            .I(N__47900));
    LocalMux I__11276 (
            .O(N__47971),
            .I(N__47900));
    LocalMux I__11275 (
            .O(N__47966),
            .I(N__47900));
    LocalMux I__11274 (
            .O(N__47963),
            .I(N__47897));
    InMux I__11273 (
            .O(N__47960),
            .I(N__47894));
    InMux I__11272 (
            .O(N__47957),
            .I(N__47891));
    InMux I__11271 (
            .O(N__47954),
            .I(N__47886));
    InMux I__11270 (
            .O(N__47951),
            .I(N__47886));
    Span4Mux_v I__11269 (
            .O(N__47948),
            .I(N__47880));
    Span4Mux_h I__11268 (
            .O(N__47943),
            .I(N__47875));
    LocalMux I__11267 (
            .O(N__47936),
            .I(N__47875));
    Span4Mux_v I__11266 (
            .O(N__47929),
            .I(N__47872));
    LocalMux I__11265 (
            .O(N__47926),
            .I(N__47865));
    LocalMux I__11264 (
            .O(N__47923),
            .I(N__47865));
    LocalMux I__11263 (
            .O(N__47918),
            .I(N__47865));
    LocalMux I__11262 (
            .O(N__47915),
            .I(N__47860));
    LocalMux I__11261 (
            .O(N__47912),
            .I(N__47860));
    Span4Mux_h I__11260 (
            .O(N__47907),
            .I(N__47853));
    Span4Mux_v I__11259 (
            .O(N__47900),
            .I(N__47853));
    Span4Mux_v I__11258 (
            .O(N__47897),
            .I(N__47853));
    LocalMux I__11257 (
            .O(N__47894),
            .I(N__47846));
    LocalMux I__11256 (
            .O(N__47891),
            .I(N__47846));
    LocalMux I__11255 (
            .O(N__47886),
            .I(N__47846));
    InMux I__11254 (
            .O(N__47885),
            .I(N__47843));
    CascadeMux I__11253 (
            .O(N__47884),
            .I(N__47839));
    CascadeMux I__11252 (
            .O(N__47883),
            .I(N__47836));
    Span4Mux_v I__11251 (
            .O(N__47880),
            .I(N__47833));
    Span4Mux_v I__11250 (
            .O(N__47875),
            .I(N__47830));
    Span4Mux_h I__11249 (
            .O(N__47872),
            .I(N__47823));
    Span4Mux_v I__11248 (
            .O(N__47865),
            .I(N__47823));
    Span4Mux_h I__11247 (
            .O(N__47860),
            .I(N__47823));
    Span4Mux_h I__11246 (
            .O(N__47853),
            .I(N__47816));
    Span4Mux_v I__11245 (
            .O(N__47846),
            .I(N__47816));
    LocalMux I__11244 (
            .O(N__47843),
            .I(N__47816));
    InMux I__11243 (
            .O(N__47842),
            .I(N__47809));
    InMux I__11242 (
            .O(N__47839),
            .I(N__47809));
    InMux I__11241 (
            .O(N__47836),
            .I(N__47809));
    Odrv4 I__11240 (
            .O(N__47833),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11239 (
            .O(N__47830),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11238 (
            .O(N__47823),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11237 (
            .O(N__47816),
            .I(CONSTANT_ONE_NET));
    LocalMux I__11236 (
            .O(N__47809),
            .I(CONSTANT_ONE_NET));
    InMux I__11235 (
            .O(N__47798),
            .I(N__47795));
    LocalMux I__11234 (
            .O(N__47795),
            .I(N__47792));
    Span4Mux_h I__11233 (
            .O(N__47792),
            .I(N__47789));
    Odrv4 I__11232 (
            .O(N__47789),
            .I(\pid_front.un1_pid_prereg_cry_11_THRU_CO ));
    InMux I__11231 (
            .O(N__47786),
            .I(\pid_front.un1_pid_prereg_cry_11 ));
    InMux I__11230 (
            .O(N__47783),
            .I(N__47780));
    LocalMux I__11229 (
            .O(N__47780),
            .I(N__47777));
    Span4Mux_h I__11228 (
            .O(N__47777),
            .I(N__47774));
    Odrv4 I__11227 (
            .O(N__47774),
            .I(\pid_front.un1_pid_prereg_cry_12_THRU_CO ));
    InMux I__11226 (
            .O(N__47771),
            .I(\pid_front.un1_pid_prereg_cry_12 ));
    InMux I__11225 (
            .O(N__47768),
            .I(N__47765));
    LocalMux I__11224 (
            .O(N__47765),
            .I(N__47762));
    Span4Mux_v I__11223 (
            .O(N__47762),
            .I(N__47759));
    Odrv4 I__11222 (
            .O(N__47759),
            .I(\pid_front.un1_pid_prereg_cry_13_THRU_CO ));
    InMux I__11221 (
            .O(N__47756),
            .I(\pid_front.un1_pid_prereg_cry_13 ));
    InMux I__11220 (
            .O(N__47753),
            .I(N__47750));
    LocalMux I__11219 (
            .O(N__47750),
            .I(N__47747));
    Odrv4 I__11218 (
            .O(N__47747),
            .I(\pid_front.un1_pid_prereg_cry_14_THRU_CO ));
    InMux I__11217 (
            .O(N__47744),
            .I(\pid_front.un1_pid_prereg_cry_14 ));
    InMux I__11216 (
            .O(N__47741),
            .I(N__47738));
    LocalMux I__11215 (
            .O(N__47738),
            .I(N__47735));
    Odrv4 I__11214 (
            .O(N__47735),
            .I(\pid_front.un1_pid_prereg_cry_15_THRU_CO ));
    InMux I__11213 (
            .O(N__47732),
            .I(\pid_front.un1_pid_prereg_cry_15 ));
    InMux I__11212 (
            .O(N__47729),
            .I(N__47726));
    LocalMux I__11211 (
            .O(N__47726),
            .I(N__47723));
    Span4Mux_h I__11210 (
            .O(N__47723),
            .I(N__47720));
    Odrv4 I__11209 (
            .O(N__47720),
            .I(\pid_front.un1_pid_prereg_cry_16_THRU_CO ));
    InMux I__11208 (
            .O(N__47717),
            .I(bfn_18_24_0_));
    SRMux I__11207 (
            .O(N__47714),
            .I(N__47705));
    SRMux I__11206 (
            .O(N__47713),
            .I(N__47705));
    SRMux I__11205 (
            .O(N__47712),
            .I(N__47705));
    GlobalMux I__11204 (
            .O(N__47705),
            .I(N__47702));
    gio2CtrlBuf I__11203 (
            .O(N__47702),
            .I(\ppm_encoder_1.N_661_g ));
    CascadeMux I__11202 (
            .O(N__47699),
            .I(N__47696));
    InMux I__11201 (
            .O(N__47696),
            .I(N__47693));
    LocalMux I__11200 (
            .O(N__47693),
            .I(N__47690));
    Span4Mux_h I__11199 (
            .O(N__47690),
            .I(N__47687));
    Odrv4 I__11198 (
            .O(N__47687),
            .I(\pid_front.un1_pid_prereg_cry_1_THRU_CO ));
    InMux I__11197 (
            .O(N__47684),
            .I(\pid_front.un1_pid_prereg_cry_1 ));
    CascadeMux I__11196 (
            .O(N__47681),
            .I(N__47678));
    InMux I__11195 (
            .O(N__47678),
            .I(N__47675));
    LocalMux I__11194 (
            .O(N__47675),
            .I(N__47672));
    Span4Mux_h I__11193 (
            .O(N__47672),
            .I(N__47669));
    Odrv4 I__11192 (
            .O(N__47669),
            .I(\pid_front.un1_pid_prereg_cry_2_THRU_CO ));
    InMux I__11191 (
            .O(N__47666),
            .I(\pid_front.un1_pid_prereg_cry_2 ));
    CascadeMux I__11190 (
            .O(N__47663),
            .I(N__47660));
    InMux I__11189 (
            .O(N__47660),
            .I(N__47657));
    LocalMux I__11188 (
            .O(N__47657),
            .I(N__47654));
    Span4Mux_v I__11187 (
            .O(N__47654),
            .I(N__47651));
    Odrv4 I__11186 (
            .O(N__47651),
            .I(\pid_front.un1_pid_prereg_cry_3_THRU_CO ));
    InMux I__11185 (
            .O(N__47648),
            .I(\pid_front.un1_pid_prereg_cry_3 ));
    CascadeMux I__11184 (
            .O(N__47645),
            .I(N__47642));
    InMux I__11183 (
            .O(N__47642),
            .I(N__47639));
    LocalMux I__11182 (
            .O(N__47639),
            .I(N__47636));
    Span4Mux_h I__11181 (
            .O(N__47636),
            .I(N__47633));
    Odrv4 I__11180 (
            .O(N__47633),
            .I(\pid_front.un1_pid_prereg_cry_4_THRU_CO ));
    InMux I__11179 (
            .O(N__47630),
            .I(\pid_front.un1_pid_prereg_cry_4 ));
    InMux I__11178 (
            .O(N__47627),
            .I(N__47624));
    LocalMux I__11177 (
            .O(N__47624),
            .I(N__47621));
    Span4Mux_h I__11176 (
            .O(N__47621),
            .I(N__47618));
    Odrv4 I__11175 (
            .O(N__47618),
            .I(\pid_front.un1_pid_prereg_cry_5_THRU_CO ));
    InMux I__11174 (
            .O(N__47615),
            .I(\pid_front.un1_pid_prereg_cry_5 ));
    InMux I__11173 (
            .O(N__47612),
            .I(N__47609));
    LocalMux I__11172 (
            .O(N__47609),
            .I(N__47606));
    Odrv12 I__11171 (
            .O(N__47606),
            .I(\pid_front.un1_pid_prereg_cry_6_THRU_CO ));
    InMux I__11170 (
            .O(N__47603),
            .I(\pid_front.un1_pid_prereg_cry_6 ));
    InMux I__11169 (
            .O(N__47600),
            .I(N__47597));
    LocalMux I__11168 (
            .O(N__47597),
            .I(\pid_front.un1_pid_prereg_cry_7_THRU_CO ));
    InMux I__11167 (
            .O(N__47594),
            .I(\pid_front.un1_pid_prereg_cry_7 ));
    InMux I__11166 (
            .O(N__47591),
            .I(N__47588));
    LocalMux I__11165 (
            .O(N__47588),
            .I(N__47585));
    Span4Mux_h I__11164 (
            .O(N__47585),
            .I(N__47582));
    Odrv4 I__11163 (
            .O(N__47582),
            .I(\pid_front.un1_pid_prereg_cry_8_THRU_CO ));
    InMux I__11162 (
            .O(N__47579),
            .I(bfn_18_23_0_));
    InMux I__11161 (
            .O(N__47576),
            .I(N__47571));
    InMux I__11160 (
            .O(N__47575),
            .I(N__47568));
    InMux I__11159 (
            .O(N__47574),
            .I(N__47565));
    LocalMux I__11158 (
            .O(N__47571),
            .I(N__47562));
    LocalMux I__11157 (
            .O(N__47568),
            .I(N__47559));
    LocalMux I__11156 (
            .O(N__47565),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__11155 (
            .O(N__47562),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    Odrv4 I__11154 (
            .O(N__47559),
            .I(\ppm_encoder_1.counterZ0Z_11 ));
    InMux I__11153 (
            .O(N__47552),
            .I(\ppm_encoder_1.un1_counter_13_cry_10 ));
    InMux I__11152 (
            .O(N__47549),
            .I(N__47544));
    InMux I__11151 (
            .O(N__47548),
            .I(N__47541));
    InMux I__11150 (
            .O(N__47547),
            .I(N__47538));
    LocalMux I__11149 (
            .O(N__47544),
            .I(N__47535));
    LocalMux I__11148 (
            .O(N__47541),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    LocalMux I__11147 (
            .O(N__47538),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    Odrv4 I__11146 (
            .O(N__47535),
            .I(\ppm_encoder_1.counterZ0Z_12 ));
    InMux I__11145 (
            .O(N__47528),
            .I(\ppm_encoder_1.un1_counter_13_cry_11 ));
    InMux I__11144 (
            .O(N__47525),
            .I(N__47520));
    InMux I__11143 (
            .O(N__47524),
            .I(N__47517));
    InMux I__11142 (
            .O(N__47523),
            .I(N__47514));
    LocalMux I__11141 (
            .O(N__47520),
            .I(N__47511));
    LocalMux I__11140 (
            .O(N__47517),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    LocalMux I__11139 (
            .O(N__47514),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    Odrv4 I__11138 (
            .O(N__47511),
            .I(\ppm_encoder_1.counterZ0Z_13 ));
    InMux I__11137 (
            .O(N__47504),
            .I(\ppm_encoder_1.un1_counter_13_cry_12 ));
    InMux I__11136 (
            .O(N__47501),
            .I(N__47498));
    LocalMux I__11135 (
            .O(N__47498),
            .I(N__47493));
    InMux I__11134 (
            .O(N__47497),
            .I(N__47490));
    InMux I__11133 (
            .O(N__47496),
            .I(N__47487));
    Span4Mux_v I__11132 (
            .O(N__47493),
            .I(N__47484));
    LocalMux I__11131 (
            .O(N__47490),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    LocalMux I__11130 (
            .O(N__47487),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    Odrv4 I__11129 (
            .O(N__47484),
            .I(\ppm_encoder_1.counterZ0Z_14 ));
    InMux I__11128 (
            .O(N__47477),
            .I(\ppm_encoder_1.un1_counter_13_cry_13 ));
    CascadeMux I__11127 (
            .O(N__47474),
            .I(N__47471));
    InMux I__11126 (
            .O(N__47471),
            .I(N__47468));
    LocalMux I__11125 (
            .O(N__47468),
            .I(N__47463));
    InMux I__11124 (
            .O(N__47467),
            .I(N__47460));
    InMux I__11123 (
            .O(N__47466),
            .I(N__47457));
    Span4Mux_v I__11122 (
            .O(N__47463),
            .I(N__47454));
    LocalMux I__11121 (
            .O(N__47460),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    LocalMux I__11120 (
            .O(N__47457),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    Odrv4 I__11119 (
            .O(N__47454),
            .I(\ppm_encoder_1.counterZ0Z_15 ));
    InMux I__11118 (
            .O(N__47447),
            .I(\ppm_encoder_1.un1_counter_13_cry_14 ));
    InMux I__11117 (
            .O(N__47444),
            .I(N__47439));
    InMux I__11116 (
            .O(N__47443),
            .I(N__47436));
    InMux I__11115 (
            .O(N__47442),
            .I(N__47433));
    LocalMux I__11114 (
            .O(N__47439),
            .I(N__47430));
    LocalMux I__11113 (
            .O(N__47436),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    LocalMux I__11112 (
            .O(N__47433),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    Odrv12 I__11111 (
            .O(N__47430),
            .I(\ppm_encoder_1.counterZ0Z_16 ));
    InMux I__11110 (
            .O(N__47423),
            .I(bfn_18_21_0_));
    InMux I__11109 (
            .O(N__47420),
            .I(N__47415));
    InMux I__11108 (
            .O(N__47419),
            .I(N__47412));
    InMux I__11107 (
            .O(N__47418),
            .I(N__47409));
    LocalMux I__11106 (
            .O(N__47415),
            .I(N__47406));
    LocalMux I__11105 (
            .O(N__47412),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    LocalMux I__11104 (
            .O(N__47409),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    Odrv12 I__11103 (
            .O(N__47406),
            .I(\ppm_encoder_1.counterZ0Z_17 ));
    InMux I__11102 (
            .O(N__47399),
            .I(\ppm_encoder_1.un1_counter_13_cry_16 ));
    InMux I__11101 (
            .O(N__47396),
            .I(\ppm_encoder_1.un1_counter_13_cry_17 ));
    CascadeMux I__11100 (
            .O(N__47393),
            .I(N__47388));
    InMux I__11099 (
            .O(N__47392),
            .I(N__47385));
    InMux I__11098 (
            .O(N__47391),
            .I(N__47382));
    InMux I__11097 (
            .O(N__47388),
            .I(N__47379));
    LocalMux I__11096 (
            .O(N__47385),
            .I(N__47376));
    LocalMux I__11095 (
            .O(N__47382),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    LocalMux I__11094 (
            .O(N__47379),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    Odrv12 I__11093 (
            .O(N__47376),
            .I(\ppm_encoder_1.counterZ0Z_18 ));
    InMux I__11092 (
            .O(N__47369),
            .I(\ppm_encoder_1.un1_counter_13_cry_1 ));
    InMux I__11091 (
            .O(N__47366),
            .I(N__47360));
    InMux I__11090 (
            .O(N__47365),
            .I(N__47355));
    InMux I__11089 (
            .O(N__47364),
            .I(N__47355));
    InMux I__11088 (
            .O(N__47363),
            .I(N__47352));
    LocalMux I__11087 (
            .O(N__47360),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__11086 (
            .O(N__47355),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    LocalMux I__11085 (
            .O(N__47352),
            .I(\ppm_encoder_1.counterZ0Z_3 ));
    InMux I__11084 (
            .O(N__47345),
            .I(\ppm_encoder_1.un1_counter_13_cry_2 ));
    InMux I__11083 (
            .O(N__47342),
            .I(N__47337));
    InMux I__11082 (
            .O(N__47341),
            .I(N__47334));
    InMux I__11081 (
            .O(N__47340),
            .I(N__47331));
    LocalMux I__11080 (
            .O(N__47337),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__11079 (
            .O(N__47334),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    LocalMux I__11078 (
            .O(N__47331),
            .I(\ppm_encoder_1.counterZ0Z_4 ));
    InMux I__11077 (
            .O(N__47324),
            .I(\ppm_encoder_1.un1_counter_13_cry_3 ));
    InMux I__11076 (
            .O(N__47321),
            .I(N__47316));
    InMux I__11075 (
            .O(N__47320),
            .I(N__47313));
    InMux I__11074 (
            .O(N__47319),
            .I(N__47310));
    LocalMux I__11073 (
            .O(N__47316),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__11072 (
            .O(N__47313),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    LocalMux I__11071 (
            .O(N__47310),
            .I(\ppm_encoder_1.counterZ0Z_5 ));
    InMux I__11070 (
            .O(N__47303),
            .I(\ppm_encoder_1.un1_counter_13_cry_4 ));
    InMux I__11069 (
            .O(N__47300),
            .I(N__47295));
    InMux I__11068 (
            .O(N__47299),
            .I(N__47292));
    InMux I__11067 (
            .O(N__47298),
            .I(N__47289));
    LocalMux I__11066 (
            .O(N__47295),
            .I(N__47286));
    LocalMux I__11065 (
            .O(N__47292),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    LocalMux I__11064 (
            .O(N__47289),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    Odrv12 I__11063 (
            .O(N__47286),
            .I(\ppm_encoder_1.counterZ0Z_6 ));
    InMux I__11062 (
            .O(N__47279),
            .I(\ppm_encoder_1.un1_counter_13_cry_5 ));
    InMux I__11061 (
            .O(N__47276),
            .I(N__47272));
    CascadeMux I__11060 (
            .O(N__47275),
            .I(N__47268));
    LocalMux I__11059 (
            .O(N__47272),
            .I(N__47265));
    InMux I__11058 (
            .O(N__47271),
            .I(N__47262));
    InMux I__11057 (
            .O(N__47268),
            .I(N__47259));
    Span4Mux_v I__11056 (
            .O(N__47265),
            .I(N__47256));
    LocalMux I__11055 (
            .O(N__47262),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    LocalMux I__11054 (
            .O(N__47259),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    Odrv4 I__11053 (
            .O(N__47256),
            .I(\ppm_encoder_1.counterZ0Z_7 ));
    InMux I__11052 (
            .O(N__47249),
            .I(\ppm_encoder_1.un1_counter_13_cry_6 ));
    InMux I__11051 (
            .O(N__47246),
            .I(N__47241));
    InMux I__11050 (
            .O(N__47245),
            .I(N__47238));
    InMux I__11049 (
            .O(N__47244),
            .I(N__47235));
    LocalMux I__11048 (
            .O(N__47241),
            .I(N__47232));
    LocalMux I__11047 (
            .O(N__47238),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    LocalMux I__11046 (
            .O(N__47235),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    Odrv4 I__11045 (
            .O(N__47232),
            .I(\ppm_encoder_1.counterZ0Z_8 ));
    InMux I__11044 (
            .O(N__47225),
            .I(bfn_18_20_0_));
    InMux I__11043 (
            .O(N__47222),
            .I(N__47215));
    InMux I__11042 (
            .O(N__47221),
            .I(N__47215));
    InMux I__11041 (
            .O(N__47220),
            .I(N__47212));
    LocalMux I__11040 (
            .O(N__47215),
            .I(N__47209));
    LocalMux I__11039 (
            .O(N__47212),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    Odrv4 I__11038 (
            .O(N__47209),
            .I(\ppm_encoder_1.counterZ0Z_9 ));
    InMux I__11037 (
            .O(N__47204),
            .I(\ppm_encoder_1.un1_counter_13_cry_8 ));
    CascadeMux I__11036 (
            .O(N__47201),
            .I(N__47198));
    InMux I__11035 (
            .O(N__47198),
            .I(N__47191));
    InMux I__11034 (
            .O(N__47197),
            .I(N__47191));
    InMux I__11033 (
            .O(N__47196),
            .I(N__47188));
    LocalMux I__11032 (
            .O(N__47191),
            .I(N__47185));
    LocalMux I__11031 (
            .O(N__47188),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    Odrv4 I__11030 (
            .O(N__47185),
            .I(\ppm_encoder_1.counterZ0Z_10 ));
    InMux I__11029 (
            .O(N__47180),
            .I(\ppm_encoder_1.un1_counter_13_cry_9 ));
    InMux I__11028 (
            .O(N__47177),
            .I(\ppm_encoder_1.counter24_0_N_2 ));
    InMux I__11027 (
            .O(N__47174),
            .I(N__47167));
    InMux I__11026 (
            .O(N__47173),
            .I(N__47167));
    CascadeMux I__11025 (
            .O(N__47172),
            .I(N__47164));
    LocalMux I__11024 (
            .O(N__47167),
            .I(N__47160));
    InMux I__11023 (
            .O(N__47164),
            .I(N__47155));
    InMux I__11022 (
            .O(N__47163),
            .I(N__47155));
    Odrv4 I__11021 (
            .O(N__47160),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    LocalMux I__11020 (
            .O(N__47155),
            .I(\ppm_encoder_1.counter24_0_N_2_THRU_CO ));
    InMux I__11019 (
            .O(N__47150),
            .I(N__47147));
    LocalMux I__11018 (
            .O(N__47147),
            .I(N__47144));
    Odrv12 I__11017 (
            .O(N__47144),
            .I(\ppm_encoder_1.pulses2countZ0Z_4 ));
    CascadeMux I__11016 (
            .O(N__47141),
            .I(N__47138));
    InMux I__11015 (
            .O(N__47138),
            .I(N__47135));
    LocalMux I__11014 (
            .O(N__47135),
            .I(N__47132));
    Span4Mux_v I__11013 (
            .O(N__47132),
            .I(N__47129));
    Odrv4 I__11012 (
            .O(N__47129),
            .I(\ppm_encoder_1.pulses2countZ0Z_5 ));
    InMux I__11011 (
            .O(N__47126),
            .I(N__47123));
    LocalMux I__11010 (
            .O(N__47123),
            .I(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ));
    InMux I__11009 (
            .O(N__47120),
            .I(N__47117));
    LocalMux I__11008 (
            .O(N__47117),
            .I(N__47114));
    Span4Mux_v I__11007 (
            .O(N__47114),
            .I(N__47111));
    Odrv4 I__11006 (
            .O(N__47111),
            .I(\ppm_encoder_1.pulses2countZ0Z_10 ));
    CascadeMux I__11005 (
            .O(N__47108),
            .I(N__47105));
    InMux I__11004 (
            .O(N__47105),
            .I(N__47102));
    LocalMux I__11003 (
            .O(N__47102),
            .I(N__47099));
    Span4Mux_v I__11002 (
            .O(N__47099),
            .I(N__47096));
    Odrv4 I__11001 (
            .O(N__47096),
            .I(\ppm_encoder_1.pulses2countZ0Z_11 ));
    InMux I__11000 (
            .O(N__47093),
            .I(N__47090));
    LocalMux I__10999 (
            .O(N__47090),
            .I(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ));
    InMux I__10998 (
            .O(N__47087),
            .I(N__47081));
    InMux I__10997 (
            .O(N__47086),
            .I(N__47081));
    LocalMux I__10996 (
            .O(N__47081),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ));
    InMux I__10995 (
            .O(N__47078),
            .I(N__47075));
    LocalMux I__10994 (
            .O(N__47075),
            .I(N__47072));
    Odrv12 I__10993 (
            .O(N__47072),
            .I(\ppm_encoder_1.pulses2countZ0Z_8 ));
    CascadeMux I__10992 (
            .O(N__47069),
            .I(N__47066));
    InMux I__10991 (
            .O(N__47066),
            .I(N__47063));
    LocalMux I__10990 (
            .O(N__47063),
            .I(N__47060));
    Span4Mux_h I__10989 (
            .O(N__47060),
            .I(N__47057));
    Odrv4 I__10988 (
            .O(N__47057),
            .I(\ppm_encoder_1.pulses2countZ0Z_9 ));
    InMux I__10987 (
            .O(N__47054),
            .I(N__47051));
    LocalMux I__10986 (
            .O(N__47051),
            .I(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ));
    InMux I__10985 (
            .O(N__47048),
            .I(N__47045));
    LocalMux I__10984 (
            .O(N__47045),
            .I(N__47042));
    Span4Mux_v I__10983 (
            .O(N__47042),
            .I(N__47039));
    Odrv4 I__10982 (
            .O(N__47039),
            .I(\ppm_encoder_1.pulses2countZ0Z_12 ));
    CascadeMux I__10981 (
            .O(N__47036),
            .I(N__47033));
    InMux I__10980 (
            .O(N__47033),
            .I(N__47030));
    LocalMux I__10979 (
            .O(N__47030),
            .I(N__47027));
    Span4Mux_v I__10978 (
            .O(N__47027),
            .I(N__47024));
    Odrv4 I__10977 (
            .O(N__47024),
            .I(\ppm_encoder_1.pulses2countZ0Z_13 ));
    InMux I__10976 (
            .O(N__47021),
            .I(N__47018));
    LocalMux I__10975 (
            .O(N__47018),
            .I(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ));
    InMux I__10974 (
            .O(N__47015),
            .I(N__47011));
    CascadeMux I__10973 (
            .O(N__47014),
            .I(N__47008));
    LocalMux I__10972 (
            .O(N__47011),
            .I(N__47005));
    InMux I__10971 (
            .O(N__47008),
            .I(N__47002));
    Odrv4 I__10970 (
            .O(N__47005),
            .I(\ppm_encoder_1.N_1818_i ));
    LocalMux I__10969 (
            .O(N__47002),
            .I(\ppm_encoder_1.N_1818_i ));
    InMux I__10968 (
            .O(N__46997),
            .I(N__46992));
    InMux I__10967 (
            .O(N__46996),
            .I(N__46989));
    InMux I__10966 (
            .O(N__46995),
            .I(N__46986));
    LocalMux I__10965 (
            .O(N__46992),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__10964 (
            .O(N__46989),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    LocalMux I__10963 (
            .O(N__46986),
            .I(\ppm_encoder_1.counterZ0Z_0 ));
    InMux I__10962 (
            .O(N__46979),
            .I(N__46973));
    InMux I__10961 (
            .O(N__46978),
            .I(N__46966));
    InMux I__10960 (
            .O(N__46977),
            .I(N__46966));
    InMux I__10959 (
            .O(N__46976),
            .I(N__46966));
    LocalMux I__10958 (
            .O(N__46973),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    LocalMux I__10957 (
            .O(N__46966),
            .I(\ppm_encoder_1.counterZ0Z_1 ));
    InMux I__10956 (
            .O(N__46961),
            .I(\ppm_encoder_1.un1_counter_13_cry_0 ));
    CascadeMux I__10955 (
            .O(N__46958),
            .I(N__46955));
    InMux I__10954 (
            .O(N__46955),
            .I(N__46950));
    CascadeMux I__10953 (
            .O(N__46954),
            .I(N__46947));
    InMux I__10952 (
            .O(N__46953),
            .I(N__46943));
    LocalMux I__10951 (
            .O(N__46950),
            .I(N__46940));
    InMux I__10950 (
            .O(N__46947),
            .I(N__46935));
    InMux I__10949 (
            .O(N__46946),
            .I(N__46935));
    LocalMux I__10948 (
            .O(N__46943),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    Odrv4 I__10947 (
            .O(N__46940),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    LocalMux I__10946 (
            .O(N__46935),
            .I(\ppm_encoder_1.counterZ0Z_2 ));
    InMux I__10945 (
            .O(N__46928),
            .I(N__46925));
    LocalMux I__10944 (
            .O(N__46925),
            .I(N__46922));
    Odrv12 I__10943 (
            .O(N__46922),
            .I(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ));
    InMux I__10942 (
            .O(N__46919),
            .I(N__46916));
    LocalMux I__10941 (
            .O(N__46916),
            .I(N__46913));
    Odrv4 I__10940 (
            .O(N__46913),
            .I(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ));
    InMux I__10939 (
            .O(N__46910),
            .I(N__46907));
    LocalMux I__10938 (
            .O(N__46907),
            .I(N__46904));
    Span4Mux_v I__10937 (
            .O(N__46904),
            .I(N__46901));
    Odrv4 I__10936 (
            .O(N__46901),
            .I(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ));
    InMux I__10935 (
            .O(N__46898),
            .I(N__46895));
    LocalMux I__10934 (
            .O(N__46895),
            .I(N__46892));
    Odrv12 I__10933 (
            .O(N__46892),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ));
    InMux I__10932 (
            .O(N__46889),
            .I(N__46886));
    LocalMux I__10931 (
            .O(N__46886),
            .I(N__46883));
    Odrv12 I__10930 (
            .O(N__46883),
            .I(\ppm_encoder_1.un2_throttle_iv_1_4 ));
    InMux I__10929 (
            .O(N__46880),
            .I(N__46877));
    LocalMux I__10928 (
            .O(N__46877),
            .I(N__46874));
    Span4Mux_v I__10927 (
            .O(N__46874),
            .I(N__46871));
    Odrv4 I__10926 (
            .O(N__46871),
            .I(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ));
    InMux I__10925 (
            .O(N__46868),
            .I(N__46864));
    InMux I__10924 (
            .O(N__46867),
            .I(N__46861));
    LocalMux I__10923 (
            .O(N__46864),
            .I(N__46858));
    LocalMux I__10922 (
            .O(N__46861),
            .I(N__46853));
    Span4Mux_v I__10921 (
            .O(N__46858),
            .I(N__46853));
    Odrv4 I__10920 (
            .O(N__46853),
            .I(side_order_4));
    CascadeMux I__10919 (
            .O(N__46850),
            .I(N__46847));
    InMux I__10918 (
            .O(N__46847),
            .I(N__46844));
    LocalMux I__10917 (
            .O(N__46844),
            .I(N__46841));
    Span4Mux_h I__10916 (
            .O(N__46841),
            .I(N__46838));
    Odrv4 I__10915 (
            .O(N__46838),
            .I(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ));
    InMux I__10914 (
            .O(N__46835),
            .I(N__46832));
    LocalMux I__10913 (
            .O(N__46832),
            .I(N__46828));
    InMux I__10912 (
            .O(N__46831),
            .I(N__46825));
    Span4Mux_v I__10911 (
            .O(N__46828),
            .I(N__46820));
    LocalMux I__10910 (
            .O(N__46825),
            .I(N__46820));
    Span4Mux_h I__10909 (
            .O(N__46820),
            .I(N__46817));
    Odrv4 I__10908 (
            .O(N__46817),
            .I(front_order_4));
    InMux I__10907 (
            .O(N__46814),
            .I(N__46808));
    CascadeMux I__10906 (
            .O(N__46813),
            .I(N__46802));
    InMux I__10905 (
            .O(N__46812),
            .I(N__46799));
    InMux I__10904 (
            .O(N__46811),
            .I(N__46796));
    LocalMux I__10903 (
            .O(N__46808),
            .I(N__46792));
    InMux I__10902 (
            .O(N__46807),
            .I(N__46789));
    InMux I__10901 (
            .O(N__46806),
            .I(N__46783));
    InMux I__10900 (
            .O(N__46805),
            .I(N__46779));
    InMux I__10899 (
            .O(N__46802),
            .I(N__46776));
    LocalMux I__10898 (
            .O(N__46799),
            .I(N__46771));
    LocalMux I__10897 (
            .O(N__46796),
            .I(N__46771));
    InMux I__10896 (
            .O(N__46795),
            .I(N__46768));
    Span4Mux_v I__10895 (
            .O(N__46792),
            .I(N__46760));
    LocalMux I__10894 (
            .O(N__46789),
            .I(N__46760));
    InMux I__10893 (
            .O(N__46788),
            .I(N__46755));
    InMux I__10892 (
            .O(N__46787),
            .I(N__46755));
    InMux I__10891 (
            .O(N__46786),
            .I(N__46749));
    LocalMux I__10890 (
            .O(N__46783),
            .I(N__46746));
    InMux I__10889 (
            .O(N__46782),
            .I(N__46742));
    LocalMux I__10888 (
            .O(N__46779),
            .I(N__46733));
    LocalMux I__10887 (
            .O(N__46776),
            .I(N__46733));
    Span4Mux_v I__10886 (
            .O(N__46771),
            .I(N__46733));
    LocalMux I__10885 (
            .O(N__46768),
            .I(N__46733));
    InMux I__10884 (
            .O(N__46767),
            .I(N__46730));
    InMux I__10883 (
            .O(N__46766),
            .I(N__46725));
    InMux I__10882 (
            .O(N__46765),
            .I(N__46725));
    Span4Mux_h I__10881 (
            .O(N__46760),
            .I(N__46720));
    LocalMux I__10880 (
            .O(N__46755),
            .I(N__46720));
    InMux I__10879 (
            .O(N__46754),
            .I(N__46713));
    InMux I__10878 (
            .O(N__46753),
            .I(N__46713));
    InMux I__10877 (
            .O(N__46752),
            .I(N__46713));
    LocalMux I__10876 (
            .O(N__46749),
            .I(N__46708));
    Span4Mux_v I__10875 (
            .O(N__46746),
            .I(N__46708));
    InMux I__10874 (
            .O(N__46745),
            .I(N__46705));
    LocalMux I__10873 (
            .O(N__46742),
            .I(N__46700));
    Span4Mux_h I__10872 (
            .O(N__46733),
            .I(N__46700));
    LocalMux I__10871 (
            .O(N__46730),
            .I(N__46693));
    LocalMux I__10870 (
            .O(N__46725),
            .I(N__46693));
    Sp12to4 I__10869 (
            .O(N__46720),
            .I(N__46693));
    LocalMux I__10868 (
            .O(N__46713),
            .I(N__46690));
    Odrv4 I__10867 (
            .O(N__46708),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    LocalMux I__10866 (
            .O(N__46705),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv4 I__10865 (
            .O(N__46700),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv12 I__10864 (
            .O(N__46693),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    Odrv12 I__10863 (
            .O(N__46690),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ));
    InMux I__10862 (
            .O(N__46679),
            .I(N__46670));
    InMux I__10861 (
            .O(N__46678),
            .I(N__46670));
    InMux I__10860 (
            .O(N__46677),
            .I(N__46670));
    LocalMux I__10859 (
            .O(N__46670),
            .I(\ppm_encoder_1.elevatorZ0Z_4 ));
    InMux I__10858 (
            .O(N__46667),
            .I(N__46659));
    CascadeMux I__10857 (
            .O(N__46666),
            .I(N__46656));
    InMux I__10856 (
            .O(N__46665),
            .I(N__46652));
    InMux I__10855 (
            .O(N__46664),
            .I(N__46649));
    InMux I__10854 (
            .O(N__46663),
            .I(N__46646));
    CascadeMux I__10853 (
            .O(N__46662),
            .I(N__46639));
    LocalMux I__10852 (
            .O(N__46659),
            .I(N__46636));
    InMux I__10851 (
            .O(N__46656),
            .I(N__46633));
    CascadeMux I__10850 (
            .O(N__46655),
            .I(N__46627));
    LocalMux I__10849 (
            .O(N__46652),
            .I(N__46624));
    LocalMux I__10848 (
            .O(N__46649),
            .I(N__46619));
    LocalMux I__10847 (
            .O(N__46646),
            .I(N__46619));
    CascadeMux I__10846 (
            .O(N__46645),
            .I(N__46616));
    InMux I__10845 (
            .O(N__46644),
            .I(N__46613));
    InMux I__10844 (
            .O(N__46643),
            .I(N__46610));
    InMux I__10843 (
            .O(N__46642),
            .I(N__46605));
    InMux I__10842 (
            .O(N__46639),
            .I(N__46605));
    Span4Mux_v I__10841 (
            .O(N__46636),
            .I(N__46602));
    LocalMux I__10840 (
            .O(N__46633),
            .I(N__46598));
    InMux I__10839 (
            .O(N__46632),
            .I(N__46593));
    InMux I__10838 (
            .O(N__46631),
            .I(N__46593));
    InMux I__10837 (
            .O(N__46630),
            .I(N__46590));
    InMux I__10836 (
            .O(N__46627),
            .I(N__46586));
    Span4Mux_v I__10835 (
            .O(N__46624),
            .I(N__46577));
    Span4Mux_v I__10834 (
            .O(N__46619),
            .I(N__46577));
    InMux I__10833 (
            .O(N__46616),
            .I(N__46574));
    LocalMux I__10832 (
            .O(N__46613),
            .I(N__46567));
    LocalMux I__10831 (
            .O(N__46610),
            .I(N__46567));
    LocalMux I__10830 (
            .O(N__46605),
            .I(N__46567));
    Span4Mux_h I__10829 (
            .O(N__46602),
            .I(N__46564));
    InMux I__10828 (
            .O(N__46601),
            .I(N__46561));
    Span4Mux_v I__10827 (
            .O(N__46598),
            .I(N__46554));
    LocalMux I__10826 (
            .O(N__46593),
            .I(N__46554));
    LocalMux I__10825 (
            .O(N__46590),
            .I(N__46554));
    InMux I__10824 (
            .O(N__46589),
            .I(N__46551));
    LocalMux I__10823 (
            .O(N__46586),
            .I(N__46548));
    InMux I__10822 (
            .O(N__46585),
            .I(N__46545));
    InMux I__10821 (
            .O(N__46584),
            .I(N__46542));
    InMux I__10820 (
            .O(N__46583),
            .I(N__46539));
    CascadeMux I__10819 (
            .O(N__46582),
            .I(N__46535));
    Span4Mux_h I__10818 (
            .O(N__46577),
            .I(N__46532));
    LocalMux I__10817 (
            .O(N__46574),
            .I(N__46523));
    Span4Mux_v I__10816 (
            .O(N__46567),
            .I(N__46523));
    Span4Mux_h I__10815 (
            .O(N__46564),
            .I(N__46523));
    LocalMux I__10814 (
            .O(N__46561),
            .I(N__46523));
    Span4Mux_v I__10813 (
            .O(N__46554),
            .I(N__46518));
    LocalMux I__10812 (
            .O(N__46551),
            .I(N__46518));
    Span4Mux_v I__10811 (
            .O(N__46548),
            .I(N__46509));
    LocalMux I__10810 (
            .O(N__46545),
            .I(N__46509));
    LocalMux I__10809 (
            .O(N__46542),
            .I(N__46509));
    LocalMux I__10808 (
            .O(N__46539),
            .I(N__46509));
    InMux I__10807 (
            .O(N__46538),
            .I(N__46506));
    InMux I__10806 (
            .O(N__46535),
            .I(N__46503));
    Span4Mux_v I__10805 (
            .O(N__46532),
            .I(N__46500));
    Span4Mux_v I__10804 (
            .O(N__46523),
            .I(N__46497));
    Span4Mux_h I__10803 (
            .O(N__46518),
            .I(N__46490));
    Span4Mux_v I__10802 (
            .O(N__46509),
            .I(N__46490));
    LocalMux I__10801 (
            .O(N__46506),
            .I(N__46490));
    LocalMux I__10800 (
            .O(N__46503),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__10799 (
            .O(N__46500),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__10798 (
            .O(N__46497),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    Odrv4 I__10797 (
            .O(N__46490),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ));
    CascadeMux I__10796 (
            .O(N__46481),
            .I(\ppm_encoder_1.N_290_cascade_ ));
    InMux I__10795 (
            .O(N__46478),
            .I(N__46469));
    InMux I__10794 (
            .O(N__46477),
            .I(N__46469));
    InMux I__10793 (
            .O(N__46476),
            .I(N__46469));
    LocalMux I__10792 (
            .O(N__46469),
            .I(\ppm_encoder_1.aileronZ0Z_4 ));
    InMux I__10791 (
            .O(N__46466),
            .I(N__46463));
    LocalMux I__10790 (
            .O(N__46463),
            .I(N__46460));
    Odrv12 I__10789 (
            .O(N__46460),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ));
    InMux I__10788 (
            .O(N__46457),
            .I(N__46454));
    LocalMux I__10787 (
            .O(N__46454),
            .I(N__46451));
    Span4Mux_v I__10786 (
            .O(N__46451),
            .I(N__46448));
    Span4Mux_h I__10785 (
            .O(N__46448),
            .I(N__46445));
    Odrv4 I__10784 (
            .O(N__46445),
            .I(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ));
    InMux I__10783 (
            .O(N__46442),
            .I(N__46439));
    LocalMux I__10782 (
            .O(N__46439),
            .I(N__46435));
    InMux I__10781 (
            .O(N__46438),
            .I(N__46432));
    Span4Mux_v I__10780 (
            .O(N__46435),
            .I(N__46429));
    LocalMux I__10779 (
            .O(N__46432),
            .I(N__46426));
    Span4Mux_h I__10778 (
            .O(N__46429),
            .I(N__46423));
    Span4Mux_v I__10777 (
            .O(N__46426),
            .I(N__46420));
    Odrv4 I__10776 (
            .O(N__46423),
            .I(throttle_order_4));
    Odrv4 I__10775 (
            .O(N__46420),
            .I(throttle_order_4));
    InMux I__10774 (
            .O(N__46415),
            .I(N__46410));
    InMux I__10773 (
            .O(N__46414),
            .I(N__46405));
    InMux I__10772 (
            .O(N__46413),
            .I(N__46405));
    LocalMux I__10771 (
            .O(N__46410),
            .I(N__46402));
    LocalMux I__10770 (
            .O(N__46405),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    Odrv4 I__10769 (
            .O(N__46402),
            .I(\ppm_encoder_1.throttleZ0Z_4 ));
    CascadeMux I__10768 (
            .O(N__46397),
            .I(N__46391));
    CascadeMux I__10767 (
            .O(N__46396),
            .I(N__46383));
    CascadeMux I__10766 (
            .O(N__46395),
            .I(N__46380));
    CascadeMux I__10765 (
            .O(N__46394),
            .I(N__46377));
    InMux I__10764 (
            .O(N__46391),
            .I(N__46371));
    CascadeMux I__10763 (
            .O(N__46390),
            .I(N__46368));
    CascadeMux I__10762 (
            .O(N__46389),
            .I(N__46362));
    CascadeMux I__10761 (
            .O(N__46388),
            .I(N__46359));
    CascadeMux I__10760 (
            .O(N__46387),
            .I(N__46356));
    InMux I__10759 (
            .O(N__46386),
            .I(N__46351));
    InMux I__10758 (
            .O(N__46383),
            .I(N__46351));
    InMux I__10757 (
            .O(N__46380),
            .I(N__46348));
    InMux I__10756 (
            .O(N__46377),
            .I(N__46343));
    InMux I__10755 (
            .O(N__46376),
            .I(N__46343));
    CascadeMux I__10754 (
            .O(N__46375),
            .I(N__46337));
    CascadeMux I__10753 (
            .O(N__46374),
            .I(N__46334));
    LocalMux I__10752 (
            .O(N__46371),
            .I(N__46329));
    InMux I__10751 (
            .O(N__46368),
            .I(N__46325));
    CascadeMux I__10750 (
            .O(N__46367),
            .I(N__46322));
    InMux I__10749 (
            .O(N__46366),
            .I(N__46312));
    InMux I__10748 (
            .O(N__46365),
            .I(N__46312));
    InMux I__10747 (
            .O(N__46362),
            .I(N__46312));
    InMux I__10746 (
            .O(N__46359),
            .I(N__46312));
    InMux I__10745 (
            .O(N__46356),
            .I(N__46301));
    LocalMux I__10744 (
            .O(N__46351),
            .I(N__46294));
    LocalMux I__10743 (
            .O(N__46348),
            .I(N__46294));
    LocalMux I__10742 (
            .O(N__46343),
            .I(N__46294));
    InMux I__10741 (
            .O(N__46342),
            .I(N__46279));
    InMux I__10740 (
            .O(N__46341),
            .I(N__46279));
    InMux I__10739 (
            .O(N__46340),
            .I(N__46279));
    InMux I__10738 (
            .O(N__46337),
            .I(N__46279));
    InMux I__10737 (
            .O(N__46334),
            .I(N__46279));
    InMux I__10736 (
            .O(N__46333),
            .I(N__46279));
    InMux I__10735 (
            .O(N__46332),
            .I(N__46279));
    Span4Mux_h I__10734 (
            .O(N__46329),
            .I(N__46276));
    InMux I__10733 (
            .O(N__46328),
            .I(N__46273));
    LocalMux I__10732 (
            .O(N__46325),
            .I(N__46270));
    InMux I__10731 (
            .O(N__46322),
            .I(N__46265));
    InMux I__10730 (
            .O(N__46321),
            .I(N__46265));
    LocalMux I__10729 (
            .O(N__46312),
            .I(N__46262));
    InMux I__10728 (
            .O(N__46311),
            .I(N__46257));
    InMux I__10727 (
            .O(N__46310),
            .I(N__46257));
    CascadeMux I__10726 (
            .O(N__46309),
            .I(N__46252));
    CascadeMux I__10725 (
            .O(N__46308),
            .I(N__46249));
    CascadeMux I__10724 (
            .O(N__46307),
            .I(N__46245));
    CascadeMux I__10723 (
            .O(N__46306),
            .I(N__46239));
    CascadeMux I__10722 (
            .O(N__46305),
            .I(N__46236));
    CascadeMux I__10721 (
            .O(N__46304),
            .I(N__46233));
    LocalMux I__10720 (
            .O(N__46301),
            .I(N__46230));
    Span4Mux_v I__10719 (
            .O(N__46294),
            .I(N__46221));
    LocalMux I__10718 (
            .O(N__46279),
            .I(N__46221));
    Span4Mux_v I__10717 (
            .O(N__46276),
            .I(N__46221));
    LocalMux I__10716 (
            .O(N__46273),
            .I(N__46221));
    Span4Mux_h I__10715 (
            .O(N__46270),
            .I(N__46212));
    LocalMux I__10714 (
            .O(N__46265),
            .I(N__46212));
    Span4Mux_h I__10713 (
            .O(N__46262),
            .I(N__46212));
    LocalMux I__10712 (
            .O(N__46257),
            .I(N__46212));
    InMux I__10711 (
            .O(N__46256),
            .I(N__46209));
    InMux I__10710 (
            .O(N__46255),
            .I(N__46200));
    InMux I__10709 (
            .O(N__46252),
            .I(N__46200));
    InMux I__10708 (
            .O(N__46249),
            .I(N__46200));
    InMux I__10707 (
            .O(N__46248),
            .I(N__46200));
    InMux I__10706 (
            .O(N__46245),
            .I(N__46195));
    InMux I__10705 (
            .O(N__46244),
            .I(N__46195));
    InMux I__10704 (
            .O(N__46243),
            .I(N__46176));
    InMux I__10703 (
            .O(N__46242),
            .I(N__46176));
    InMux I__10702 (
            .O(N__46239),
            .I(N__46176));
    InMux I__10701 (
            .O(N__46236),
            .I(N__46176));
    InMux I__10700 (
            .O(N__46233),
            .I(N__46176));
    Span4Mux_v I__10699 (
            .O(N__46230),
            .I(N__46171));
    Span4Mux_v I__10698 (
            .O(N__46221),
            .I(N__46171));
    Span4Mux_v I__10697 (
            .O(N__46212),
            .I(N__46161));
    LocalMux I__10696 (
            .O(N__46209),
            .I(N__46161));
    LocalMux I__10695 (
            .O(N__46200),
            .I(N__46161));
    LocalMux I__10694 (
            .O(N__46195),
            .I(N__46161));
    InMux I__10693 (
            .O(N__46194),
            .I(N__46158));
    CascadeMux I__10692 (
            .O(N__46193),
            .I(N__46152));
    CascadeMux I__10691 (
            .O(N__46192),
            .I(N__46148));
    CascadeMux I__10690 (
            .O(N__46191),
            .I(N__46145));
    InMux I__10689 (
            .O(N__46190),
            .I(N__46141));
    CascadeMux I__10688 (
            .O(N__46189),
            .I(N__46137));
    CascadeMux I__10687 (
            .O(N__46188),
            .I(N__46134));
    CascadeMux I__10686 (
            .O(N__46187),
            .I(N__46131));
    LocalMux I__10685 (
            .O(N__46176),
            .I(N__46128));
    Span4Mux_h I__10684 (
            .O(N__46171),
            .I(N__46125));
    CascadeMux I__10683 (
            .O(N__46170),
            .I(N__46122));
    Span4Mux_v I__10682 (
            .O(N__46161),
            .I(N__46119));
    LocalMux I__10681 (
            .O(N__46158),
            .I(N__46116));
    InMux I__10680 (
            .O(N__46157),
            .I(N__46113));
    InMux I__10679 (
            .O(N__46156),
            .I(N__46106));
    InMux I__10678 (
            .O(N__46155),
            .I(N__46106));
    InMux I__10677 (
            .O(N__46152),
            .I(N__46106));
    InMux I__10676 (
            .O(N__46151),
            .I(N__46097));
    InMux I__10675 (
            .O(N__46148),
            .I(N__46097));
    InMux I__10674 (
            .O(N__46145),
            .I(N__46097));
    InMux I__10673 (
            .O(N__46144),
            .I(N__46097));
    LocalMux I__10672 (
            .O(N__46141),
            .I(N__46094));
    InMux I__10671 (
            .O(N__46140),
            .I(N__46085));
    InMux I__10670 (
            .O(N__46137),
            .I(N__46085));
    InMux I__10669 (
            .O(N__46134),
            .I(N__46085));
    InMux I__10668 (
            .O(N__46131),
            .I(N__46085));
    Span4Mux_v I__10667 (
            .O(N__46128),
            .I(N__46082));
    Span4Mux_h I__10666 (
            .O(N__46125),
            .I(N__46079));
    InMux I__10665 (
            .O(N__46122),
            .I(N__46076));
    Span4Mux_h I__10664 (
            .O(N__46119),
            .I(N__46069));
    Span4Mux_v I__10663 (
            .O(N__46116),
            .I(N__46069));
    LocalMux I__10662 (
            .O(N__46113),
            .I(N__46069));
    LocalMux I__10661 (
            .O(N__46106),
            .I(N__46062));
    LocalMux I__10660 (
            .O(N__46097),
            .I(N__46062));
    Sp12to4 I__10659 (
            .O(N__46094),
            .I(N__46062));
    LocalMux I__10658 (
            .O(N__46085),
            .I(N__46059));
    Span4Mux_h I__10657 (
            .O(N__46082),
            .I(N__46054));
    Span4Mux_v I__10656 (
            .O(N__46079),
            .I(N__46054));
    LocalMux I__10655 (
            .O(N__46076),
            .I(N__46049));
    Span4Mux_v I__10654 (
            .O(N__46069),
            .I(N__46049));
    Span12Mux_v I__10653 (
            .O(N__46062),
            .I(N__46046));
    Span4Mux_v I__10652 (
            .O(N__46059),
            .I(N__46041));
    Span4Mux_v I__10651 (
            .O(N__46054),
            .I(N__46041));
    Span4Mux_v I__10650 (
            .O(N__46049),
            .I(N__46038));
    Odrv12 I__10649 (
            .O(N__46046),
            .I(pid_altitude_dv));
    Odrv4 I__10648 (
            .O(N__46041),
            .I(pid_altitude_dv));
    Odrv4 I__10647 (
            .O(N__46038),
            .I(pid_altitude_dv));
    InMux I__10646 (
            .O(N__46031),
            .I(N__46027));
    CascadeMux I__10645 (
            .O(N__46030),
            .I(N__46023));
    LocalMux I__10644 (
            .O(N__46027),
            .I(N__46020));
    InMux I__10643 (
            .O(N__46026),
            .I(N__46017));
    InMux I__10642 (
            .O(N__46023),
            .I(N__46014));
    Span4Mux_v I__10641 (
            .O(N__46020),
            .I(N__46011));
    LocalMux I__10640 (
            .O(N__46017),
            .I(N__46008));
    LocalMux I__10639 (
            .O(N__46014),
            .I(side_order_0));
    Odrv4 I__10638 (
            .O(N__46011),
            .I(side_order_0));
    Odrv4 I__10637 (
            .O(N__46008),
            .I(side_order_0));
    InMux I__10636 (
            .O(N__46001),
            .I(N__45998));
    LocalMux I__10635 (
            .O(N__45998),
            .I(N__45994));
    InMux I__10634 (
            .O(N__45997),
            .I(N__45990));
    Span4Mux_v I__10633 (
            .O(N__45994),
            .I(N__45987));
    InMux I__10632 (
            .O(N__45993),
            .I(N__45984));
    LocalMux I__10631 (
            .O(N__45990),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    Odrv4 I__10630 (
            .O(N__45987),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    LocalMux I__10629 (
            .O(N__45984),
            .I(\ppm_encoder_1.aileronZ0Z_0 ));
    InMux I__10628 (
            .O(N__45977),
            .I(N__45974));
    LocalMux I__10627 (
            .O(N__45974),
            .I(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ));
    InMux I__10626 (
            .O(N__45971),
            .I(N__45968));
    LocalMux I__10625 (
            .O(N__45968),
            .I(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ));
    InMux I__10624 (
            .O(N__45965),
            .I(N__45961));
    CascadeMux I__10623 (
            .O(N__45964),
            .I(N__45958));
    LocalMux I__10622 (
            .O(N__45961),
            .I(N__45955));
    InMux I__10621 (
            .O(N__45958),
            .I(N__45951));
    Span4Mux_v I__10620 (
            .O(N__45955),
            .I(N__45948));
    InMux I__10619 (
            .O(N__45954),
            .I(N__45945));
    LocalMux I__10618 (
            .O(N__45951),
            .I(N__45940));
    Span4Mux_h I__10617 (
            .O(N__45948),
            .I(N__45940));
    LocalMux I__10616 (
            .O(N__45945),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    Odrv4 I__10615 (
            .O(N__45940),
            .I(\ppm_encoder_1.rudderZ0Z_7 ));
    CascadeMux I__10614 (
            .O(N__45935),
            .I(N__45929));
    CascadeMux I__10613 (
            .O(N__45934),
            .I(N__45926));
    InMux I__10612 (
            .O(N__45933),
            .I(N__45921));
    CascadeMux I__10611 (
            .O(N__45932),
            .I(N__45918));
    InMux I__10610 (
            .O(N__45929),
            .I(N__45915));
    InMux I__10609 (
            .O(N__45926),
            .I(N__45912));
    InMux I__10608 (
            .O(N__45925),
            .I(N__45909));
    InMux I__10607 (
            .O(N__45924),
            .I(N__45906));
    LocalMux I__10606 (
            .O(N__45921),
            .I(N__45902));
    InMux I__10605 (
            .O(N__45918),
            .I(N__45899));
    LocalMux I__10604 (
            .O(N__45915),
            .I(N__45894));
    LocalMux I__10603 (
            .O(N__45912),
            .I(N__45891));
    LocalMux I__10602 (
            .O(N__45909),
            .I(N__45884));
    LocalMux I__10601 (
            .O(N__45906),
            .I(N__45884));
    InMux I__10600 (
            .O(N__45905),
            .I(N__45881));
    Span4Mux_h I__10599 (
            .O(N__45902),
            .I(N__45876));
    LocalMux I__10598 (
            .O(N__45899),
            .I(N__45876));
    InMux I__10597 (
            .O(N__45898),
            .I(N__45873));
    InMux I__10596 (
            .O(N__45897),
            .I(N__45870));
    Span4Mux_v I__10595 (
            .O(N__45894),
            .I(N__45865));
    Span4Mux_v I__10594 (
            .O(N__45891),
            .I(N__45865));
    InMux I__10593 (
            .O(N__45890),
            .I(N__45862));
    InMux I__10592 (
            .O(N__45889),
            .I(N__45859));
    Odrv4 I__10591 (
            .O(N__45884),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__10590 (
            .O(N__45881),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__10589 (
            .O(N__45876),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__10588 (
            .O(N__45873),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__10587 (
            .O(N__45870),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    Odrv4 I__10586 (
            .O(N__45865),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__10585 (
            .O(N__45862),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    LocalMux I__10584 (
            .O(N__45859),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ));
    CascadeMux I__10583 (
            .O(N__45842),
            .I(N__45836));
    CascadeMux I__10582 (
            .O(N__45841),
            .I(N__45833));
    CascadeMux I__10581 (
            .O(N__45840),
            .I(N__45826));
    InMux I__10580 (
            .O(N__45839),
            .I(N__45823));
    InMux I__10579 (
            .O(N__45836),
            .I(N__45820));
    InMux I__10578 (
            .O(N__45833),
            .I(N__45817));
    CascadeMux I__10577 (
            .O(N__45832),
            .I(N__45814));
    CascadeMux I__10576 (
            .O(N__45831),
            .I(N__45810));
    InMux I__10575 (
            .O(N__45830),
            .I(N__45807));
    InMux I__10574 (
            .O(N__45829),
            .I(N__45804));
    InMux I__10573 (
            .O(N__45826),
            .I(N__45799));
    LocalMux I__10572 (
            .O(N__45823),
            .I(N__45796));
    LocalMux I__10571 (
            .O(N__45820),
            .I(N__45793));
    LocalMux I__10570 (
            .O(N__45817),
            .I(N__45790));
    InMux I__10569 (
            .O(N__45814),
            .I(N__45787));
    CascadeMux I__10568 (
            .O(N__45813),
            .I(N__45782));
    InMux I__10567 (
            .O(N__45810),
            .I(N__45779));
    LocalMux I__10566 (
            .O(N__45807),
            .I(N__45774));
    LocalMux I__10565 (
            .O(N__45804),
            .I(N__45774));
    InMux I__10564 (
            .O(N__45803),
            .I(N__45771));
    InMux I__10563 (
            .O(N__45802),
            .I(N__45768));
    LocalMux I__10562 (
            .O(N__45799),
            .I(N__45765));
    Span4Mux_v I__10561 (
            .O(N__45796),
            .I(N__45756));
    Span4Mux_v I__10560 (
            .O(N__45793),
            .I(N__45756));
    Span4Mux_v I__10559 (
            .O(N__45790),
            .I(N__45756));
    LocalMux I__10558 (
            .O(N__45787),
            .I(N__45756));
    InMux I__10557 (
            .O(N__45786),
            .I(N__45753));
    InMux I__10556 (
            .O(N__45785),
            .I(N__45748));
    InMux I__10555 (
            .O(N__45782),
            .I(N__45748));
    LocalMux I__10554 (
            .O(N__45779),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__10553 (
            .O(N__45774),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__10552 (
            .O(N__45771),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__10551 (
            .O(N__45768),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__10550 (
            .O(N__45765),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    Odrv4 I__10549 (
            .O(N__45756),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__10548 (
            .O(N__45753),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    LocalMux I__10547 (
            .O(N__45748),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ));
    InMux I__10546 (
            .O(N__45731),
            .I(N__45728));
    LocalMux I__10545 (
            .O(N__45728),
            .I(N__45724));
    InMux I__10544 (
            .O(N__45727),
            .I(N__45721));
    Span4Mux_v I__10543 (
            .O(N__45724),
            .I(N__45718));
    LocalMux I__10542 (
            .O(N__45721),
            .I(N__45715));
    Odrv4 I__10541 (
            .O(N__45718),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    Odrv4 I__10540 (
            .O(N__45715),
            .I(\ppm_encoder_1.un1_init_pulses_0_7 ));
    CascadeMux I__10539 (
            .O(N__45710),
            .I(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ));
    CascadeMux I__10538 (
            .O(N__45707),
            .I(N__45704));
    InMux I__10537 (
            .O(N__45704),
            .I(N__45701));
    LocalMux I__10536 (
            .O(N__45701),
            .I(N__45698));
    Span4Mux_h I__10535 (
            .O(N__45698),
            .I(N__45695));
    Odrv4 I__10534 (
            .O(N__45695),
            .I(\ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ));
    InMux I__10533 (
            .O(N__45692),
            .I(N__45689));
    LocalMux I__10532 (
            .O(N__45689),
            .I(\ppm_encoder_1.un2_throttle_iv_1_7 ));
    CascadeMux I__10531 (
            .O(N__45686),
            .I(\ppm_encoder_1.N_293_cascade_ ));
    InMux I__10530 (
            .O(N__45683),
            .I(N__45680));
    LocalMux I__10529 (
            .O(N__45680),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ));
    InMux I__10528 (
            .O(N__45677),
            .I(N__45674));
    LocalMux I__10527 (
            .O(N__45674),
            .I(N__45671));
    Span4Mux_h I__10526 (
            .O(N__45671),
            .I(N__45668));
    Span4Mux_h I__10525 (
            .O(N__45668),
            .I(N__45665));
    Odrv4 I__10524 (
            .O(N__45665),
            .I(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ));
    CascadeMux I__10523 (
            .O(N__45662),
            .I(N__45659));
    InMux I__10522 (
            .O(N__45659),
            .I(N__45655));
    CascadeMux I__10521 (
            .O(N__45658),
            .I(N__45651));
    LocalMux I__10520 (
            .O(N__45655),
            .I(N__45648));
    InMux I__10519 (
            .O(N__45654),
            .I(N__45645));
    InMux I__10518 (
            .O(N__45651),
            .I(N__45642));
    Span12Mux_s11_h I__10517 (
            .O(N__45648),
            .I(N__45639));
    LocalMux I__10516 (
            .O(N__45645),
            .I(N__45636));
    LocalMux I__10515 (
            .O(N__45642),
            .I(side_order_7));
    Odrv12 I__10514 (
            .O(N__45639),
            .I(side_order_7));
    Odrv4 I__10513 (
            .O(N__45636),
            .I(side_order_7));
    InMux I__10512 (
            .O(N__45629),
            .I(N__45620));
    InMux I__10511 (
            .O(N__45628),
            .I(N__45620));
    InMux I__10510 (
            .O(N__45627),
            .I(N__45620));
    LocalMux I__10509 (
            .O(N__45620),
            .I(\ppm_encoder_1.aileronZ0Z_7 ));
    InMux I__10508 (
            .O(N__45617),
            .I(N__45614));
    LocalMux I__10507 (
            .O(N__45614),
            .I(N__45611));
    Span4Mux_h I__10506 (
            .O(N__45611),
            .I(N__45608));
    Odrv4 I__10505 (
            .O(N__45608),
            .I(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ));
    InMux I__10504 (
            .O(N__45605),
            .I(N__45602));
    LocalMux I__10503 (
            .O(N__45602),
            .I(N__45598));
    CascadeMux I__10502 (
            .O(N__45601),
            .I(N__45594));
    Span4Mux_h I__10501 (
            .O(N__45598),
            .I(N__45591));
    InMux I__10500 (
            .O(N__45597),
            .I(N__45588));
    InMux I__10499 (
            .O(N__45594),
            .I(N__45585));
    Span4Mux_h I__10498 (
            .O(N__45591),
            .I(N__45582));
    LocalMux I__10497 (
            .O(N__45588),
            .I(N__45579));
    LocalMux I__10496 (
            .O(N__45585),
            .I(front_order_7));
    Odrv4 I__10495 (
            .O(N__45582),
            .I(front_order_7));
    Odrv4 I__10494 (
            .O(N__45579),
            .I(front_order_7));
    InMux I__10493 (
            .O(N__45572),
            .I(N__45563));
    InMux I__10492 (
            .O(N__45571),
            .I(N__45563));
    InMux I__10491 (
            .O(N__45570),
            .I(N__45563));
    LocalMux I__10490 (
            .O(N__45563),
            .I(\ppm_encoder_1.elevatorZ0Z_7 ));
    InMux I__10489 (
            .O(N__45560),
            .I(N__45557));
    LocalMux I__10488 (
            .O(N__45557),
            .I(N__45554));
    Span4Mux_v I__10487 (
            .O(N__45554),
            .I(N__45551));
    Span4Mux_h I__10486 (
            .O(N__45551),
            .I(N__45548));
    Odrv4 I__10485 (
            .O(N__45548),
            .I(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ));
    CascadeMux I__10484 (
            .O(N__45545),
            .I(N__45541));
    CascadeMux I__10483 (
            .O(N__45544),
            .I(N__45538));
    InMux I__10482 (
            .O(N__45541),
            .I(N__45535));
    InMux I__10481 (
            .O(N__45538),
            .I(N__45531));
    LocalMux I__10480 (
            .O(N__45535),
            .I(N__45528));
    InMux I__10479 (
            .O(N__45534),
            .I(N__45525));
    LocalMux I__10478 (
            .O(N__45531),
            .I(N__45520));
    Span4Mux_h I__10477 (
            .O(N__45528),
            .I(N__45520));
    LocalMux I__10476 (
            .O(N__45525),
            .I(N__45517));
    Odrv4 I__10475 (
            .O(N__45520),
            .I(throttle_order_7));
    Odrv12 I__10474 (
            .O(N__45517),
            .I(throttle_order_7));
    InMux I__10473 (
            .O(N__45512),
            .I(N__45503));
    InMux I__10472 (
            .O(N__45511),
            .I(N__45503));
    InMux I__10471 (
            .O(N__45510),
            .I(N__45503));
    LocalMux I__10470 (
            .O(N__45503),
            .I(\ppm_encoder_1.throttleZ0Z_7 ));
    InMux I__10469 (
            .O(N__45500),
            .I(N__45495));
    CascadeMux I__10468 (
            .O(N__45499),
            .I(N__45491));
    CascadeMux I__10467 (
            .O(N__45498),
            .I(N__45488));
    LocalMux I__10466 (
            .O(N__45495),
            .I(N__45485));
    CascadeMux I__10465 (
            .O(N__45494),
            .I(N__45482));
    InMux I__10464 (
            .O(N__45491),
            .I(N__45479));
    InMux I__10463 (
            .O(N__45488),
            .I(N__45473));
    Span4Mux_h I__10462 (
            .O(N__45485),
            .I(N__45470));
    InMux I__10461 (
            .O(N__45482),
            .I(N__45467));
    LocalMux I__10460 (
            .O(N__45479),
            .I(N__45464));
    InMux I__10459 (
            .O(N__45478),
            .I(N__45461));
    InMux I__10458 (
            .O(N__45477),
            .I(N__45458));
    InMux I__10457 (
            .O(N__45476),
            .I(N__45455));
    LocalMux I__10456 (
            .O(N__45473),
            .I(N__45449));
    Span4Mux_v I__10455 (
            .O(N__45470),
            .I(N__45444));
    LocalMux I__10454 (
            .O(N__45467),
            .I(N__45441));
    Span4Mux_v I__10453 (
            .O(N__45464),
            .I(N__45435));
    LocalMux I__10452 (
            .O(N__45461),
            .I(N__45435));
    LocalMux I__10451 (
            .O(N__45458),
            .I(N__45430));
    LocalMux I__10450 (
            .O(N__45455),
            .I(N__45430));
    InMux I__10449 (
            .O(N__45454),
            .I(N__45425));
    InMux I__10448 (
            .O(N__45453),
            .I(N__45425));
    CascadeMux I__10447 (
            .O(N__45452),
            .I(N__45419));
    Span4Mux_h I__10446 (
            .O(N__45449),
            .I(N__45416));
    InMux I__10445 (
            .O(N__45448),
            .I(N__45411));
    InMux I__10444 (
            .O(N__45447),
            .I(N__45411));
    Span4Mux_h I__10443 (
            .O(N__45444),
            .I(N__45406));
    Span4Mux_h I__10442 (
            .O(N__45441),
            .I(N__45406));
    InMux I__10441 (
            .O(N__45440),
            .I(N__45403));
    Span4Mux_h I__10440 (
            .O(N__45435),
            .I(N__45396));
    Span4Mux_h I__10439 (
            .O(N__45430),
            .I(N__45396));
    LocalMux I__10438 (
            .O(N__45425),
            .I(N__45396));
    InMux I__10437 (
            .O(N__45424),
            .I(N__45393));
    InMux I__10436 (
            .O(N__45423),
            .I(N__45388));
    InMux I__10435 (
            .O(N__45422),
            .I(N__45388));
    InMux I__10434 (
            .O(N__45419),
            .I(N__45385));
    Odrv4 I__10433 (
            .O(N__45416),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__10432 (
            .O(N__45411),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__10431 (
            .O(N__45406),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__10430 (
            .O(N__45403),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    Odrv4 I__10429 (
            .O(N__45396),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__10428 (
            .O(N__45393),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__10427 (
            .O(N__45388),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    LocalMux I__10426 (
            .O(N__45385),
            .I(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ));
    CascadeMux I__10425 (
            .O(N__45368),
            .I(N__45363));
    InMux I__10424 (
            .O(N__45367),
            .I(N__45357));
    InMux I__10423 (
            .O(N__45366),
            .I(N__45354));
    InMux I__10422 (
            .O(N__45363),
            .I(N__45349));
    CascadeMux I__10421 (
            .O(N__45362),
            .I(N__45346));
    CascadeMux I__10420 (
            .O(N__45361),
            .I(N__45343));
    CascadeMux I__10419 (
            .O(N__45360),
            .I(N__45340));
    LocalMux I__10418 (
            .O(N__45357),
            .I(N__45333));
    LocalMux I__10417 (
            .O(N__45354),
            .I(N__45333));
    InMux I__10416 (
            .O(N__45353),
            .I(N__45330));
    InMux I__10415 (
            .O(N__45352),
            .I(N__45327));
    LocalMux I__10414 (
            .O(N__45349),
            .I(N__45324));
    InMux I__10413 (
            .O(N__45346),
            .I(N__45321));
    InMux I__10412 (
            .O(N__45343),
            .I(N__45318));
    InMux I__10411 (
            .O(N__45340),
            .I(N__45315));
    CascadeMux I__10410 (
            .O(N__45339),
            .I(N__45311));
    CascadeMux I__10409 (
            .O(N__45338),
            .I(N__45305));
    Span4Mux_v I__10408 (
            .O(N__45333),
            .I(N__45299));
    LocalMux I__10407 (
            .O(N__45330),
            .I(N__45299));
    LocalMux I__10406 (
            .O(N__45327),
            .I(N__45288));
    Span4Mux_h I__10405 (
            .O(N__45324),
            .I(N__45288));
    LocalMux I__10404 (
            .O(N__45321),
            .I(N__45288));
    LocalMux I__10403 (
            .O(N__45318),
            .I(N__45288));
    LocalMux I__10402 (
            .O(N__45315),
            .I(N__45288));
    InMux I__10401 (
            .O(N__45314),
            .I(N__45285));
    InMux I__10400 (
            .O(N__45311),
            .I(N__45282));
    InMux I__10399 (
            .O(N__45310),
            .I(N__45277));
    InMux I__10398 (
            .O(N__45309),
            .I(N__45277));
    InMux I__10397 (
            .O(N__45308),
            .I(N__45274));
    InMux I__10396 (
            .O(N__45305),
            .I(N__45269));
    InMux I__10395 (
            .O(N__45304),
            .I(N__45269));
    Odrv4 I__10394 (
            .O(N__45299),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    Odrv4 I__10393 (
            .O(N__45288),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__10392 (
            .O(N__45285),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__10391 (
            .O(N__45282),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__10390 (
            .O(N__45277),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__10389 (
            .O(N__45274),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    LocalMux I__10388 (
            .O(N__45269),
            .I(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ));
    InMux I__10387 (
            .O(N__45254),
            .I(N__45250));
    CascadeMux I__10386 (
            .O(N__45253),
            .I(N__45247));
    LocalMux I__10385 (
            .O(N__45250),
            .I(N__45244));
    InMux I__10384 (
            .O(N__45247),
            .I(N__45241));
    Span4Mux_h I__10383 (
            .O(N__45244),
            .I(N__45237));
    LocalMux I__10382 (
            .O(N__45241),
            .I(N__45234));
    InMux I__10381 (
            .O(N__45240),
            .I(N__45231));
    Span4Mux_h I__10380 (
            .O(N__45237),
            .I(N__45226));
    Span4Mux_h I__10379 (
            .O(N__45234),
            .I(N__45226));
    LocalMux I__10378 (
            .O(N__45231),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    Odrv4 I__10377 (
            .O(N__45226),
            .I(\ppm_encoder_1.init_pulsesZ0Z_18 ));
    CascadeMux I__10376 (
            .O(N__45221),
            .I(N__45215));
    CascadeMux I__10375 (
            .O(N__45220),
            .I(N__45212));
    InMux I__10374 (
            .O(N__45219),
            .I(N__45202));
    InMux I__10373 (
            .O(N__45218),
            .I(N__45202));
    InMux I__10372 (
            .O(N__45215),
            .I(N__45202));
    InMux I__10371 (
            .O(N__45212),
            .I(N__45202));
    InMux I__10370 (
            .O(N__45211),
            .I(N__45199));
    LocalMux I__10369 (
            .O(N__45202),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ));
    LocalMux I__10368 (
            .O(N__45199),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ));
    CascadeMux I__10367 (
            .O(N__45194),
            .I(N__45191));
    InMux I__10366 (
            .O(N__45191),
            .I(N__45185));
    InMux I__10365 (
            .O(N__45190),
            .I(N__45185));
    LocalMux I__10364 (
            .O(N__45185),
            .I(\ppm_encoder_1.pulses2countZ0Z_18 ));
    InMux I__10363 (
            .O(N__45182),
            .I(N__45175));
    InMux I__10362 (
            .O(N__45181),
            .I(N__45175));
    InMux I__10361 (
            .O(N__45180),
            .I(N__45172));
    LocalMux I__10360 (
            .O(N__45175),
            .I(N__45169));
    LocalMux I__10359 (
            .O(N__45172),
            .I(N__45164));
    Span4Mux_v I__10358 (
            .O(N__45169),
            .I(N__45164));
    Odrv4 I__10357 (
            .O(N__45164),
            .I(\ppm_encoder_1.init_pulsesZ0Z_16 ));
    InMux I__10356 (
            .O(N__45161),
            .I(N__45153));
    CascadeMux I__10355 (
            .O(N__45160),
            .I(N__45149));
    CascadeMux I__10354 (
            .O(N__45159),
            .I(N__45145));
    CascadeMux I__10353 (
            .O(N__45158),
            .I(N__45141));
    CascadeMux I__10352 (
            .O(N__45157),
            .I(N__45137));
    InMux I__10351 (
            .O(N__45156),
            .I(N__45128));
    LocalMux I__10350 (
            .O(N__45153),
            .I(N__45118));
    InMux I__10349 (
            .O(N__45152),
            .I(N__45111));
    InMux I__10348 (
            .O(N__45149),
            .I(N__45111));
    InMux I__10347 (
            .O(N__45148),
            .I(N__45111));
    InMux I__10346 (
            .O(N__45145),
            .I(N__45106));
    InMux I__10345 (
            .O(N__45144),
            .I(N__45106));
    InMux I__10344 (
            .O(N__45141),
            .I(N__45101));
    InMux I__10343 (
            .O(N__45140),
            .I(N__45101));
    InMux I__10342 (
            .O(N__45137),
            .I(N__45092));
    InMux I__10341 (
            .O(N__45136),
            .I(N__45092));
    InMux I__10340 (
            .O(N__45135),
            .I(N__45092));
    InMux I__10339 (
            .O(N__45134),
            .I(N__45092));
    CascadeMux I__10338 (
            .O(N__45133),
            .I(N__45086));
    InMux I__10337 (
            .O(N__45132),
            .I(N__45082));
    CascadeMux I__10336 (
            .O(N__45131),
            .I(N__45079));
    LocalMux I__10335 (
            .O(N__45128),
            .I(N__45075));
    InMux I__10334 (
            .O(N__45127),
            .I(N__45066));
    InMux I__10333 (
            .O(N__45126),
            .I(N__45066));
    InMux I__10332 (
            .O(N__45125),
            .I(N__45066));
    InMux I__10331 (
            .O(N__45124),
            .I(N__45066));
    CascadeMux I__10330 (
            .O(N__45123),
            .I(N__45063));
    CascadeMux I__10329 (
            .O(N__45122),
            .I(N__45057));
    CascadeMux I__10328 (
            .O(N__45121),
            .I(N__45053));
    Span4Mux_h I__10327 (
            .O(N__45118),
            .I(N__45046));
    LocalMux I__10326 (
            .O(N__45111),
            .I(N__45046));
    LocalMux I__10325 (
            .O(N__45106),
            .I(N__45043));
    LocalMux I__10324 (
            .O(N__45101),
            .I(N__45038));
    LocalMux I__10323 (
            .O(N__45092),
            .I(N__45038));
    CascadeMux I__10322 (
            .O(N__45091),
            .I(N__45035));
    CascadeMux I__10321 (
            .O(N__45090),
            .I(N__45032));
    CascadeMux I__10320 (
            .O(N__45089),
            .I(N__45025));
    InMux I__10319 (
            .O(N__45086),
            .I(N__45020));
    InMux I__10318 (
            .O(N__45085),
            .I(N__45017));
    LocalMux I__10317 (
            .O(N__45082),
            .I(N__45014));
    InMux I__10316 (
            .O(N__45079),
            .I(N__45009));
    InMux I__10315 (
            .O(N__45078),
            .I(N__45009));
    Span4Mux_v I__10314 (
            .O(N__45075),
            .I(N__45004));
    LocalMux I__10313 (
            .O(N__45066),
            .I(N__45004));
    InMux I__10312 (
            .O(N__45063),
            .I(N__44995));
    InMux I__10311 (
            .O(N__45062),
            .I(N__44995));
    InMux I__10310 (
            .O(N__45061),
            .I(N__44995));
    InMux I__10309 (
            .O(N__45060),
            .I(N__44995));
    InMux I__10308 (
            .O(N__45057),
            .I(N__44984));
    InMux I__10307 (
            .O(N__45056),
            .I(N__44984));
    InMux I__10306 (
            .O(N__45053),
            .I(N__44984));
    InMux I__10305 (
            .O(N__45052),
            .I(N__44984));
    InMux I__10304 (
            .O(N__45051),
            .I(N__44984));
    Span4Mux_v I__10303 (
            .O(N__45046),
            .I(N__44977));
    Span4Mux_v I__10302 (
            .O(N__45043),
            .I(N__44977));
    Span4Mux_v I__10301 (
            .O(N__45038),
            .I(N__44977));
    InMux I__10300 (
            .O(N__45035),
            .I(N__44968));
    InMux I__10299 (
            .O(N__45032),
            .I(N__44968));
    InMux I__10298 (
            .O(N__45031),
            .I(N__44968));
    InMux I__10297 (
            .O(N__45030),
            .I(N__44968));
    InMux I__10296 (
            .O(N__45029),
            .I(N__44959));
    InMux I__10295 (
            .O(N__45028),
            .I(N__44959));
    InMux I__10294 (
            .O(N__45025),
            .I(N__44959));
    InMux I__10293 (
            .O(N__45024),
            .I(N__44959));
    InMux I__10292 (
            .O(N__45023),
            .I(N__44956));
    LocalMux I__10291 (
            .O(N__45020),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10290 (
            .O(N__45017),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10289 (
            .O(N__45014),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10288 (
            .O(N__45009),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10287 (
            .O(N__45004),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10286 (
            .O(N__44995),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10285 (
            .O(N__44984),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    Odrv4 I__10284 (
            .O(N__44977),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10283 (
            .O(N__44968),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10282 (
            .O(N__44959),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    LocalMux I__10281 (
            .O(N__44956),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ));
    CascadeMux I__10280 (
            .O(N__44933),
            .I(N__44927));
    InMux I__10279 (
            .O(N__44932),
            .I(N__44904));
    InMux I__10278 (
            .O(N__44931),
            .I(N__44904));
    CascadeMux I__10277 (
            .O(N__44930),
            .I(N__44901));
    InMux I__10276 (
            .O(N__44927),
            .I(N__44893));
    InMux I__10275 (
            .O(N__44926),
            .I(N__44888));
    InMux I__10274 (
            .O(N__44925),
            .I(N__44888));
    InMux I__10273 (
            .O(N__44924),
            .I(N__44879));
    InMux I__10272 (
            .O(N__44923),
            .I(N__44879));
    InMux I__10271 (
            .O(N__44922),
            .I(N__44879));
    InMux I__10270 (
            .O(N__44921),
            .I(N__44879));
    InMux I__10269 (
            .O(N__44920),
            .I(N__44874));
    InMux I__10268 (
            .O(N__44919),
            .I(N__44874));
    InMux I__10267 (
            .O(N__44918),
            .I(N__44865));
    InMux I__10266 (
            .O(N__44917),
            .I(N__44865));
    InMux I__10265 (
            .O(N__44916),
            .I(N__44865));
    InMux I__10264 (
            .O(N__44915),
            .I(N__44865));
    InMux I__10263 (
            .O(N__44914),
            .I(N__44862));
    CascadeMux I__10262 (
            .O(N__44913),
            .I(N__44854));
    CascadeMux I__10261 (
            .O(N__44912),
            .I(N__44836));
    InMux I__10260 (
            .O(N__44911),
            .I(N__44819));
    InMux I__10259 (
            .O(N__44910),
            .I(N__44819));
    InMux I__10258 (
            .O(N__44909),
            .I(N__44819));
    LocalMux I__10257 (
            .O(N__44904),
            .I(N__44816));
    InMux I__10256 (
            .O(N__44901),
            .I(N__44811));
    InMux I__10255 (
            .O(N__44900),
            .I(N__44811));
    InMux I__10254 (
            .O(N__44899),
            .I(N__44806));
    InMux I__10253 (
            .O(N__44898),
            .I(N__44806));
    InMux I__10252 (
            .O(N__44897),
            .I(N__44801));
    InMux I__10251 (
            .O(N__44896),
            .I(N__44801));
    LocalMux I__10250 (
            .O(N__44893),
            .I(N__44796));
    LocalMux I__10249 (
            .O(N__44888),
            .I(N__44796));
    LocalMux I__10248 (
            .O(N__44879),
            .I(N__44793));
    LocalMux I__10247 (
            .O(N__44874),
            .I(N__44788));
    LocalMux I__10246 (
            .O(N__44865),
            .I(N__44788));
    LocalMux I__10245 (
            .O(N__44862),
            .I(N__44783));
    InMux I__10244 (
            .O(N__44861),
            .I(N__44772));
    InMux I__10243 (
            .O(N__44860),
            .I(N__44772));
    InMux I__10242 (
            .O(N__44859),
            .I(N__44772));
    InMux I__10241 (
            .O(N__44858),
            .I(N__44772));
    InMux I__10240 (
            .O(N__44857),
            .I(N__44772));
    InMux I__10239 (
            .O(N__44854),
            .I(N__44757));
    InMux I__10238 (
            .O(N__44853),
            .I(N__44757));
    InMux I__10237 (
            .O(N__44852),
            .I(N__44757));
    InMux I__10236 (
            .O(N__44851),
            .I(N__44757));
    InMux I__10235 (
            .O(N__44850),
            .I(N__44757));
    InMux I__10234 (
            .O(N__44849),
            .I(N__44757));
    InMux I__10233 (
            .O(N__44848),
            .I(N__44757));
    InMux I__10232 (
            .O(N__44847),
            .I(N__44748));
    InMux I__10231 (
            .O(N__44846),
            .I(N__44748));
    InMux I__10230 (
            .O(N__44845),
            .I(N__44748));
    InMux I__10229 (
            .O(N__44844),
            .I(N__44748));
    InMux I__10228 (
            .O(N__44843),
            .I(N__44739));
    InMux I__10227 (
            .O(N__44842),
            .I(N__44739));
    InMux I__10226 (
            .O(N__44841),
            .I(N__44739));
    InMux I__10225 (
            .O(N__44840),
            .I(N__44739));
    InMux I__10224 (
            .O(N__44839),
            .I(N__44726));
    InMux I__10223 (
            .O(N__44836),
            .I(N__44726));
    InMux I__10222 (
            .O(N__44835),
            .I(N__44726));
    InMux I__10221 (
            .O(N__44834),
            .I(N__44726));
    InMux I__10220 (
            .O(N__44833),
            .I(N__44726));
    InMux I__10219 (
            .O(N__44832),
            .I(N__44726));
    InMux I__10218 (
            .O(N__44831),
            .I(N__44711));
    InMux I__10217 (
            .O(N__44830),
            .I(N__44711));
    InMux I__10216 (
            .O(N__44829),
            .I(N__44711));
    InMux I__10215 (
            .O(N__44828),
            .I(N__44711));
    InMux I__10214 (
            .O(N__44827),
            .I(N__44711));
    InMux I__10213 (
            .O(N__44826),
            .I(N__44708));
    LocalMux I__10212 (
            .O(N__44819),
            .I(N__44703));
    Span4Mux_v I__10211 (
            .O(N__44816),
            .I(N__44703));
    LocalMux I__10210 (
            .O(N__44811),
            .I(N__44700));
    LocalMux I__10209 (
            .O(N__44806),
            .I(N__44689));
    LocalMux I__10208 (
            .O(N__44801),
            .I(N__44689));
    Span4Mux_v I__10207 (
            .O(N__44796),
            .I(N__44689));
    Span4Mux_h I__10206 (
            .O(N__44793),
            .I(N__44689));
    Span4Mux_h I__10205 (
            .O(N__44788),
            .I(N__44689));
    InMux I__10204 (
            .O(N__44787),
            .I(N__44684));
    InMux I__10203 (
            .O(N__44786),
            .I(N__44684));
    Span4Mux_v I__10202 (
            .O(N__44783),
            .I(N__44679));
    LocalMux I__10201 (
            .O(N__44772),
            .I(N__44679));
    LocalMux I__10200 (
            .O(N__44757),
            .I(N__44670));
    LocalMux I__10199 (
            .O(N__44748),
            .I(N__44670));
    LocalMux I__10198 (
            .O(N__44739),
            .I(N__44670));
    LocalMux I__10197 (
            .O(N__44726),
            .I(N__44670));
    CascadeMux I__10196 (
            .O(N__44725),
            .I(N__44663));
    CascadeMux I__10195 (
            .O(N__44724),
            .I(N__44660));
    InMux I__10194 (
            .O(N__44723),
            .I(N__44655));
    InMux I__10193 (
            .O(N__44722),
            .I(N__44655));
    LocalMux I__10192 (
            .O(N__44711),
            .I(N__44652));
    LocalMux I__10191 (
            .O(N__44708),
            .I(N__44649));
    Span4Mux_v I__10190 (
            .O(N__44703),
            .I(N__44646));
    Span4Mux_h I__10189 (
            .O(N__44700),
            .I(N__44641));
    Span4Mux_v I__10188 (
            .O(N__44689),
            .I(N__44641));
    LocalMux I__10187 (
            .O(N__44684),
            .I(N__44634));
    Span4Mux_h I__10186 (
            .O(N__44679),
            .I(N__44634));
    Span4Mux_v I__10185 (
            .O(N__44670),
            .I(N__44634));
    InMux I__10184 (
            .O(N__44669),
            .I(N__44627));
    InMux I__10183 (
            .O(N__44668),
            .I(N__44627));
    InMux I__10182 (
            .O(N__44667),
            .I(N__44627));
    InMux I__10181 (
            .O(N__44666),
            .I(N__44624));
    InMux I__10180 (
            .O(N__44663),
            .I(N__44621));
    InMux I__10179 (
            .O(N__44660),
            .I(N__44618));
    LocalMux I__10178 (
            .O(N__44655),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10177 (
            .O(N__44652),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10176 (
            .O(N__44649),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10175 (
            .O(N__44646),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10174 (
            .O(N__44641),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    Odrv4 I__10173 (
            .O(N__44634),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10172 (
            .O(N__44627),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10171 (
            .O(N__44624),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10170 (
            .O(N__44621),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    LocalMux I__10169 (
            .O(N__44618),
            .I(\ppm_encoder_1.PPM_STATE_53_d ));
    InMux I__10168 (
            .O(N__44597),
            .I(N__44594));
    LocalMux I__10167 (
            .O(N__44594),
            .I(N__44591));
    Odrv4 I__10166 (
            .O(N__44591),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_16 ));
    InMux I__10165 (
            .O(N__44588),
            .I(N__44585));
    LocalMux I__10164 (
            .O(N__44585),
            .I(N__44582));
    Odrv12 I__10163 (
            .O(N__44582),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ));
    InMux I__10162 (
            .O(N__44579),
            .I(N__44576));
    LocalMux I__10161 (
            .O(N__44576),
            .I(N__44573));
    Span4Mux_v I__10160 (
            .O(N__44573),
            .I(N__44570));
    Span4Mux_h I__10159 (
            .O(N__44570),
            .I(N__44567));
    Odrv4 I__10158 (
            .O(N__44567),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ));
    InMux I__10157 (
            .O(N__44564),
            .I(N__44561));
    LocalMux I__10156 (
            .O(N__44561),
            .I(\ppm_encoder_1.pulses2countZ0Z_6 ));
    InMux I__10155 (
            .O(N__44558),
            .I(N__44555));
    LocalMux I__10154 (
            .O(N__44555),
            .I(N__44552));
    Span4Mux_v I__10153 (
            .O(N__44552),
            .I(N__44549));
    Span4Mux_h I__10152 (
            .O(N__44549),
            .I(N__44546));
    Odrv4 I__10151 (
            .O(N__44546),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ));
    CascadeMux I__10150 (
            .O(N__44543),
            .I(N__44540));
    InMux I__10149 (
            .O(N__44540),
            .I(N__44537));
    LocalMux I__10148 (
            .O(N__44537),
            .I(\ppm_encoder_1.pulses2countZ0Z_7 ));
    InMux I__10147 (
            .O(N__44534),
            .I(N__44531));
    LocalMux I__10146 (
            .O(N__44531),
            .I(N__44528));
    Span4Mux_h I__10145 (
            .O(N__44528),
            .I(N__44525));
    Odrv4 I__10144 (
            .O(N__44525),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ));
    InMux I__10143 (
            .O(N__44522),
            .I(N__44519));
    LocalMux I__10142 (
            .O(N__44519),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ));
    InMux I__10141 (
            .O(N__44516),
            .I(N__44513));
    LocalMux I__10140 (
            .O(N__44513),
            .I(N__44510));
    Span4Mux_v I__10139 (
            .O(N__44510),
            .I(N__44507));
    Odrv4 I__10138 (
            .O(N__44507),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ));
    CascadeMux I__10137 (
            .O(N__44504),
            .I(N__44495));
    InMux I__10136 (
            .O(N__44503),
            .I(N__44477));
    InMux I__10135 (
            .O(N__44502),
            .I(N__44477));
    InMux I__10134 (
            .O(N__44501),
            .I(N__44477));
    InMux I__10133 (
            .O(N__44500),
            .I(N__44477));
    InMux I__10132 (
            .O(N__44499),
            .I(N__44477));
    InMux I__10131 (
            .O(N__44498),
            .I(N__44474));
    InMux I__10130 (
            .O(N__44495),
            .I(N__44464));
    InMux I__10129 (
            .O(N__44494),
            .I(N__44464));
    InMux I__10128 (
            .O(N__44493),
            .I(N__44464));
    InMux I__10127 (
            .O(N__44492),
            .I(N__44464));
    InMux I__10126 (
            .O(N__44491),
            .I(N__44455));
    InMux I__10125 (
            .O(N__44490),
            .I(N__44455));
    InMux I__10124 (
            .O(N__44489),
            .I(N__44455));
    InMux I__10123 (
            .O(N__44488),
            .I(N__44455));
    LocalMux I__10122 (
            .O(N__44477),
            .I(N__44452));
    LocalMux I__10121 (
            .O(N__44474),
            .I(N__44449));
    InMux I__10120 (
            .O(N__44473),
            .I(N__44446));
    LocalMux I__10119 (
            .O(N__44464),
            .I(N__44443));
    LocalMux I__10118 (
            .O(N__44455),
            .I(N__44440));
    Span4Mux_v I__10117 (
            .O(N__44452),
            .I(N__44437));
    Span12Mux_v I__10116 (
            .O(N__44449),
            .I(N__44434));
    LocalMux I__10115 (
            .O(N__44446),
            .I(N__44427));
    Span12Mux_s8_h I__10114 (
            .O(N__44443),
            .I(N__44427));
    Span12Mux_v I__10113 (
            .O(N__44440),
            .I(N__44427));
    Odrv4 I__10112 (
            .O(N__44437),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv12 I__10111 (
            .O(N__44434),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    Odrv12 I__10110 (
            .O(N__44427),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ));
    InMux I__10109 (
            .O(N__44420),
            .I(N__44417));
    LocalMux I__10108 (
            .O(N__44417),
            .I(N__44414));
    Odrv4 I__10107 (
            .O(N__44414),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ));
    CEMux I__10106 (
            .O(N__44411),
            .I(N__44405));
    CEMux I__10105 (
            .O(N__44410),
            .I(N__44401));
    CEMux I__10104 (
            .O(N__44409),
            .I(N__44398));
    CEMux I__10103 (
            .O(N__44408),
            .I(N__44395));
    LocalMux I__10102 (
            .O(N__44405),
            .I(N__44392));
    CEMux I__10101 (
            .O(N__44404),
            .I(N__44389));
    LocalMux I__10100 (
            .O(N__44401),
            .I(N__44386));
    LocalMux I__10099 (
            .O(N__44398),
            .I(N__44383));
    LocalMux I__10098 (
            .O(N__44395),
            .I(N__44378));
    Span4Mux_v I__10097 (
            .O(N__44392),
            .I(N__44378));
    LocalMux I__10096 (
            .O(N__44389),
            .I(N__44375));
    Span4Mux_h I__10095 (
            .O(N__44386),
            .I(N__44372));
    Span4Mux_h I__10094 (
            .O(N__44383),
            .I(N__44369));
    Span4Mux_v I__10093 (
            .O(N__44378),
            .I(N__44366));
    Odrv12 I__10092 (
            .O(N__44375),
            .I(\ppm_encoder_1.N_1818_0 ));
    Odrv4 I__10091 (
            .O(N__44372),
            .I(\ppm_encoder_1.N_1818_0 ));
    Odrv4 I__10090 (
            .O(N__44369),
            .I(\ppm_encoder_1.N_1818_0 ));
    Odrv4 I__10089 (
            .O(N__44366),
            .I(\ppm_encoder_1.N_1818_0 ));
    InMux I__10088 (
            .O(N__44357),
            .I(N__44354));
    LocalMux I__10087 (
            .O(N__44354),
            .I(N__44351));
    Odrv4 I__10086 (
            .O(N__44351),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ));
    InMux I__10085 (
            .O(N__44348),
            .I(N__44345));
    LocalMux I__10084 (
            .O(N__44345),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ));
    InMux I__10083 (
            .O(N__44342),
            .I(N__44339));
    LocalMux I__10082 (
            .O(N__44339),
            .I(N__44336));
    Span4Mux_h I__10081 (
            .O(N__44336),
            .I(N__44333));
    Span4Mux_h I__10080 (
            .O(N__44333),
            .I(N__44330));
    Odrv4 I__10079 (
            .O(N__44330),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ));
    InMux I__10078 (
            .O(N__44327),
            .I(N__44324));
    LocalMux I__10077 (
            .O(N__44324),
            .I(N__44321));
    Span4Mux_h I__10076 (
            .O(N__44321),
            .I(N__44318));
    Odrv4 I__10075 (
            .O(N__44318),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ));
    InMux I__10074 (
            .O(N__44315),
            .I(N__44312));
    LocalMux I__10073 (
            .O(N__44312),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ));
    InMux I__10072 (
            .O(N__44309),
            .I(N__44306));
    LocalMux I__10071 (
            .O(N__44306),
            .I(N__44303));
    Odrv12 I__10070 (
            .O(N__44303),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ));
    InMux I__10069 (
            .O(N__44300),
            .I(N__44297));
    LocalMux I__10068 (
            .O(N__44297),
            .I(N__44294));
    Span4Mux_h I__10067 (
            .O(N__44294),
            .I(N__44291));
    Odrv4 I__10066 (
            .O(N__44291),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ));
    InMux I__10065 (
            .O(N__44288),
            .I(N__44285));
    LocalMux I__10064 (
            .O(N__44285),
            .I(N__44282));
    Span12Mux_v I__10063 (
            .O(N__44282),
            .I(N__44279));
    Odrv12 I__10062 (
            .O(N__44279),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ));
    InMux I__10061 (
            .O(N__44276),
            .I(N__44273));
    LocalMux I__10060 (
            .O(N__44273),
            .I(N__44270));
    Span4Mux_h I__10059 (
            .O(N__44270),
            .I(N__44267));
    Span4Mux_h I__10058 (
            .O(N__44267),
            .I(N__44264));
    Odrv4 I__10057 (
            .O(N__44264),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ));
    InMux I__10056 (
            .O(N__44261),
            .I(N__44255));
    InMux I__10055 (
            .O(N__44260),
            .I(N__44255));
    LocalMux I__10054 (
            .O(N__44255),
            .I(\ppm_encoder_1.pulses2countZ0Z_16 ));
    InMux I__10053 (
            .O(N__44252),
            .I(N__44249));
    LocalMux I__10052 (
            .O(N__44249),
            .I(N__44246));
    Span4Mux_h I__10051 (
            .O(N__44246),
            .I(N__44241));
    InMux I__10050 (
            .O(N__44245),
            .I(N__44236));
    InMux I__10049 (
            .O(N__44244),
            .I(N__44236));
    Odrv4 I__10048 (
            .O(N__44241),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    LocalMux I__10047 (
            .O(N__44236),
            .I(\ppm_encoder_1.init_pulsesZ0Z_17 ));
    CascadeMux I__10046 (
            .O(N__44231),
            .I(N__44227));
    CascadeMux I__10045 (
            .O(N__44230),
            .I(N__44224));
    InMux I__10044 (
            .O(N__44227),
            .I(N__44219));
    InMux I__10043 (
            .O(N__44224),
            .I(N__44219));
    LocalMux I__10042 (
            .O(N__44219),
            .I(\ppm_encoder_1.pulses2countZ0Z_17 ));
    InMux I__10041 (
            .O(N__44216),
            .I(N__44212));
    InMux I__10040 (
            .O(N__44215),
            .I(N__44209));
    LocalMux I__10039 (
            .O(N__44212),
            .I(N__44206));
    LocalMux I__10038 (
            .O(N__44209),
            .I(N__44203));
    Span4Mux_v I__10037 (
            .O(N__44206),
            .I(N__44197));
    Span4Mux_v I__10036 (
            .O(N__44203),
            .I(N__44197));
    InMux I__10035 (
            .O(N__44202),
            .I(N__44194));
    Odrv4 I__10034 (
            .O(N__44197),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    LocalMux I__10033 (
            .O(N__44194),
            .I(\ppm_encoder_1.init_pulsesZ0Z_15 ));
    InMux I__10032 (
            .O(N__44189),
            .I(N__44185));
    InMux I__10031 (
            .O(N__44188),
            .I(N__44182));
    LocalMux I__10030 (
            .O(N__44185),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    LocalMux I__10029 (
            .O(N__44182),
            .I(\ppm_encoder_1.pulses2countZ0Z_15 ));
    InMux I__10028 (
            .O(N__44177),
            .I(N__44174));
    LocalMux I__10027 (
            .O(N__44174),
            .I(N__44171));
    Span4Mux_v I__10026 (
            .O(N__44171),
            .I(N__44167));
    InMux I__10025 (
            .O(N__44170),
            .I(N__44164));
    Span4Mux_v I__10024 (
            .O(N__44167),
            .I(N__44158));
    LocalMux I__10023 (
            .O(N__44164),
            .I(N__44158));
    InMux I__10022 (
            .O(N__44163),
            .I(N__44155));
    Odrv4 I__10021 (
            .O(N__44158),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    LocalMux I__10020 (
            .O(N__44155),
            .I(\ppm_encoder_1.init_pulsesZ0Z_9 ));
    InMux I__10019 (
            .O(N__44150),
            .I(N__44147));
    LocalMux I__10018 (
            .O(N__44147),
            .I(N__44143));
    InMux I__10017 (
            .O(N__44146),
            .I(N__44140));
    Span4Mux_v I__10016 (
            .O(N__44143),
            .I(N__44135));
    LocalMux I__10015 (
            .O(N__44140),
            .I(N__44135));
    Span4Mux_v I__10014 (
            .O(N__44135),
            .I(N__44132));
    Span4Mux_h I__10013 (
            .O(N__44132),
            .I(N__44129));
    Odrv4 I__10012 (
            .O(N__44129),
            .I(\ppm_encoder_1.un1_init_pulses_0_9 ));
    InMux I__10011 (
            .O(N__44126),
            .I(N__44123));
    LocalMux I__10010 (
            .O(N__44123),
            .I(N__44119));
    InMux I__10009 (
            .O(N__44122),
            .I(N__44116));
    Span4Mux_v I__10008 (
            .O(N__44119),
            .I(N__44111));
    LocalMux I__10007 (
            .O(N__44116),
            .I(N__44111));
    Span4Mux_v I__10006 (
            .O(N__44111),
            .I(N__44108));
    Odrv4 I__10005 (
            .O(N__44108),
            .I(\ppm_encoder_1.un1_init_pulses_0_5 ));
    InMux I__10004 (
            .O(N__44105),
            .I(N__44102));
    LocalMux I__10003 (
            .O(N__44102),
            .I(N__44097));
    InMux I__10002 (
            .O(N__44101),
            .I(N__44094));
    InMux I__10001 (
            .O(N__44100),
            .I(N__44091));
    Span4Mux_v I__10000 (
            .O(N__44097),
            .I(N__44088));
    LocalMux I__9999 (
            .O(N__44094),
            .I(N__44083));
    LocalMux I__9998 (
            .O(N__44091),
            .I(N__44083));
    Odrv4 I__9997 (
            .O(N__44088),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    Odrv12 I__9996 (
            .O(N__44083),
            .I(\ppm_encoder_1.init_pulsesZ0Z_8 ));
    InMux I__9995 (
            .O(N__44078),
            .I(N__44074));
    InMux I__9994 (
            .O(N__44077),
            .I(N__44071));
    LocalMux I__9993 (
            .O(N__44074),
            .I(N__44068));
    LocalMux I__9992 (
            .O(N__44071),
            .I(N__44065));
    Span4Mux_v I__9991 (
            .O(N__44068),
            .I(N__44062));
    Span4Mux_h I__9990 (
            .O(N__44065),
            .I(N__44059));
    Odrv4 I__9989 (
            .O(N__44062),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    Odrv4 I__9988 (
            .O(N__44059),
            .I(\ppm_encoder_1.un1_init_pulses_0_8 ));
    InMux I__9987 (
            .O(N__44054),
            .I(N__44051));
    LocalMux I__9986 (
            .O(N__44051),
            .I(N__44048));
    Span4Mux_h I__9985 (
            .O(N__44048),
            .I(N__44045));
    Odrv4 I__9984 (
            .O(N__44045),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_15 ));
    InMux I__9983 (
            .O(N__44042),
            .I(N__44039));
    LocalMux I__9982 (
            .O(N__44039),
            .I(N__44035));
    CascadeMux I__9981 (
            .O(N__44038),
            .I(N__44031));
    Span4Mux_h I__9980 (
            .O(N__44035),
            .I(N__44028));
    InMux I__9979 (
            .O(N__44034),
            .I(N__44025));
    InMux I__9978 (
            .O(N__44031),
            .I(N__44022));
    Span4Mux_h I__9977 (
            .O(N__44028),
            .I(N__44017));
    LocalMux I__9976 (
            .O(N__44025),
            .I(N__44017));
    LocalMux I__9975 (
            .O(N__44022),
            .I(throttle_order_0));
    Odrv4 I__9974 (
            .O(N__44017),
            .I(throttle_order_0));
    InMux I__9973 (
            .O(N__44012),
            .I(N__44007));
    InMux I__9972 (
            .O(N__44011),
            .I(N__44004));
    InMux I__9971 (
            .O(N__44010),
            .I(N__44000));
    LocalMux I__9970 (
            .O(N__44007),
            .I(N__43995));
    LocalMux I__9969 (
            .O(N__44004),
            .I(N__43995));
    InMux I__9968 (
            .O(N__44003),
            .I(N__43992));
    LocalMux I__9967 (
            .O(N__44000),
            .I(N__43987));
    Span4Mux_v I__9966 (
            .O(N__43995),
            .I(N__43987));
    LocalMux I__9965 (
            .O(N__43992),
            .I(N__43982));
    Span4Mux_h I__9964 (
            .O(N__43987),
            .I(N__43982));
    Odrv4 I__9963 (
            .O(N__43982),
            .I(\ppm_encoder_1.elevatorZ0Z_0 ));
    InMux I__9962 (
            .O(N__43979),
            .I(N__43974));
    InMux I__9961 (
            .O(N__43978),
            .I(N__43969));
    InMux I__9960 (
            .O(N__43977),
            .I(N__43969));
    LocalMux I__9959 (
            .O(N__43974),
            .I(N__43966));
    LocalMux I__9958 (
            .O(N__43969),
            .I(N__43961));
    Span4Mux_v I__9957 (
            .O(N__43966),
            .I(N__43961));
    Odrv4 I__9956 (
            .O(N__43961),
            .I(\ppm_encoder_1.throttleZ0Z_0 ));
    InMux I__9955 (
            .O(N__43958),
            .I(N__43955));
    LocalMux I__9954 (
            .O(N__43955),
            .I(N__43950));
    InMux I__9953 (
            .O(N__43954),
            .I(N__43947));
    InMux I__9952 (
            .O(N__43953),
            .I(N__43941));
    Span4Mux_h I__9951 (
            .O(N__43950),
            .I(N__43936));
    LocalMux I__9950 (
            .O(N__43947),
            .I(N__43936));
    InMux I__9949 (
            .O(N__43946),
            .I(N__43929));
    InMux I__9948 (
            .O(N__43945),
            .I(N__43929));
    InMux I__9947 (
            .O(N__43944),
            .I(N__43929));
    LocalMux I__9946 (
            .O(N__43941),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    Odrv4 I__9945 (
            .O(N__43936),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    LocalMux I__9944 (
            .O(N__43929),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ));
    CascadeMux I__9943 (
            .O(N__43922),
            .I(\ppm_encoder_1.N_286_cascade_ ));
    InMux I__9942 (
            .O(N__43919),
            .I(N__43916));
    LocalMux I__9941 (
            .O(N__43916),
            .I(N__43913));
    Span4Mux_h I__9940 (
            .O(N__43913),
            .I(N__43910));
    Span4Mux_v I__9939 (
            .O(N__43910),
            .I(N__43907));
    Odrv4 I__9938 (
            .O(N__43907),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ));
    InMux I__9937 (
            .O(N__43904),
            .I(N__43899));
    InMux I__9936 (
            .O(N__43903),
            .I(N__43896));
    InMux I__9935 (
            .O(N__43902),
            .I(N__43893));
    LocalMux I__9934 (
            .O(N__43899),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    LocalMux I__9933 (
            .O(N__43896),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    LocalMux I__9932 (
            .O(N__43893),
            .I(\ppm_encoder_1.init_pulsesZ0Z_5 ));
    CascadeMux I__9931 (
            .O(N__43886),
            .I(N__43883));
    InMux I__9930 (
            .O(N__43883),
            .I(N__43875));
    InMux I__9929 (
            .O(N__43882),
            .I(N__43875));
    InMux I__9928 (
            .O(N__43881),
            .I(N__43872));
    InMux I__9927 (
            .O(N__43880),
            .I(N__43866));
    LocalMux I__9926 (
            .O(N__43875),
            .I(N__43861));
    LocalMux I__9925 (
            .O(N__43872),
            .I(N__43861));
    InMux I__9924 (
            .O(N__43871),
            .I(N__43856));
    InMux I__9923 (
            .O(N__43870),
            .I(N__43856));
    InMux I__9922 (
            .O(N__43869),
            .I(N__43853));
    LocalMux I__9921 (
            .O(N__43866),
            .I(N__43849));
    Span4Mux_v I__9920 (
            .O(N__43861),
            .I(N__43844));
    LocalMux I__9919 (
            .O(N__43856),
            .I(N__43844));
    LocalMux I__9918 (
            .O(N__43853),
            .I(N__43841));
    CascadeMux I__9917 (
            .O(N__43852),
            .I(N__43836));
    Span12Mux_v I__9916 (
            .O(N__43849),
            .I(N__43828));
    Span4Mux_v I__9915 (
            .O(N__43844),
            .I(N__43825));
    Span4Mux_h I__9914 (
            .O(N__43841),
            .I(N__43822));
    InMux I__9913 (
            .O(N__43840),
            .I(N__43819));
    InMux I__9912 (
            .O(N__43839),
            .I(N__43816));
    InMux I__9911 (
            .O(N__43836),
            .I(N__43811));
    InMux I__9910 (
            .O(N__43835),
            .I(N__43811));
    InMux I__9909 (
            .O(N__43834),
            .I(N__43806));
    InMux I__9908 (
            .O(N__43833),
            .I(N__43806));
    InMux I__9907 (
            .O(N__43832),
            .I(N__43801));
    InMux I__9906 (
            .O(N__43831),
            .I(N__43801));
    Odrv12 I__9905 (
            .O(N__43828),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9904 (
            .O(N__43825),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    Odrv4 I__9903 (
            .O(N__43822),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9902 (
            .O(N__43819),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9901 (
            .O(N__43816),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9900 (
            .O(N__43811),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9899 (
            .O(N__43806),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    LocalMux I__9898 (
            .O(N__43801),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_7 ));
    CascadeMux I__9897 (
            .O(N__43784),
            .I(N__43779));
    CascadeMux I__9896 (
            .O(N__43783),
            .I(N__43773));
    InMux I__9895 (
            .O(N__43782),
            .I(N__43767));
    InMux I__9894 (
            .O(N__43779),
            .I(N__43767));
    CascadeMux I__9893 (
            .O(N__43778),
            .I(N__43763));
    CascadeMux I__9892 (
            .O(N__43777),
            .I(N__43758));
    CascadeMux I__9891 (
            .O(N__43776),
            .I(N__43754));
    InMux I__9890 (
            .O(N__43773),
            .I(N__43750));
    CascadeMux I__9889 (
            .O(N__43772),
            .I(N__43746));
    LocalMux I__9888 (
            .O(N__43767),
            .I(N__43743));
    InMux I__9887 (
            .O(N__43766),
            .I(N__43740));
    InMux I__9886 (
            .O(N__43763),
            .I(N__43736));
    InMux I__9885 (
            .O(N__43762),
            .I(N__43729));
    InMux I__9884 (
            .O(N__43761),
            .I(N__43729));
    InMux I__9883 (
            .O(N__43758),
            .I(N__43729));
    InMux I__9882 (
            .O(N__43757),
            .I(N__43723));
    InMux I__9881 (
            .O(N__43754),
            .I(N__43723));
    InMux I__9880 (
            .O(N__43753),
            .I(N__43720));
    LocalMux I__9879 (
            .O(N__43750),
            .I(N__43717));
    InMux I__9878 (
            .O(N__43749),
            .I(N__43712));
    InMux I__9877 (
            .O(N__43746),
            .I(N__43712));
    Span4Mux_v I__9876 (
            .O(N__43743),
            .I(N__43705));
    LocalMux I__9875 (
            .O(N__43740),
            .I(N__43705));
    CascadeMux I__9874 (
            .O(N__43739),
            .I(N__43702));
    LocalMux I__9873 (
            .O(N__43736),
            .I(N__43696));
    LocalMux I__9872 (
            .O(N__43729),
            .I(N__43696));
    InMux I__9871 (
            .O(N__43728),
            .I(N__43693));
    LocalMux I__9870 (
            .O(N__43723),
            .I(N__43688));
    LocalMux I__9869 (
            .O(N__43720),
            .I(N__43688));
    Span4Mux_v I__9868 (
            .O(N__43717),
            .I(N__43683));
    LocalMux I__9867 (
            .O(N__43712),
            .I(N__43683));
    InMux I__9866 (
            .O(N__43711),
            .I(N__43678));
    InMux I__9865 (
            .O(N__43710),
            .I(N__43678));
    Span4Mux_v I__9864 (
            .O(N__43705),
            .I(N__43675));
    InMux I__9863 (
            .O(N__43702),
            .I(N__43672));
    InMux I__9862 (
            .O(N__43701),
            .I(N__43669));
    Span4Mux_h I__9861 (
            .O(N__43696),
            .I(N__43662));
    LocalMux I__9860 (
            .O(N__43693),
            .I(N__43662));
    Span4Mux_v I__9859 (
            .O(N__43688),
            .I(N__43662));
    Span4Mux_v I__9858 (
            .O(N__43683),
            .I(N__43655));
    LocalMux I__9857 (
            .O(N__43678),
            .I(N__43655));
    Span4Mux_h I__9856 (
            .O(N__43675),
            .I(N__43655));
    LocalMux I__9855 (
            .O(N__43672),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    LocalMux I__9854 (
            .O(N__43669),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9853 (
            .O(N__43662),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    Odrv4 I__9852 (
            .O(N__43655),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ));
    InMux I__9851 (
            .O(N__43646),
            .I(N__43643));
    LocalMux I__9850 (
            .O(N__43643),
            .I(N__43639));
    InMux I__9849 (
            .O(N__43642),
            .I(N__43636));
    Span4Mux_v I__9848 (
            .O(N__43639),
            .I(N__43633));
    LocalMux I__9847 (
            .O(N__43636),
            .I(N__43630));
    Odrv4 I__9846 (
            .O(N__43633),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    Odrv12 I__9845 (
            .O(N__43630),
            .I(\ppm_encoder_1.rudderZ0Z_5 ));
    InMux I__9844 (
            .O(N__43625),
            .I(N__43622));
    LocalMux I__9843 (
            .O(N__43622),
            .I(drone_H_disp_front_i_9));
    CascadeMux I__9842 (
            .O(N__43619),
            .I(N__43616));
    InMux I__9841 (
            .O(N__43616),
            .I(N__43613));
    LocalMux I__9840 (
            .O(N__43613),
            .I(front_command_5));
    InMux I__9839 (
            .O(N__43610),
            .I(N__43607));
    LocalMux I__9838 (
            .O(N__43607),
            .I(N__43604));
    Span12Mux_s8_h I__9837 (
            .O(N__43604),
            .I(N__43601));
    Odrv12 I__9836 (
            .O(N__43601),
            .I(\pid_front.error_9 ));
    InMux I__9835 (
            .O(N__43598),
            .I(\pid_front.error_cry_4 ));
    InMux I__9834 (
            .O(N__43595),
            .I(N__43592));
    LocalMux I__9833 (
            .O(N__43592),
            .I(N__43589));
    Odrv4 I__9832 (
            .O(N__43589),
            .I(front_command_6));
    CascadeMux I__9831 (
            .O(N__43586),
            .I(N__43583));
    InMux I__9830 (
            .O(N__43583),
            .I(N__43580));
    LocalMux I__9829 (
            .O(N__43580),
            .I(drone_H_disp_front_i_10));
    InMux I__9828 (
            .O(N__43577),
            .I(N__43574));
    LocalMux I__9827 (
            .O(N__43574),
            .I(N__43571));
    Span4Mux_s3_h I__9826 (
            .O(N__43571),
            .I(N__43568));
    Span4Mux_h I__9825 (
            .O(N__43568),
            .I(N__43565));
    Odrv4 I__9824 (
            .O(N__43565),
            .I(\pid_front.error_10 ));
    InMux I__9823 (
            .O(N__43562),
            .I(\pid_front.error_cry_5 ));
    InMux I__9822 (
            .O(N__43559),
            .I(N__43556));
    LocalMux I__9821 (
            .O(N__43556),
            .I(\pid_front.error_axbZ0Z_7 ));
    InMux I__9820 (
            .O(N__43553),
            .I(N__43550));
    LocalMux I__9819 (
            .O(N__43550),
            .I(N__43547));
    Span4Mux_v I__9818 (
            .O(N__43547),
            .I(N__43544));
    Span4Mux_h I__9817 (
            .O(N__43544),
            .I(N__43541));
    Odrv4 I__9816 (
            .O(N__43541),
            .I(\pid_front.error_11 ));
    InMux I__9815 (
            .O(N__43538),
            .I(\pid_front.error_cry_6 ));
    InMux I__9814 (
            .O(N__43535),
            .I(N__43532));
    LocalMux I__9813 (
            .O(N__43532),
            .I(\pid_front.error_axb_8_l_ofx_0 ));
    CascadeMux I__9812 (
            .O(N__43529),
            .I(N__43526));
    InMux I__9811 (
            .O(N__43526),
            .I(N__43522));
    InMux I__9810 (
            .O(N__43525),
            .I(N__43519));
    LocalMux I__9809 (
            .O(N__43522),
            .I(N__43515));
    LocalMux I__9808 (
            .O(N__43519),
            .I(N__43512));
    InMux I__9807 (
            .O(N__43518),
            .I(N__43509));
    Span4Mux_h I__9806 (
            .O(N__43515),
            .I(N__43504));
    Span4Mux_h I__9805 (
            .O(N__43512),
            .I(N__43504));
    LocalMux I__9804 (
            .O(N__43509),
            .I(drone_H_disp_front_12));
    Odrv4 I__9803 (
            .O(N__43504),
            .I(drone_H_disp_front_12));
    InMux I__9802 (
            .O(N__43499),
            .I(N__43496));
    LocalMux I__9801 (
            .O(N__43496),
            .I(N__43493));
    Span4Mux_v I__9800 (
            .O(N__43493),
            .I(N__43490));
    Span4Mux_h I__9799 (
            .O(N__43490),
            .I(N__43487));
    Odrv4 I__9798 (
            .O(N__43487),
            .I(\pid_front.error_12 ));
    InMux I__9797 (
            .O(N__43484),
            .I(\pid_front.error_cry_7 ));
    InMux I__9796 (
            .O(N__43481),
            .I(N__43478));
    LocalMux I__9795 (
            .O(N__43478),
            .I(N__43475));
    Odrv12 I__9794 (
            .O(N__43475),
            .I(drone_H_disp_front_i_12));
    CascadeMux I__9793 (
            .O(N__43472),
            .I(N__43469));
    InMux I__9792 (
            .O(N__43469),
            .I(N__43465));
    InMux I__9791 (
            .O(N__43468),
            .I(N__43462));
    LocalMux I__9790 (
            .O(N__43465),
            .I(N__43459));
    LocalMux I__9789 (
            .O(N__43462),
            .I(N__43456));
    Odrv4 I__9788 (
            .O(N__43459),
            .I(drone_H_disp_front_13));
    Odrv4 I__9787 (
            .O(N__43456),
            .I(drone_H_disp_front_13));
    InMux I__9786 (
            .O(N__43451),
            .I(N__43448));
    LocalMux I__9785 (
            .O(N__43448),
            .I(N__43445));
    Span4Mux_v I__9784 (
            .O(N__43445),
            .I(N__43442));
    Span4Mux_h I__9783 (
            .O(N__43442),
            .I(N__43439));
    Odrv4 I__9782 (
            .O(N__43439),
            .I(\pid_front.error_13 ));
    InMux I__9781 (
            .O(N__43436),
            .I(\pid_front.error_cry_8 ));
    InMux I__9780 (
            .O(N__43433),
            .I(N__43430));
    LocalMux I__9779 (
            .O(N__43430),
            .I(N__43427));
    Odrv4 I__9778 (
            .O(N__43427),
            .I(drone_H_disp_front_i_13));
    InMux I__9777 (
            .O(N__43424),
            .I(N__43421));
    LocalMux I__9776 (
            .O(N__43421),
            .I(N__43418));
    Span4Mux_s3_h I__9775 (
            .O(N__43418),
            .I(N__43415));
    Span4Mux_h I__9774 (
            .O(N__43415),
            .I(N__43412));
    Odrv4 I__9773 (
            .O(N__43412),
            .I(\pid_front.error_14 ));
    InMux I__9772 (
            .O(N__43409),
            .I(\pid_front.error_cry_9 ));
    InMux I__9771 (
            .O(N__43406),
            .I(N__43403));
    LocalMux I__9770 (
            .O(N__43403),
            .I(N__43400));
    Span4Mux_h I__9769 (
            .O(N__43400),
            .I(N__43397));
    Odrv4 I__9768 (
            .O(N__43397),
            .I(drone_H_disp_front_15));
    InMux I__9767 (
            .O(N__43394),
            .I(\pid_front.error_cry_10 ));
    InMux I__9766 (
            .O(N__43391),
            .I(N__43388));
    LocalMux I__9765 (
            .O(N__43388),
            .I(N__43385));
    Span4Mux_s3_h I__9764 (
            .O(N__43385),
            .I(N__43382));
    Span4Mux_h I__9763 (
            .O(N__43382),
            .I(N__43379));
    Odrv4 I__9762 (
            .O(N__43379),
            .I(\pid_front.error_15 ));
    InMux I__9761 (
            .O(N__43376),
            .I(N__43367));
    InMux I__9760 (
            .O(N__43375),
            .I(N__43367));
    CascadeMux I__9759 (
            .O(N__43374),
            .I(N__43363));
    CascadeMux I__9758 (
            .O(N__43373),
            .I(N__43355));
    InMux I__9757 (
            .O(N__43372),
            .I(N__43347));
    LocalMux I__9756 (
            .O(N__43367),
            .I(N__43344));
    InMux I__9755 (
            .O(N__43366),
            .I(N__43341));
    InMux I__9754 (
            .O(N__43363),
            .I(N__43338));
    InMux I__9753 (
            .O(N__43362),
            .I(N__43331));
    InMux I__9752 (
            .O(N__43361),
            .I(N__43331));
    InMux I__9751 (
            .O(N__43360),
            .I(N__43331));
    InMux I__9750 (
            .O(N__43359),
            .I(N__43326));
    InMux I__9749 (
            .O(N__43358),
            .I(N__43326));
    InMux I__9748 (
            .O(N__43355),
            .I(N__43323));
    InMux I__9747 (
            .O(N__43354),
            .I(N__43318));
    InMux I__9746 (
            .O(N__43353),
            .I(N__43318));
    InMux I__9745 (
            .O(N__43352),
            .I(N__43311));
    InMux I__9744 (
            .O(N__43351),
            .I(N__43311));
    InMux I__9743 (
            .O(N__43350),
            .I(N__43311));
    LocalMux I__9742 (
            .O(N__43347),
            .I(N__43305));
    Span4Mux_v I__9741 (
            .O(N__43344),
            .I(N__43300));
    LocalMux I__9740 (
            .O(N__43341),
            .I(N__43300));
    LocalMux I__9739 (
            .O(N__43338),
            .I(N__43287));
    LocalMux I__9738 (
            .O(N__43331),
            .I(N__43287));
    LocalMux I__9737 (
            .O(N__43326),
            .I(N__43287));
    LocalMux I__9736 (
            .O(N__43323),
            .I(N__43287));
    LocalMux I__9735 (
            .O(N__43318),
            .I(N__43287));
    LocalMux I__9734 (
            .O(N__43311),
            .I(N__43287));
    InMux I__9733 (
            .O(N__43310),
            .I(N__43280));
    InMux I__9732 (
            .O(N__43309),
            .I(N__43280));
    InMux I__9731 (
            .O(N__43308),
            .I(N__43280));
    Span4Mux_v I__9730 (
            .O(N__43305),
            .I(N__43275));
    Span4Mux_h I__9729 (
            .O(N__43300),
            .I(N__43275));
    Span4Mux_v I__9728 (
            .O(N__43287),
            .I(N__43272));
    LocalMux I__9727 (
            .O(N__43280),
            .I(N__43269));
    Span4Mux_v I__9726 (
            .O(N__43275),
            .I(N__43266));
    Span4Mux_v I__9725 (
            .O(N__43272),
            .I(N__43263));
    Odrv12 I__9724 (
            .O(N__43269),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__9723 (
            .O(N__43266),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    Odrv4 I__9722 (
            .O(N__43263),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ));
    InMux I__9721 (
            .O(N__43256),
            .I(N__43253));
    LocalMux I__9720 (
            .O(N__43253),
            .I(N__43250));
    Span4Mux_h I__9719 (
            .O(N__43250),
            .I(N__43247));
    Odrv4 I__9718 (
            .O(N__43247),
            .I(\ppm_encoder_1.un1_init_pulses_11_9 ));
    CascadeMux I__9717 (
            .O(N__43244),
            .I(N__43233));
    CascadeMux I__9716 (
            .O(N__43243),
            .I(N__43230));
    CascadeMux I__9715 (
            .O(N__43242),
            .I(N__43227));
    CascadeMux I__9714 (
            .O(N__43241),
            .I(N__43224));
    CascadeMux I__9713 (
            .O(N__43240),
            .I(N__43215));
    CascadeMux I__9712 (
            .O(N__43239),
            .I(N__43212));
    CascadeMux I__9711 (
            .O(N__43238),
            .I(N__43209));
    InMux I__9710 (
            .O(N__43237),
            .I(N__43204));
    InMux I__9709 (
            .O(N__43236),
            .I(N__43204));
    InMux I__9708 (
            .O(N__43233),
            .I(N__43201));
    InMux I__9707 (
            .O(N__43230),
            .I(N__43196));
    InMux I__9706 (
            .O(N__43227),
            .I(N__43196));
    InMux I__9705 (
            .O(N__43224),
            .I(N__43193));
    InMux I__9704 (
            .O(N__43223),
            .I(N__43190));
    InMux I__9703 (
            .O(N__43222),
            .I(N__43185));
    InMux I__9702 (
            .O(N__43221),
            .I(N__43185));
    CascadeMux I__9701 (
            .O(N__43220),
            .I(N__43182));
    CascadeMux I__9700 (
            .O(N__43219),
            .I(N__43179));
    CascadeMux I__9699 (
            .O(N__43218),
            .I(N__43172));
    InMux I__9698 (
            .O(N__43215),
            .I(N__43167));
    InMux I__9697 (
            .O(N__43212),
            .I(N__43167));
    InMux I__9696 (
            .O(N__43209),
            .I(N__43164));
    LocalMux I__9695 (
            .O(N__43204),
            .I(N__43161));
    LocalMux I__9694 (
            .O(N__43201),
            .I(N__43156));
    LocalMux I__9693 (
            .O(N__43196),
            .I(N__43156));
    LocalMux I__9692 (
            .O(N__43193),
            .I(N__43149));
    LocalMux I__9691 (
            .O(N__43190),
            .I(N__43149));
    LocalMux I__9690 (
            .O(N__43185),
            .I(N__43149));
    InMux I__9689 (
            .O(N__43182),
            .I(N__43146));
    InMux I__9688 (
            .O(N__43179),
            .I(N__43141));
    InMux I__9687 (
            .O(N__43178),
            .I(N__43141));
    InMux I__9686 (
            .O(N__43177),
            .I(N__43136));
    InMux I__9685 (
            .O(N__43176),
            .I(N__43136));
    InMux I__9684 (
            .O(N__43175),
            .I(N__43133));
    InMux I__9683 (
            .O(N__43172),
            .I(N__43130));
    LocalMux I__9682 (
            .O(N__43167),
            .I(N__43125));
    LocalMux I__9681 (
            .O(N__43164),
            .I(N__43125));
    Span4Mux_h I__9680 (
            .O(N__43161),
            .I(N__43122));
    Span4Mux_h I__9679 (
            .O(N__43156),
            .I(N__43117));
    Span4Mux_h I__9678 (
            .O(N__43149),
            .I(N__43117));
    LocalMux I__9677 (
            .O(N__43146),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9676 (
            .O(N__43141),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9675 (
            .O(N__43136),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9674 (
            .O(N__43133),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    LocalMux I__9673 (
            .O(N__43130),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv12 I__9672 (
            .O(N__43125),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__9671 (
            .O(N__43122),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    Odrv4 I__9670 (
            .O(N__43117),
            .I(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ));
    InMux I__9669 (
            .O(N__43100),
            .I(N__43097));
    LocalMux I__9668 (
            .O(N__43097),
            .I(N__43094));
    Span4Mux_h I__9667 (
            .O(N__43094),
            .I(N__43091));
    Odrv4 I__9666 (
            .O(N__43091),
            .I(\ppm_encoder_1.un1_init_pulses_10_9 ));
    InMux I__9665 (
            .O(N__43088),
            .I(N__43085));
    LocalMux I__9664 (
            .O(N__43085),
            .I(N__43082));
    Span12Mux_s9_v I__9663 (
            .O(N__43082),
            .I(N__43079));
    Odrv12 I__9662 (
            .O(N__43079),
            .I(\pid_front.error_axbZ0Z_2 ));
    InMux I__9661 (
            .O(N__43076),
            .I(N__43073));
    LocalMux I__9660 (
            .O(N__43073),
            .I(N__43070));
    Span12Mux_s8_h I__9659 (
            .O(N__43070),
            .I(N__43067));
    Odrv12 I__9658 (
            .O(N__43067),
            .I(\pid_front.error_2 ));
    InMux I__9657 (
            .O(N__43064),
            .I(\pid_front.error_cry_1 ));
    InMux I__9656 (
            .O(N__43061),
            .I(N__43058));
    LocalMux I__9655 (
            .O(N__43058),
            .I(N__43055));
    Span4Mux_h I__9654 (
            .O(N__43055),
            .I(N__43052));
    Span4Mux_h I__9653 (
            .O(N__43052),
            .I(N__43049));
    Odrv4 I__9652 (
            .O(N__43049),
            .I(\pid_front.error_axbZ0Z_3 ));
    InMux I__9651 (
            .O(N__43046),
            .I(N__43043));
    LocalMux I__9650 (
            .O(N__43043),
            .I(N__43040));
    Span4Mux_v I__9649 (
            .O(N__43040),
            .I(N__43037));
    Span4Mux_h I__9648 (
            .O(N__43037),
            .I(N__43034));
    Odrv4 I__9647 (
            .O(N__43034),
            .I(\pid_front.error_3 ));
    InMux I__9646 (
            .O(N__43031),
            .I(\pid_front.error_cry_2 ));
    InMux I__9645 (
            .O(N__43028),
            .I(N__43025));
    LocalMux I__9644 (
            .O(N__43025),
            .I(front_command_0));
    CascadeMux I__9643 (
            .O(N__43022),
            .I(N__43019));
    InMux I__9642 (
            .O(N__43019),
            .I(N__43016));
    LocalMux I__9641 (
            .O(N__43016),
            .I(drone_H_disp_front_i_4));
    InMux I__9640 (
            .O(N__43013),
            .I(N__43010));
    LocalMux I__9639 (
            .O(N__43010),
            .I(N__43007));
    Span4Mux_v I__9638 (
            .O(N__43007),
            .I(N__43004));
    Span4Mux_h I__9637 (
            .O(N__43004),
            .I(N__43001));
    Odrv4 I__9636 (
            .O(N__43001),
            .I(\pid_front.error_4 ));
    InMux I__9635 (
            .O(N__42998),
            .I(\pid_front.error_cry_3 ));
    InMux I__9634 (
            .O(N__42995),
            .I(N__42992));
    LocalMux I__9633 (
            .O(N__42992),
            .I(drone_H_disp_front_i_5));
    CascadeMux I__9632 (
            .O(N__42989),
            .I(N__42986));
    InMux I__9631 (
            .O(N__42986),
            .I(N__42983));
    LocalMux I__9630 (
            .O(N__42983),
            .I(front_command_1));
    InMux I__9629 (
            .O(N__42980),
            .I(N__42977));
    LocalMux I__9628 (
            .O(N__42977),
            .I(N__42974));
    Span4Mux_s3_h I__9627 (
            .O(N__42974),
            .I(N__42971));
    Span4Mux_h I__9626 (
            .O(N__42971),
            .I(N__42968));
    Odrv4 I__9625 (
            .O(N__42968),
            .I(\pid_front.error_5 ));
    InMux I__9624 (
            .O(N__42965),
            .I(\pid_front.error_cry_0_0 ));
    InMux I__9623 (
            .O(N__42962),
            .I(N__42959));
    LocalMux I__9622 (
            .O(N__42959),
            .I(drone_H_disp_front_i_6));
    CascadeMux I__9621 (
            .O(N__42956),
            .I(N__42953));
    InMux I__9620 (
            .O(N__42953),
            .I(N__42950));
    LocalMux I__9619 (
            .O(N__42950),
            .I(front_command_2));
    InMux I__9618 (
            .O(N__42947),
            .I(N__42944));
    LocalMux I__9617 (
            .O(N__42944),
            .I(N__42941));
    Span4Mux_s3_h I__9616 (
            .O(N__42941),
            .I(N__42938));
    Span4Mux_h I__9615 (
            .O(N__42938),
            .I(N__42935));
    Odrv4 I__9614 (
            .O(N__42935),
            .I(\pid_front.error_6 ));
    InMux I__9613 (
            .O(N__42932),
            .I(\pid_front.error_cry_1_0 ));
    InMux I__9612 (
            .O(N__42929),
            .I(N__42926));
    LocalMux I__9611 (
            .O(N__42926),
            .I(drone_H_disp_front_i_7));
    CascadeMux I__9610 (
            .O(N__42923),
            .I(N__42920));
    InMux I__9609 (
            .O(N__42920),
            .I(N__42917));
    LocalMux I__9608 (
            .O(N__42917),
            .I(front_command_3));
    InMux I__9607 (
            .O(N__42914),
            .I(N__42911));
    LocalMux I__9606 (
            .O(N__42911),
            .I(N__42908));
    Span4Mux_s3_h I__9605 (
            .O(N__42908),
            .I(N__42905));
    Span4Mux_h I__9604 (
            .O(N__42905),
            .I(N__42902));
    Odrv4 I__9603 (
            .O(N__42902),
            .I(\pid_front.error_7 ));
    InMux I__9602 (
            .O(N__42899),
            .I(\pid_front.error_cry_2_0 ));
    InMux I__9601 (
            .O(N__42896),
            .I(N__42893));
    LocalMux I__9600 (
            .O(N__42893),
            .I(front_command_4));
    CascadeMux I__9599 (
            .O(N__42890),
            .I(N__42887));
    InMux I__9598 (
            .O(N__42887),
            .I(N__42884));
    LocalMux I__9597 (
            .O(N__42884),
            .I(N__42881));
    Span4Mux_h I__9596 (
            .O(N__42881),
            .I(N__42878));
    Odrv4 I__9595 (
            .O(N__42878),
            .I(drone_H_disp_front_i_8));
    InMux I__9594 (
            .O(N__42875),
            .I(N__42872));
    LocalMux I__9593 (
            .O(N__42872),
            .I(N__42869));
    Span4Mux_s3_h I__9592 (
            .O(N__42869),
            .I(N__42866));
    Span4Mux_h I__9591 (
            .O(N__42866),
            .I(N__42863));
    Odrv4 I__9590 (
            .O(N__42863),
            .I(\pid_front.error_8 ));
    InMux I__9589 (
            .O(N__42860),
            .I(bfn_17_24_0_));
    CascadeMux I__9588 (
            .O(N__42857),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ));
    CascadeMux I__9587 (
            .O(N__42854),
            .I(N__42850));
    InMux I__9586 (
            .O(N__42853),
            .I(N__42847));
    InMux I__9585 (
            .O(N__42850),
            .I(N__42844));
    LocalMux I__9584 (
            .O(N__42847),
            .I(N__42839));
    LocalMux I__9583 (
            .O(N__42844),
            .I(N__42839));
    Odrv4 I__9582 (
            .O(N__42839),
            .I(\ppm_encoder_1.N_139_17 ));
    InMux I__9581 (
            .O(N__42836),
            .I(N__42833));
    LocalMux I__9580 (
            .O(N__42833),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ));
    InMux I__9579 (
            .O(N__42830),
            .I(N__42824));
    InMux I__9578 (
            .O(N__42829),
            .I(N__42824));
    LocalMux I__9577 (
            .O(N__42824),
            .I(N__42821));
    Odrv12 I__9576 (
            .O(N__42821),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ));
    CascadeMux I__9575 (
            .O(N__42818),
            .I(N__42811));
    CascadeMux I__9574 (
            .O(N__42817),
            .I(N__42806));
    CascadeMux I__9573 (
            .O(N__42816),
            .I(N__42795));
    CascadeMux I__9572 (
            .O(N__42815),
            .I(N__42792));
    InMux I__9571 (
            .O(N__42814),
            .I(N__42788));
    InMux I__9570 (
            .O(N__42811),
            .I(N__42785));
    InMux I__9569 (
            .O(N__42810),
            .I(N__42780));
    InMux I__9568 (
            .O(N__42809),
            .I(N__42780));
    InMux I__9567 (
            .O(N__42806),
            .I(N__42777));
    CascadeMux I__9566 (
            .O(N__42805),
            .I(N__42772));
    CascadeMux I__9565 (
            .O(N__42804),
            .I(N__42768));
    CascadeMux I__9564 (
            .O(N__42803),
            .I(N__42765));
    InMux I__9563 (
            .O(N__42802),
            .I(N__42761));
    InMux I__9562 (
            .O(N__42801),
            .I(N__42756));
    InMux I__9561 (
            .O(N__42800),
            .I(N__42756));
    InMux I__9560 (
            .O(N__42799),
            .I(N__42751));
    InMux I__9559 (
            .O(N__42798),
            .I(N__42751));
    InMux I__9558 (
            .O(N__42795),
            .I(N__42744));
    InMux I__9557 (
            .O(N__42792),
            .I(N__42744));
    InMux I__9556 (
            .O(N__42791),
            .I(N__42744));
    LocalMux I__9555 (
            .O(N__42788),
            .I(N__42737));
    LocalMux I__9554 (
            .O(N__42785),
            .I(N__42737));
    LocalMux I__9553 (
            .O(N__42780),
            .I(N__42737));
    LocalMux I__9552 (
            .O(N__42777),
            .I(N__42734));
    InMux I__9551 (
            .O(N__42776),
            .I(N__42727));
    InMux I__9550 (
            .O(N__42775),
            .I(N__42727));
    InMux I__9549 (
            .O(N__42772),
            .I(N__42727));
    CascadeMux I__9548 (
            .O(N__42771),
            .I(N__42723));
    InMux I__9547 (
            .O(N__42768),
            .I(N__42716));
    InMux I__9546 (
            .O(N__42765),
            .I(N__42716));
    InMux I__9545 (
            .O(N__42764),
            .I(N__42716));
    LocalMux I__9544 (
            .O(N__42761),
            .I(N__42713));
    LocalMux I__9543 (
            .O(N__42756),
            .I(N__42704));
    LocalMux I__9542 (
            .O(N__42751),
            .I(N__42704));
    LocalMux I__9541 (
            .O(N__42744),
            .I(N__42704));
    Span4Mux_v I__9540 (
            .O(N__42737),
            .I(N__42704));
    Span4Mux_v I__9539 (
            .O(N__42734),
            .I(N__42699));
    LocalMux I__9538 (
            .O(N__42727),
            .I(N__42699));
    InMux I__9537 (
            .O(N__42726),
            .I(N__42696));
    InMux I__9536 (
            .O(N__42723),
            .I(N__42691));
    LocalMux I__9535 (
            .O(N__42716),
            .I(N__42688));
    Span4Mux_h I__9534 (
            .O(N__42713),
            .I(N__42683));
    Span4Mux_h I__9533 (
            .O(N__42704),
            .I(N__42683));
    Sp12to4 I__9532 (
            .O(N__42699),
            .I(N__42678));
    LocalMux I__9531 (
            .O(N__42696),
            .I(N__42678));
    InMux I__9530 (
            .O(N__42695),
            .I(N__42675));
    InMux I__9529 (
            .O(N__42694),
            .I(N__42672));
    LocalMux I__9528 (
            .O(N__42691),
            .I(N__42662));
    Span12Mux_h I__9527 (
            .O(N__42688),
            .I(N__42662));
    Sp12to4 I__9526 (
            .O(N__42683),
            .I(N__42662));
    Span12Mux_h I__9525 (
            .O(N__42678),
            .I(N__42662));
    LocalMux I__9524 (
            .O(N__42675),
            .I(N__42657));
    LocalMux I__9523 (
            .O(N__42672),
            .I(N__42657));
    InMux I__9522 (
            .O(N__42671),
            .I(N__42654));
    Span12Mux_v I__9521 (
            .O(N__42662),
            .I(N__42651));
    Span4Mux_v I__9520 (
            .O(N__42657),
            .I(N__42648));
    LocalMux I__9519 (
            .O(N__42654),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv12 I__9518 (
            .O(N__42651),
            .I(\pid_front.stateZ0Z_0 ));
    Odrv4 I__9517 (
            .O(N__42648),
            .I(\pid_front.stateZ0Z_0 ));
    InMux I__9516 (
            .O(N__42641),
            .I(N__42634));
    InMux I__9515 (
            .O(N__42640),
            .I(N__42634));
    InMux I__9514 (
            .O(N__42639),
            .I(N__42631));
    LocalMux I__9513 (
            .O(N__42634),
            .I(N__42627));
    LocalMux I__9512 (
            .O(N__42631),
            .I(N__42624));
    InMux I__9511 (
            .O(N__42630),
            .I(N__42621));
    Span4Mux_h I__9510 (
            .O(N__42627),
            .I(N__42616));
    Span4Mux_h I__9509 (
            .O(N__42624),
            .I(N__42616));
    LocalMux I__9508 (
            .O(N__42621),
            .I(\pid_front.pid_preregZ0Z_8 ));
    Odrv4 I__9507 (
            .O(N__42616),
            .I(\pid_front.pid_preregZ0Z_8 ));
    InMux I__9506 (
            .O(N__42611),
            .I(N__42607));
    InMux I__9505 (
            .O(N__42610),
            .I(N__42602));
    LocalMux I__9504 (
            .O(N__42607),
            .I(N__42598));
    InMux I__9503 (
            .O(N__42606),
            .I(N__42595));
    InMux I__9502 (
            .O(N__42605),
            .I(N__42592));
    LocalMux I__9501 (
            .O(N__42602),
            .I(N__42589));
    InMux I__9500 (
            .O(N__42601),
            .I(N__42586));
    Span4Mux_h I__9499 (
            .O(N__42598),
            .I(N__42581));
    LocalMux I__9498 (
            .O(N__42595),
            .I(N__42581));
    LocalMux I__9497 (
            .O(N__42592),
            .I(N__42578));
    Span4Mux_v I__9496 (
            .O(N__42589),
            .I(N__42575));
    LocalMux I__9495 (
            .O(N__42586),
            .I(N__42572));
    Span4Mux_v I__9494 (
            .O(N__42581),
            .I(N__42567));
    Span4Mux_v I__9493 (
            .O(N__42578),
            .I(N__42564));
    Span4Mux_h I__9492 (
            .O(N__42575),
            .I(N__42559));
    Span4Mux_v I__9491 (
            .O(N__42572),
            .I(N__42559));
    InMux I__9490 (
            .O(N__42571),
            .I(N__42556));
    InMux I__9489 (
            .O(N__42570),
            .I(N__42553));
    Span4Mux_h I__9488 (
            .O(N__42567),
            .I(N__42548));
    Span4Mux_v I__9487 (
            .O(N__42564),
            .I(N__42548));
    Span4Mux_v I__9486 (
            .O(N__42559),
            .I(N__42543));
    LocalMux I__9485 (
            .O(N__42556),
            .I(N__42543));
    LocalMux I__9484 (
            .O(N__42553),
            .I(N__42540));
    Span4Mux_v I__9483 (
            .O(N__42548),
            .I(N__42535));
    Span4Mux_v I__9482 (
            .O(N__42543),
            .I(N__42535));
    Span4Mux_h I__9481 (
            .O(N__42540),
            .I(N__42532));
    Odrv4 I__9480 (
            .O(N__42535),
            .I(uart_drone_data_0));
    Odrv4 I__9479 (
            .O(N__42532),
            .I(uart_drone_data_0));
    CEMux I__9478 (
            .O(N__42527),
            .I(N__42523));
    CEMux I__9477 (
            .O(N__42526),
            .I(N__42520));
    LocalMux I__9476 (
            .O(N__42523),
            .I(N__42516));
    LocalMux I__9475 (
            .O(N__42520),
            .I(N__42513));
    CEMux I__9474 (
            .O(N__42519),
            .I(N__42510));
    Span4Mux_h I__9473 (
            .O(N__42516),
            .I(N__42506));
    Span4Mux_h I__9472 (
            .O(N__42513),
            .I(N__42501));
    LocalMux I__9471 (
            .O(N__42510),
            .I(N__42501));
    CEMux I__9470 (
            .O(N__42509),
            .I(N__42498));
    Span4Mux_h I__9469 (
            .O(N__42506),
            .I(N__42495));
    Span4Mux_h I__9468 (
            .O(N__42501),
            .I(N__42492));
    LocalMux I__9467 (
            .O(N__42498),
            .I(N__42489));
    Odrv4 I__9466 (
            .O(N__42495),
            .I(\dron_frame_decoder_1.N_731_0 ));
    Odrv4 I__9465 (
            .O(N__42492),
            .I(\dron_frame_decoder_1.N_731_0 ));
    Odrv4 I__9464 (
            .O(N__42489),
            .I(\dron_frame_decoder_1.N_731_0 ));
    InMux I__9463 (
            .O(N__42482),
            .I(N__42479));
    LocalMux I__9462 (
            .O(N__42479),
            .I(N__42476));
    Span4Mux_s3_h I__9461 (
            .O(N__42476),
            .I(N__42473));
    Span4Mux_h I__9460 (
            .O(N__42473),
            .I(N__42469));
    InMux I__9459 (
            .O(N__42472),
            .I(N__42466));
    Odrv4 I__9458 (
            .O(N__42469),
            .I(drone_H_disp_front_0));
    LocalMux I__9457 (
            .O(N__42466),
            .I(drone_H_disp_front_0));
    InMux I__9456 (
            .O(N__42461),
            .I(N__42458));
    LocalMux I__9455 (
            .O(N__42458),
            .I(\pid_front.error_axb_0 ));
    InMux I__9454 (
            .O(N__42455),
            .I(N__42452));
    LocalMux I__9453 (
            .O(N__42452),
            .I(N__42449));
    Span4Mux_v I__9452 (
            .O(N__42449),
            .I(N__42446));
    Odrv4 I__9451 (
            .O(N__42446),
            .I(\pid_front.error_axbZ0Z_1 ));
    InMux I__9450 (
            .O(N__42443),
            .I(N__42440));
    LocalMux I__9449 (
            .O(N__42440),
            .I(N__42437));
    Span4Mux_v I__9448 (
            .O(N__42437),
            .I(N__42434));
    Span4Mux_h I__9447 (
            .O(N__42434),
            .I(N__42431));
    Odrv4 I__9446 (
            .O(N__42431),
            .I(\pid_front.error_1 ));
    InMux I__9445 (
            .O(N__42428),
            .I(\pid_front.error_cry_0 ));
    InMux I__9444 (
            .O(N__42425),
            .I(N__42412));
    InMux I__9443 (
            .O(N__42424),
            .I(N__42412));
    InMux I__9442 (
            .O(N__42423),
            .I(N__42412));
    InMux I__9441 (
            .O(N__42422),
            .I(N__42409));
    InMux I__9440 (
            .O(N__42421),
            .I(N__42402));
    InMux I__9439 (
            .O(N__42420),
            .I(N__42402));
    InMux I__9438 (
            .O(N__42419),
            .I(N__42402));
    LocalMux I__9437 (
            .O(N__42412),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__9436 (
            .O(N__42409),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    LocalMux I__9435 (
            .O(N__42402),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_0 ));
    CascadeMux I__9434 (
            .O(N__42395),
            .I(N__42392));
    InMux I__9433 (
            .O(N__42392),
            .I(N__42389));
    LocalMux I__9432 (
            .O(N__42389),
            .I(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ));
    InMux I__9431 (
            .O(N__42386),
            .I(N__42383));
    LocalMux I__9430 (
            .O(N__42383),
            .I(N__42380));
    Span4Mux_v I__9429 (
            .O(N__42380),
            .I(N__42377));
    Span4Mux_h I__9428 (
            .O(N__42377),
            .I(N__42374));
    Odrv4 I__9427 (
            .O(N__42374),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ));
    InMux I__9426 (
            .O(N__42371),
            .I(N__42368));
    LocalMux I__9425 (
            .O(N__42368),
            .I(N__42365));
    Span4Mux_v I__9424 (
            .O(N__42365),
            .I(N__42362));
    Odrv4 I__9423 (
            .O(N__42362),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ));
    InMux I__9422 (
            .O(N__42359),
            .I(N__42356));
    LocalMux I__9421 (
            .O(N__42356),
            .I(\ppm_encoder_1.pulses2countZ0Z_2 ));
    InMux I__9420 (
            .O(N__42353),
            .I(N__42350));
    LocalMux I__9419 (
            .O(N__42350),
            .I(N__42347));
    Span4Mux_v I__9418 (
            .O(N__42347),
            .I(N__42344));
    Odrv4 I__9417 (
            .O(N__42344),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ));
    CascadeMux I__9416 (
            .O(N__42341),
            .I(N__42338));
    InMux I__9415 (
            .O(N__42338),
            .I(N__42335));
    LocalMux I__9414 (
            .O(N__42335),
            .I(\ppm_encoder_1.pulses2countZ0Z_3 ));
    InMux I__9413 (
            .O(N__42332),
            .I(N__42329));
    LocalMux I__9412 (
            .O(N__42329),
            .I(N__42326));
    Span4Mux_v I__9411 (
            .O(N__42326),
            .I(N__42323));
    Odrv4 I__9410 (
            .O(N__42323),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ));
    InMux I__9409 (
            .O(N__42320),
            .I(N__42317));
    LocalMux I__9408 (
            .O(N__42317),
            .I(\ppm_encoder_1.pulses2countZ0Z_0 ));
    InMux I__9407 (
            .O(N__42314),
            .I(N__42311));
    LocalMux I__9406 (
            .O(N__42311),
            .I(N__42308));
    Span4Mux_v I__9405 (
            .O(N__42308),
            .I(N__42305));
    Odrv4 I__9404 (
            .O(N__42305),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ));
    InMux I__9403 (
            .O(N__42302),
            .I(N__42299));
    LocalMux I__9402 (
            .O(N__42299),
            .I(N__42296));
    Span4Mux_h I__9401 (
            .O(N__42296),
            .I(N__42293));
    Span4Mux_v I__9400 (
            .O(N__42293),
            .I(N__42290));
    Odrv4 I__9399 (
            .O(N__42290),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ));
    CascadeMux I__9398 (
            .O(N__42287),
            .I(N__42284));
    InMux I__9397 (
            .O(N__42284),
            .I(N__42281));
    LocalMux I__9396 (
            .O(N__42281),
            .I(\ppm_encoder_1.pulses2countZ0Z_1 ));
    InMux I__9395 (
            .O(N__42278),
            .I(N__42273));
    InMux I__9394 (
            .O(N__42277),
            .I(N__42270));
    InMux I__9393 (
            .O(N__42276),
            .I(N__42267));
    LocalMux I__9392 (
            .O(N__42273),
            .I(N__42264));
    LocalMux I__9391 (
            .O(N__42270),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    LocalMux I__9390 (
            .O(N__42267),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    Odrv4 I__9389 (
            .O(N__42264),
            .I(\ppm_encoder_1.aileronZ0Z_3 ));
    InMux I__9388 (
            .O(N__42257),
            .I(N__42254));
    LocalMux I__9387 (
            .O(N__42254),
            .I(N__42251));
    Span4Mux_v I__9386 (
            .O(N__42251),
            .I(N__42248));
    Span4Mux_h I__9385 (
            .O(N__42248),
            .I(N__42245));
    Odrv4 I__9384 (
            .O(N__42245),
            .I(\ppm_encoder_1.N_289 ));
    InMux I__9383 (
            .O(N__42242),
            .I(N__42239));
    LocalMux I__9382 (
            .O(N__42239),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ));
    CascadeMux I__9381 (
            .O(N__42236),
            .I(\ppm_encoder_1.PPM_STATE_53_d_cascade_ ));
    InMux I__9380 (
            .O(N__42233),
            .I(N__42230));
    LocalMux I__9379 (
            .O(N__42230),
            .I(N__42227));
    Span4Mux_h I__9378 (
            .O(N__42227),
            .I(N__42224));
    Odrv4 I__9377 (
            .O(N__42224),
            .I(\ppm_encoder_1.N_134_0 ));
    InMux I__9376 (
            .O(N__42221),
            .I(N__42214));
    InMux I__9375 (
            .O(N__42220),
            .I(N__42209));
    InMux I__9374 (
            .O(N__42219),
            .I(N__42209));
    CascadeMux I__9373 (
            .O(N__42218),
            .I(N__42206));
    InMux I__9372 (
            .O(N__42217),
            .I(N__42201));
    LocalMux I__9371 (
            .O(N__42214),
            .I(N__42196));
    LocalMux I__9370 (
            .O(N__42209),
            .I(N__42196));
    InMux I__9369 (
            .O(N__42206),
            .I(N__42189));
    InMux I__9368 (
            .O(N__42205),
            .I(N__42189));
    InMux I__9367 (
            .O(N__42204),
            .I(N__42189));
    LocalMux I__9366 (
            .O(N__42201),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    Odrv12 I__9365 (
            .O(N__42196),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    LocalMux I__9364 (
            .O(N__42189),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ));
    InMux I__9363 (
            .O(N__42182),
            .I(N__42179));
    LocalMux I__9362 (
            .O(N__42179),
            .I(N__42176));
    Span12Mux_v I__9361 (
            .O(N__42176),
            .I(N__42168));
    InMux I__9360 (
            .O(N__42175),
            .I(N__42165));
    InMux I__9359 (
            .O(N__42174),
            .I(N__42162));
    InMux I__9358 (
            .O(N__42173),
            .I(N__42155));
    InMux I__9357 (
            .O(N__42172),
            .I(N__42155));
    InMux I__9356 (
            .O(N__42171),
            .I(N__42155));
    Odrv12 I__9355 (
            .O(N__42168),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__9354 (
            .O(N__42165),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__9353 (
            .O(N__42162),
            .I(\ppm_encoder_1.N_221 ));
    LocalMux I__9352 (
            .O(N__42155),
            .I(\ppm_encoder_1.N_221 ));
    CascadeMux I__9351 (
            .O(N__42146),
            .I(\ppm_encoder_1.N_232_cascade_ ));
    IoInMux I__9350 (
            .O(N__42143),
            .I(N__42140));
    LocalMux I__9349 (
            .O(N__42140),
            .I(N__42137));
    Span12Mux_s1_v I__9348 (
            .O(N__42137),
            .I(N__42134));
    Span12Mux_v I__9347 (
            .O(N__42134),
            .I(N__42131));
    Odrv12 I__9346 (
            .O(N__42131),
            .I(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ));
    InMux I__9345 (
            .O(N__42128),
            .I(N__42125));
    LocalMux I__9344 (
            .O(N__42125),
            .I(N__42122));
    Span4Mux_h I__9343 (
            .O(N__42122),
            .I(N__42119));
    Span4Mux_h I__9342 (
            .O(N__42119),
            .I(N__42116));
    Odrv4 I__9341 (
            .O(N__42116),
            .I(\ppm_encoder_1.N_139 ));
    InMux I__9340 (
            .O(N__42113),
            .I(N__42107));
    InMux I__9339 (
            .O(N__42112),
            .I(N__42107));
    LocalMux I__9338 (
            .O(N__42107),
            .I(\ppm_encoder_1.N_232 ));
    InMux I__9337 (
            .O(N__42104),
            .I(N__42101));
    LocalMux I__9336 (
            .O(N__42101),
            .I(N__42098));
    Span4Mux_h I__9335 (
            .O(N__42098),
            .I(N__42094));
    InMux I__9334 (
            .O(N__42097),
            .I(N__42091));
    Span4Mux_v I__9333 (
            .O(N__42094),
            .I(N__42088));
    LocalMux I__9332 (
            .O(N__42091),
            .I(N__42081));
    Span4Mux_h I__9331 (
            .O(N__42088),
            .I(N__42081));
    InMux I__9330 (
            .O(N__42087),
            .I(N__42078));
    InMux I__9329 (
            .O(N__42086),
            .I(N__42075));
    Odrv4 I__9328 (
            .O(N__42081),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__9327 (
            .O(N__42078),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    LocalMux I__9326 (
            .O(N__42075),
            .I(\ppm_encoder_1.PPM_STATEZ0Z_1 ));
    InMux I__9325 (
            .O(N__42068),
            .I(N__42065));
    LocalMux I__9324 (
            .O(N__42065),
            .I(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ));
    CascadeMux I__9323 (
            .O(N__42062),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ));
    CascadeMux I__9322 (
            .O(N__42059),
            .I(N__42055));
    InMux I__9321 (
            .O(N__42058),
            .I(N__42052));
    InMux I__9320 (
            .O(N__42055),
            .I(N__42049));
    LocalMux I__9319 (
            .O(N__42052),
            .I(N__42046));
    LocalMux I__9318 (
            .O(N__42049),
            .I(N__42040));
    Span4Mux_v I__9317 (
            .O(N__42046),
            .I(N__42040));
    InMux I__9316 (
            .O(N__42045),
            .I(N__42037));
    Odrv4 I__9315 (
            .O(N__42040),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    LocalMux I__9314 (
            .O(N__42037),
            .I(\ppm_encoder_1.un1_init_pulses_0 ));
    InMux I__9313 (
            .O(N__42032),
            .I(N__42029));
    LocalMux I__9312 (
            .O(N__42029),
            .I(N__42026));
    Span4Mux_h I__9311 (
            .O(N__42026),
            .I(N__42023));
    Odrv4 I__9310 (
            .O(N__42023),
            .I(\ppm_encoder_1.un1_init_pulses_10_0 ));
    InMux I__9309 (
            .O(N__42020),
            .I(N__42017));
    LocalMux I__9308 (
            .O(N__42017),
            .I(N__42012));
    InMux I__9307 (
            .O(N__42016),
            .I(N__42009));
    InMux I__9306 (
            .O(N__42015),
            .I(N__42006));
    Span4Mux_v I__9305 (
            .O(N__42012),
            .I(N__42003));
    LocalMux I__9304 (
            .O(N__42009),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    LocalMux I__9303 (
            .O(N__42006),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    Odrv4 I__9302 (
            .O(N__42003),
            .I(\ppm_encoder_1.throttleZ0Z_3 ));
    InMux I__9301 (
            .O(N__41996),
            .I(N__41992));
    InMux I__9300 (
            .O(N__41995),
            .I(N__41989));
    LocalMux I__9299 (
            .O(N__41992),
            .I(N__41986));
    LocalMux I__9298 (
            .O(N__41989),
            .I(N__41983));
    Span4Mux_h I__9297 (
            .O(N__41986),
            .I(N__41980));
    Odrv12 I__9296 (
            .O(N__41983),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    Odrv4 I__9295 (
            .O(N__41980),
            .I(\ppm_encoder_1.un1_init_pulses_0_3 ));
    InMux I__9294 (
            .O(N__41975),
            .I(N__41972));
    LocalMux I__9293 (
            .O(N__41972),
            .I(N__41967));
    CascadeMux I__9292 (
            .O(N__41971),
            .I(N__41964));
    InMux I__9291 (
            .O(N__41970),
            .I(N__41961));
    Span4Mux_v I__9290 (
            .O(N__41967),
            .I(N__41958));
    InMux I__9289 (
            .O(N__41964),
            .I(N__41955));
    LocalMux I__9288 (
            .O(N__41961),
            .I(N__41952));
    Span4Mux_h I__9287 (
            .O(N__41958),
            .I(N__41949));
    LocalMux I__9286 (
            .O(N__41955),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    Odrv4 I__9285 (
            .O(N__41952),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    Odrv4 I__9284 (
            .O(N__41949),
            .I(\ppm_encoder_1.elevatorZ0Z_3 ));
    CascadeMux I__9283 (
            .O(N__41942),
            .I(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ));
    CascadeMux I__9282 (
            .O(N__41939),
            .I(N__41936));
    InMux I__9281 (
            .O(N__41936),
            .I(N__41933));
    LocalMux I__9280 (
            .O(N__41933),
            .I(N__41930));
    Span4Mux_h I__9279 (
            .O(N__41930),
            .I(N__41927));
    Span4Mux_v I__9278 (
            .O(N__41927),
            .I(N__41924));
    Odrv4 I__9277 (
            .O(N__41924),
            .I(\ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ));
    InMux I__9276 (
            .O(N__41921),
            .I(N__41916));
    InMux I__9275 (
            .O(N__41920),
            .I(N__41913));
    InMux I__9274 (
            .O(N__41919),
            .I(N__41910));
    LocalMux I__9273 (
            .O(N__41916),
            .I(N__41905));
    LocalMux I__9272 (
            .O(N__41913),
            .I(N__41905));
    LocalMux I__9271 (
            .O(N__41910),
            .I(N__41902));
    Span4Mux_v I__9270 (
            .O(N__41905),
            .I(N__41899));
    Span4Mux_h I__9269 (
            .O(N__41902),
            .I(N__41896));
    Odrv4 I__9268 (
            .O(N__41899),
            .I(\pid_side.pid_preregZ0Z_0 ));
    Odrv4 I__9267 (
            .O(N__41896),
            .I(\pid_side.pid_preregZ0Z_0 ));
    CEMux I__9266 (
            .O(N__41891),
            .I(N__41887));
    CEMux I__9265 (
            .O(N__41890),
            .I(N__41884));
    LocalMux I__9264 (
            .O(N__41887),
            .I(N__41881));
    LocalMux I__9263 (
            .O(N__41884),
            .I(N__41878));
    Span4Mux_h I__9262 (
            .O(N__41881),
            .I(N__41875));
    Span4Mux_h I__9261 (
            .O(N__41878),
            .I(N__41872));
    Span4Mux_v I__9260 (
            .O(N__41875),
            .I(N__41869));
    Span4Mux_h I__9259 (
            .O(N__41872),
            .I(N__41866));
    Odrv4 I__9258 (
            .O(N__41869),
            .I(\pid_side.state_0_0 ));
    Odrv4 I__9257 (
            .O(N__41866),
            .I(\pid_side.state_0_0 ));
    CascadeMux I__9256 (
            .O(N__41861),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ));
    InMux I__9255 (
            .O(N__41858),
            .I(N__41855));
    LocalMux I__9254 (
            .O(N__41855),
            .I(N__41852));
    Span4Mux_h I__9253 (
            .O(N__41852),
            .I(N__41848));
    InMux I__9252 (
            .O(N__41851),
            .I(N__41845));
    Odrv4 I__9251 (
            .O(N__41848),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    LocalMux I__9250 (
            .O(N__41845),
            .I(\ppm_encoder_1.un1_init_pulses_0_14 ));
    CascadeMux I__9249 (
            .O(N__41840),
            .I(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ));
    CascadeMux I__9248 (
            .O(N__41837),
            .I(N__41834));
    InMux I__9247 (
            .O(N__41834),
            .I(N__41831));
    LocalMux I__9246 (
            .O(N__41831),
            .I(N__41828));
    Span4Mux_h I__9245 (
            .O(N__41828),
            .I(N__41825));
    Odrv4 I__9244 (
            .O(N__41825),
            .I(\ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ));
    InMux I__9243 (
            .O(N__41822),
            .I(N__41819));
    LocalMux I__9242 (
            .O(N__41819),
            .I(\ppm_encoder_1.un2_throttle_iv_1_14 ));
    InMux I__9241 (
            .O(N__41816),
            .I(N__41810));
    InMux I__9240 (
            .O(N__41815),
            .I(N__41810));
    LocalMux I__9239 (
            .O(N__41810),
            .I(N__41807));
    Span4Mux_h I__9238 (
            .O(N__41807),
            .I(N__41804));
    Span4Mux_h I__9237 (
            .O(N__41804),
            .I(N__41801));
    Odrv4 I__9236 (
            .O(N__41801),
            .I(\ppm_encoder_1.throttleZ0Z_14 ));
    InMux I__9235 (
            .O(N__41798),
            .I(N__41792));
    InMux I__9234 (
            .O(N__41797),
            .I(N__41792));
    LocalMux I__9233 (
            .O(N__41792),
            .I(N__41789));
    Span12Mux_v I__9232 (
            .O(N__41789),
            .I(N__41786));
    Odrv12 I__9231 (
            .O(N__41786),
            .I(\ppm_encoder_1.elevatorZ0Z_14 ));
    CascadeMux I__9230 (
            .O(N__41783),
            .I(\ppm_encoder_1.N_300_cascade_ ));
    InMux I__9229 (
            .O(N__41780),
            .I(N__41774));
    InMux I__9228 (
            .O(N__41779),
            .I(N__41774));
    LocalMux I__9227 (
            .O(N__41774),
            .I(N__41771));
    Span4Mux_h I__9226 (
            .O(N__41771),
            .I(N__41768));
    Odrv4 I__9225 (
            .O(N__41768),
            .I(\ppm_encoder_1.aileronZ0Z_14 ));
    CascadeMux I__9224 (
            .O(N__41765),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_ ));
    InMux I__9223 (
            .O(N__41762),
            .I(N__41759));
    LocalMux I__9222 (
            .O(N__41759),
            .I(N__41756));
    Odrv4 I__9221 (
            .O(N__41756),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ));
    InMux I__9220 (
            .O(N__41753),
            .I(N__41750));
    LocalMux I__9219 (
            .O(N__41750),
            .I(\ppm_encoder_1.pulses2countZ0Z_14 ));
    CascadeMux I__9218 (
            .O(N__41747),
            .I(N__41742));
    InMux I__9217 (
            .O(N__41746),
            .I(N__41738));
    InMux I__9216 (
            .O(N__41745),
            .I(N__41735));
    InMux I__9215 (
            .O(N__41742),
            .I(N__41730));
    InMux I__9214 (
            .O(N__41741),
            .I(N__41730));
    LocalMux I__9213 (
            .O(N__41738),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__9212 (
            .O(N__41735),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    LocalMux I__9211 (
            .O(N__41730),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ));
    InMux I__9210 (
            .O(N__41723),
            .I(N__41717));
    InMux I__9209 (
            .O(N__41722),
            .I(N__41714));
    InMux I__9208 (
            .O(N__41721),
            .I(N__41709));
    InMux I__9207 (
            .O(N__41720),
            .I(N__41709));
    LocalMux I__9206 (
            .O(N__41717),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__9205 (
            .O(N__41714),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    LocalMux I__9204 (
            .O(N__41709),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ));
    CascadeMux I__9203 (
            .O(N__41702),
            .I(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ));
    InMux I__9202 (
            .O(N__41699),
            .I(N__41696));
    LocalMux I__9201 (
            .O(N__41696),
            .I(\ppm_encoder_1.un2_throttle_iv_0_0 ));
    InMux I__9200 (
            .O(N__41693),
            .I(N__41688));
    InMux I__9199 (
            .O(N__41692),
            .I(N__41685));
    CascadeMux I__9198 (
            .O(N__41691),
            .I(N__41682));
    LocalMux I__9197 (
            .O(N__41688),
            .I(N__41679));
    LocalMux I__9196 (
            .O(N__41685),
            .I(N__41676));
    InMux I__9195 (
            .O(N__41682),
            .I(N__41673));
    Span4Mux_v I__9194 (
            .O(N__41679),
            .I(N__41668));
    Span4Mux_v I__9193 (
            .O(N__41676),
            .I(N__41668));
    LocalMux I__9192 (
            .O(N__41673),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    Odrv4 I__9191 (
            .O(N__41668),
            .I(\ppm_encoder_1.rudderZ0Z_13 ));
    InMux I__9190 (
            .O(N__41663),
            .I(N__41660));
    LocalMux I__9189 (
            .O(N__41660),
            .I(N__41656));
    InMux I__9188 (
            .O(N__41659),
            .I(N__41653));
    Odrv4 I__9187 (
            .O(N__41656),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    LocalMux I__9186 (
            .O(N__41653),
            .I(\ppm_encoder_1.un1_init_pulses_0_13 ));
    CascadeMux I__9185 (
            .O(N__41648),
            .I(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ));
    CascadeMux I__9184 (
            .O(N__41645),
            .I(N__41642));
    InMux I__9183 (
            .O(N__41642),
            .I(N__41639));
    LocalMux I__9182 (
            .O(N__41639),
            .I(N__41636));
    Span4Mux_v I__9181 (
            .O(N__41636),
            .I(N__41633));
    Odrv4 I__9180 (
            .O(N__41633),
            .I(\ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ));
    InMux I__9179 (
            .O(N__41630),
            .I(N__41627));
    LocalMux I__9178 (
            .O(N__41627),
            .I(\ppm_encoder_1.un2_throttle_iv_1_13 ));
    CascadeMux I__9177 (
            .O(N__41624),
            .I(\ppm_encoder_1.N_299_cascade_ ));
    CascadeMux I__9176 (
            .O(N__41621),
            .I(N__41617));
    CascadeMux I__9175 (
            .O(N__41620),
            .I(N__41614));
    InMux I__9174 (
            .O(N__41617),
            .I(N__41611));
    InMux I__9173 (
            .O(N__41614),
            .I(N__41608));
    LocalMux I__9172 (
            .O(N__41611),
            .I(N__41605));
    LocalMux I__9171 (
            .O(N__41608),
            .I(N__41602));
    Span4Mux_v I__9170 (
            .O(N__41605),
            .I(N__41599));
    Odrv4 I__9169 (
            .O(N__41602),
            .I(side_order_13));
    Odrv4 I__9168 (
            .O(N__41599),
            .I(side_order_13));
    InMux I__9167 (
            .O(N__41594),
            .I(N__41591));
    LocalMux I__9166 (
            .O(N__41591),
            .I(N__41588));
    Span4Mux_h I__9165 (
            .O(N__41588),
            .I(N__41585));
    Odrv4 I__9164 (
            .O(N__41585),
            .I(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ));
    InMux I__9163 (
            .O(N__41582),
            .I(N__41573));
    InMux I__9162 (
            .O(N__41581),
            .I(N__41573));
    InMux I__9161 (
            .O(N__41580),
            .I(N__41573));
    LocalMux I__9160 (
            .O(N__41573),
            .I(\ppm_encoder_1.aileronZ0Z_13 ));
    InMux I__9159 (
            .O(N__41570),
            .I(N__41567));
    LocalMux I__9158 (
            .O(N__41567),
            .I(N__41564));
    Span4Mux_v I__9157 (
            .O(N__41564),
            .I(N__41561));
    Span4Mux_v I__9156 (
            .O(N__41561),
            .I(N__41557));
    InMux I__9155 (
            .O(N__41560),
            .I(N__41554));
    Sp12to4 I__9154 (
            .O(N__41557),
            .I(N__41549));
    LocalMux I__9153 (
            .O(N__41554),
            .I(N__41549));
    Odrv12 I__9152 (
            .O(N__41549),
            .I(front_order_13));
    InMux I__9151 (
            .O(N__41546),
            .I(N__41543));
    LocalMux I__9150 (
            .O(N__41543),
            .I(N__41540));
    Span4Mux_h I__9149 (
            .O(N__41540),
            .I(N__41537));
    Span4Mux_v I__9148 (
            .O(N__41537),
            .I(N__41534));
    Odrv4 I__9147 (
            .O(N__41534),
            .I(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ));
    InMux I__9146 (
            .O(N__41531),
            .I(N__41522));
    InMux I__9145 (
            .O(N__41530),
            .I(N__41522));
    InMux I__9144 (
            .O(N__41529),
            .I(N__41522));
    LocalMux I__9143 (
            .O(N__41522),
            .I(\ppm_encoder_1.elevatorZ0Z_13 ));
    InMux I__9142 (
            .O(N__41519),
            .I(N__41516));
    LocalMux I__9141 (
            .O(N__41516),
            .I(N__41513));
    Span4Mux_h I__9140 (
            .O(N__41513),
            .I(N__41509));
    CascadeMux I__9139 (
            .O(N__41512),
            .I(N__41506));
    Span4Mux_h I__9138 (
            .O(N__41509),
            .I(N__41503));
    InMux I__9137 (
            .O(N__41506),
            .I(N__41500));
    Odrv4 I__9136 (
            .O(N__41503),
            .I(throttle_order_13));
    LocalMux I__9135 (
            .O(N__41500),
            .I(throttle_order_13));
    InMux I__9134 (
            .O(N__41495),
            .I(N__41492));
    LocalMux I__9133 (
            .O(N__41492),
            .I(N__41489));
    Odrv12 I__9132 (
            .O(N__41489),
            .I(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ));
    CascadeMux I__9131 (
            .O(N__41486),
            .I(N__41481));
    InMux I__9130 (
            .O(N__41485),
            .I(N__41476));
    InMux I__9129 (
            .O(N__41484),
            .I(N__41476));
    InMux I__9128 (
            .O(N__41481),
            .I(N__41473));
    LocalMux I__9127 (
            .O(N__41476),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    LocalMux I__9126 (
            .O(N__41473),
            .I(\ppm_encoder_1.throttleZ0Z_13 ));
    InMux I__9125 (
            .O(N__41468),
            .I(N__41464));
    InMux I__9124 (
            .O(N__41467),
            .I(N__41461));
    LocalMux I__9123 (
            .O(N__41464),
            .I(N__41458));
    LocalMux I__9122 (
            .O(N__41461),
            .I(N__41453));
    Span4Mux_v I__9121 (
            .O(N__41458),
            .I(N__41453));
    Span4Mux_h I__9120 (
            .O(N__41453),
            .I(N__41450));
    Odrv4 I__9119 (
            .O(N__41450),
            .I(\ppm_encoder_1.rudderZ0Z_14 ));
    InMux I__9118 (
            .O(N__41447),
            .I(N__41444));
    LocalMux I__9117 (
            .O(N__41444),
            .I(N__41436));
    InMux I__9116 (
            .O(N__41443),
            .I(N__41433));
    InMux I__9115 (
            .O(N__41442),
            .I(N__41424));
    InMux I__9114 (
            .O(N__41441),
            .I(N__41424));
    InMux I__9113 (
            .O(N__41440),
            .I(N__41424));
    InMux I__9112 (
            .O(N__41439),
            .I(N__41424));
    Odrv4 I__9111 (
            .O(N__41436),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__9110 (
            .O(N__41433),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    LocalMux I__9109 (
            .O(N__41424),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ));
    CascadeMux I__9108 (
            .O(N__41417),
            .I(N__41413));
    InMux I__9107 (
            .O(N__41416),
            .I(N__41410));
    InMux I__9106 (
            .O(N__41413),
            .I(N__41406));
    LocalMux I__9105 (
            .O(N__41410),
            .I(N__41402));
    InMux I__9104 (
            .O(N__41409),
            .I(N__41399));
    LocalMux I__9103 (
            .O(N__41406),
            .I(N__41396));
    InMux I__9102 (
            .O(N__41405),
            .I(N__41393));
    Span4Mux_v I__9101 (
            .O(N__41402),
            .I(N__41388));
    LocalMux I__9100 (
            .O(N__41399),
            .I(N__41388));
    Odrv4 I__9099 (
            .O(N__41396),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    LocalMux I__9098 (
            .O(N__41393),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    Odrv4 I__9097 (
            .O(N__41388),
            .I(\ppm_encoder_1.init_pulsesZ0Z_0 ));
    CascadeMux I__9096 (
            .O(N__41381),
            .I(N__41378));
    InMux I__9095 (
            .O(N__41378),
            .I(N__41375));
    LocalMux I__9094 (
            .O(N__41375),
            .I(\ppm_encoder_1.un1_init_pulses_11_0 ));
    InMux I__9093 (
            .O(N__41372),
            .I(N__41369));
    LocalMux I__9092 (
            .O(N__41369),
            .I(N__41364));
    InMux I__9091 (
            .O(N__41368),
            .I(N__41361));
    CascadeMux I__9090 (
            .O(N__41367),
            .I(N__41358));
    Span4Mux_v I__9089 (
            .O(N__41364),
            .I(N__41353));
    LocalMux I__9088 (
            .O(N__41361),
            .I(N__41353));
    InMux I__9087 (
            .O(N__41358),
            .I(N__41350));
    Odrv4 I__9086 (
            .O(N__41353),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    LocalMux I__9085 (
            .O(N__41350),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_6 ));
    InMux I__9084 (
            .O(N__41345),
            .I(N__41341));
    CascadeMux I__9083 (
            .O(N__41344),
            .I(N__41338));
    LocalMux I__9082 (
            .O(N__41341),
            .I(N__41334));
    InMux I__9081 (
            .O(N__41338),
            .I(N__41329));
    InMux I__9080 (
            .O(N__41337),
            .I(N__41329));
    Span4Mux_v I__9079 (
            .O(N__41334),
            .I(N__41318));
    LocalMux I__9078 (
            .O(N__41329),
            .I(N__41318));
    InMux I__9077 (
            .O(N__41328),
            .I(N__41309));
    InMux I__9076 (
            .O(N__41327),
            .I(N__41309));
    InMux I__9075 (
            .O(N__41326),
            .I(N__41309));
    InMux I__9074 (
            .O(N__41325),
            .I(N__41309));
    InMux I__9073 (
            .O(N__41324),
            .I(N__41306));
    InMux I__9072 (
            .O(N__41323),
            .I(N__41303));
    Span4Mux_h I__9071 (
            .O(N__41318),
            .I(N__41298));
    LocalMux I__9070 (
            .O(N__41309),
            .I(N__41298));
    LocalMux I__9069 (
            .O(N__41306),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    LocalMux I__9068 (
            .O(N__41303),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    Odrv4 I__9067 (
            .O(N__41298),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ));
    CascadeMux I__9066 (
            .O(N__41291),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ));
    InMux I__9065 (
            .O(N__41288),
            .I(N__41285));
    LocalMux I__9064 (
            .O(N__41285),
            .I(N__41282));
    Span4Mux_h I__9063 (
            .O(N__41282),
            .I(N__41279));
    Odrv4 I__9062 (
            .O(N__41279),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ));
    CascadeMux I__9061 (
            .O(N__41276),
            .I(N__41271));
    CascadeMux I__9060 (
            .O(N__41275),
            .I(N__41267));
    CascadeMux I__9059 (
            .O(N__41274),
            .I(N__41264));
    InMux I__9058 (
            .O(N__41271),
            .I(N__41256));
    InMux I__9057 (
            .O(N__41270),
            .I(N__41256));
    InMux I__9056 (
            .O(N__41267),
            .I(N__41251));
    InMux I__9055 (
            .O(N__41264),
            .I(N__41251));
    InMux I__9054 (
            .O(N__41263),
            .I(N__41248));
    InMux I__9053 (
            .O(N__41262),
            .I(N__41243));
    InMux I__9052 (
            .O(N__41261),
            .I(N__41243));
    LocalMux I__9051 (
            .O(N__41256),
            .I(N__41240));
    LocalMux I__9050 (
            .O(N__41251),
            .I(N__41237));
    LocalMux I__9049 (
            .O(N__41248),
            .I(N__41234));
    LocalMux I__9048 (
            .O(N__41243),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__9047 (
            .O(N__41240),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv4 I__9046 (
            .O(N__41237),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    Odrv12 I__9045 (
            .O(N__41234),
            .I(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ));
    InMux I__9044 (
            .O(N__41225),
            .I(N__41222));
    LocalMux I__9043 (
            .O(N__41222),
            .I(N__41217));
    InMux I__9042 (
            .O(N__41221),
            .I(N__41212));
    InMux I__9041 (
            .O(N__41220),
            .I(N__41212));
    Odrv12 I__9040 (
            .O(N__41217),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    LocalMux I__9039 (
            .O(N__41212),
            .I(\ppm_encoder_1.init_pulsesZ0Z_3 ));
    InMux I__9038 (
            .O(N__41207),
            .I(N__41204));
    LocalMux I__9037 (
            .O(N__41204),
            .I(N__41199));
    InMux I__9036 (
            .O(N__41203),
            .I(N__41196));
    CascadeMux I__9035 (
            .O(N__41202),
            .I(N__41193));
    Span4Mux_v I__9034 (
            .O(N__41199),
            .I(N__41189));
    LocalMux I__9033 (
            .O(N__41196),
            .I(N__41186));
    InMux I__9032 (
            .O(N__41193),
            .I(N__41183));
    InMux I__9031 (
            .O(N__41192),
            .I(N__41180));
    Span4Mux_h I__9030 (
            .O(N__41189),
            .I(N__41175));
    Span4Mux_h I__9029 (
            .O(N__41186),
            .I(N__41175));
    LocalMux I__9028 (
            .O(N__41183),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    LocalMux I__9027 (
            .O(N__41180),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    Odrv4 I__9026 (
            .O(N__41175),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ));
    InMux I__9025 (
            .O(N__41168),
            .I(N__41163));
    InMux I__9024 (
            .O(N__41167),
            .I(N__41160));
    InMux I__9023 (
            .O(N__41166),
            .I(N__41157));
    LocalMux I__9022 (
            .O(N__41163),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    LocalMux I__9021 (
            .O(N__41160),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    LocalMux I__9020 (
            .O(N__41157),
            .I(\ppm_encoder_1.init_pulsesZ0Z_10 ));
    InMux I__9019 (
            .O(N__41150),
            .I(N__41145));
    InMux I__9018 (
            .O(N__41149),
            .I(N__41142));
    CascadeMux I__9017 (
            .O(N__41148),
            .I(N__41139));
    LocalMux I__9016 (
            .O(N__41145),
            .I(N__41136));
    LocalMux I__9015 (
            .O(N__41142),
            .I(N__41133));
    InMux I__9014 (
            .O(N__41139),
            .I(N__41130));
    Span4Mux_h I__9013 (
            .O(N__41136),
            .I(N__41127));
    Span4Mux_v I__9012 (
            .O(N__41133),
            .I(N__41124));
    LocalMux I__9011 (
            .O(N__41130),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__9010 (
            .O(N__41127),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    Odrv4 I__9009 (
            .O(N__41124),
            .I(\ppm_encoder_1.rudderZ0Z_10 ));
    CascadeMux I__9008 (
            .O(N__41117),
            .I(N__41114));
    InMux I__9007 (
            .O(N__41114),
            .I(N__41108));
    InMux I__9006 (
            .O(N__41113),
            .I(N__41108));
    LocalMux I__9005 (
            .O(N__41108),
            .I(N__41104));
    CascadeMux I__9004 (
            .O(N__41107),
            .I(N__41101));
    Span4Mux_h I__9003 (
            .O(N__41104),
            .I(N__41098));
    InMux I__9002 (
            .O(N__41101),
            .I(N__41095));
    Span4Mux_v I__9001 (
            .O(N__41098),
            .I(N__41092));
    LocalMux I__9000 (
            .O(N__41095),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    Odrv4 I__8999 (
            .O(N__41092),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ));
    InMux I__8998 (
            .O(N__41087),
            .I(N__41084));
    LocalMux I__8997 (
            .O(N__41084),
            .I(N__41078));
    InMux I__8996 (
            .O(N__41083),
            .I(N__41074));
    InMux I__8995 (
            .O(N__41082),
            .I(N__41069));
    InMux I__8994 (
            .O(N__41081),
            .I(N__41069));
    Span4Mux_v I__8993 (
            .O(N__41078),
            .I(N__41066));
    InMux I__8992 (
            .O(N__41077),
            .I(N__41063));
    LocalMux I__8991 (
            .O(N__41074),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__8990 (
            .O(N__41069),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    Odrv4 I__8989 (
            .O(N__41066),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    LocalMux I__8988 (
            .O(N__41063),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ));
    InMux I__8987 (
            .O(N__41054),
            .I(N__41045));
    InMux I__8986 (
            .O(N__41053),
            .I(N__41045));
    InMux I__8985 (
            .O(N__41052),
            .I(N__41045));
    LocalMux I__8984 (
            .O(N__41045),
            .I(\ppm_encoder_1.init_pulsesZ0Z_4 ));
    InMux I__8983 (
            .O(N__41042),
            .I(N__41038));
    InMux I__8982 (
            .O(N__41041),
            .I(N__41035));
    LocalMux I__8981 (
            .O(N__41038),
            .I(N__41032));
    LocalMux I__8980 (
            .O(N__41035),
            .I(N__41029));
    Span4Mux_v I__8979 (
            .O(N__41032),
            .I(N__41026));
    Span12Mux_v I__8978 (
            .O(N__41029),
            .I(N__41023));
    Odrv4 I__8977 (
            .O(N__41026),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    Odrv12 I__8976 (
            .O(N__41023),
            .I(\ppm_encoder_1.rudderZ0Z_4 ));
    InMux I__8975 (
            .O(N__41018),
            .I(N__41015));
    LocalMux I__8974 (
            .O(N__41015),
            .I(N__41012));
    Span4Mux_h I__8973 (
            .O(N__41012),
            .I(N__41009));
    Odrv4 I__8972 (
            .O(N__41009),
            .I(\ppm_encoder_1.un1_init_pulses_10_5 ));
    CascadeMux I__8971 (
            .O(N__41006),
            .I(N__41003));
    InMux I__8970 (
            .O(N__41003),
            .I(N__41000));
    LocalMux I__8969 (
            .O(N__41000),
            .I(N__40997));
    Odrv4 I__8968 (
            .O(N__40997),
            .I(\ppm_encoder_1.un1_init_pulses_11_5 ));
    InMux I__8967 (
            .O(N__40994),
            .I(N__40990));
    CascadeMux I__8966 (
            .O(N__40993),
            .I(N__40987));
    LocalMux I__8965 (
            .O(N__40990),
            .I(N__40984));
    InMux I__8964 (
            .O(N__40987),
            .I(N__40980));
    Span4Mux_h I__8963 (
            .O(N__40984),
            .I(N__40977));
    InMux I__8962 (
            .O(N__40983),
            .I(N__40974));
    LocalMux I__8961 (
            .O(N__40980),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    Odrv4 I__8960 (
            .O(N__40977),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    LocalMux I__8959 (
            .O(N__40974),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ));
    InMux I__8958 (
            .O(N__40967),
            .I(N__40964));
    LocalMux I__8957 (
            .O(N__40964),
            .I(N__40959));
    InMux I__8956 (
            .O(N__40963),
            .I(N__40954));
    InMux I__8955 (
            .O(N__40962),
            .I(N__40954));
    Span4Mux_h I__8954 (
            .O(N__40959),
            .I(N__40951));
    LocalMux I__8953 (
            .O(N__40954),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    Odrv4 I__8952 (
            .O(N__40951),
            .I(\ppm_encoder_1.init_pulsesZ0Z_7 ));
    CascadeMux I__8951 (
            .O(N__40946),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ));
    InMux I__8950 (
            .O(N__40943),
            .I(N__40938));
    InMux I__8949 (
            .O(N__40942),
            .I(N__40933));
    InMux I__8948 (
            .O(N__40941),
            .I(N__40933));
    LocalMux I__8947 (
            .O(N__40938),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    LocalMux I__8946 (
            .O(N__40933),
            .I(\ppm_encoder_1.init_pulsesZ0Z_1 ));
    CascadeMux I__8945 (
            .O(N__40928),
            .I(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ));
    InMux I__8944 (
            .O(N__40925),
            .I(N__40921));
    InMux I__8943 (
            .O(N__40924),
            .I(N__40918));
    LocalMux I__8942 (
            .O(N__40921),
            .I(N__40915));
    LocalMux I__8941 (
            .O(N__40918),
            .I(N__40912));
    Span4Mux_h I__8940 (
            .O(N__40915),
            .I(N__40908));
    Span4Mux_h I__8939 (
            .O(N__40912),
            .I(N__40905));
    InMux I__8938 (
            .O(N__40911),
            .I(N__40902));
    Odrv4 I__8937 (
            .O(N__40908),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    Odrv4 I__8936 (
            .O(N__40905),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    LocalMux I__8935 (
            .O(N__40902),
            .I(\ppm_encoder_1.init_pulsesZ0Z_2 ));
    InMux I__8934 (
            .O(N__40895),
            .I(N__40892));
    LocalMux I__8933 (
            .O(N__40892),
            .I(N__40889));
    Sp12to4 I__8932 (
            .O(N__40889),
            .I(N__40884));
    InMux I__8931 (
            .O(N__40888),
            .I(N__40881));
    InMux I__8930 (
            .O(N__40887),
            .I(N__40878));
    Span12Mux_v I__8929 (
            .O(N__40884),
            .I(N__40873));
    LocalMux I__8928 (
            .O(N__40881),
            .I(N__40873));
    LocalMux I__8927 (
            .O(N__40878),
            .I(N__40870));
    Odrv12 I__8926 (
            .O(N__40873),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    Odrv12 I__8925 (
            .O(N__40870),
            .I(\ppm_encoder_1.init_pulsesZ0Z_12 ));
    InMux I__8924 (
            .O(N__40865),
            .I(N__40862));
    LocalMux I__8923 (
            .O(N__40862),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_12 ));
    InMux I__8922 (
            .O(N__40859),
            .I(N__40856));
    LocalMux I__8921 (
            .O(N__40856),
            .I(N__40853));
    Span4Mux_v I__8920 (
            .O(N__40853),
            .I(N__40850));
    Odrv4 I__8919 (
            .O(N__40850),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_18 ));
    InMux I__8918 (
            .O(N__40847),
            .I(N__40844));
    LocalMux I__8917 (
            .O(N__40844),
            .I(N__40841));
    Odrv4 I__8916 (
            .O(N__40841),
            .I(\ppm_encoder_1.un1_init_pulses_11_3 ));
    InMux I__8915 (
            .O(N__40838),
            .I(N__40835));
    LocalMux I__8914 (
            .O(N__40835),
            .I(N__40832));
    Span4Mux_h I__8913 (
            .O(N__40832),
            .I(N__40829));
    Odrv4 I__8912 (
            .O(N__40829),
            .I(\ppm_encoder_1.un1_init_pulses_10_3 ));
    CascadeMux I__8911 (
            .O(N__40826),
            .I(N__40823));
    InMux I__8910 (
            .O(N__40823),
            .I(N__40820));
    LocalMux I__8909 (
            .O(N__40820),
            .I(N__40817));
    Odrv4 I__8908 (
            .O(N__40817),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_3 ));
    InMux I__8907 (
            .O(N__40814),
            .I(N__40811));
    LocalMux I__8906 (
            .O(N__40811),
            .I(N__40808));
    Span4Mux_h I__8905 (
            .O(N__40808),
            .I(N__40805));
    Odrv4 I__8904 (
            .O(N__40805),
            .I(\ppm_encoder_1.un1_init_pulses_10_4 ));
    InMux I__8903 (
            .O(N__40802),
            .I(N__40799));
    LocalMux I__8902 (
            .O(N__40799),
            .I(N__40796));
    Odrv4 I__8901 (
            .O(N__40796),
            .I(\ppm_encoder_1.un1_init_pulses_11_4 ));
    InMux I__8900 (
            .O(N__40793),
            .I(N__40790));
    LocalMux I__8899 (
            .O(N__40790),
            .I(N__40786));
    InMux I__8898 (
            .O(N__40789),
            .I(N__40783));
    Span4Mux_v I__8897 (
            .O(N__40786),
            .I(N__40778));
    LocalMux I__8896 (
            .O(N__40783),
            .I(N__40778));
    Span4Mux_v I__8895 (
            .O(N__40778),
            .I(N__40775));
    Sp12to4 I__8894 (
            .O(N__40775),
            .I(N__40772));
    Odrv12 I__8893 (
            .O(N__40772),
            .I(\ppm_encoder_1.un1_init_pulses_0_4 ));
    InMux I__8892 (
            .O(N__40769),
            .I(N__40766));
    LocalMux I__8891 (
            .O(N__40766),
            .I(N__40763));
    Odrv4 I__8890 (
            .O(N__40763),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_4 ));
    InMux I__8889 (
            .O(N__40760),
            .I(N__40752));
    InMux I__8888 (
            .O(N__40759),
            .I(N__40752));
    InMux I__8887 (
            .O(N__40758),
            .I(N__40743));
    InMux I__8886 (
            .O(N__40757),
            .I(N__40743));
    LocalMux I__8885 (
            .O(N__40752),
            .I(N__40740));
    InMux I__8884 (
            .O(N__40751),
            .I(N__40731));
    InMux I__8883 (
            .O(N__40750),
            .I(N__40731));
    InMux I__8882 (
            .O(N__40749),
            .I(N__40731));
    InMux I__8881 (
            .O(N__40748),
            .I(N__40731));
    LocalMux I__8880 (
            .O(N__40743),
            .I(N__40728));
    Span4Mux_h I__8879 (
            .O(N__40740),
            .I(N__40725));
    LocalMux I__8878 (
            .O(N__40731),
            .I(N__40722));
    Span4Mux_h I__8877 (
            .O(N__40728),
            .I(N__40719));
    Odrv4 I__8876 (
            .O(N__40725),
            .I(\uart_pc.un1_state_2_0 ));
    Odrv4 I__8875 (
            .O(N__40722),
            .I(\uart_pc.un1_state_2_0 ));
    Odrv4 I__8874 (
            .O(N__40719),
            .I(\uart_pc.un1_state_2_0 ));
    CascadeMux I__8873 (
            .O(N__40712),
            .I(N__40708));
    CascadeMux I__8872 (
            .O(N__40711),
            .I(N__40701));
    InMux I__8871 (
            .O(N__40708),
            .I(N__40695));
    InMux I__8870 (
            .O(N__40707),
            .I(N__40695));
    IoInMux I__8869 (
            .O(N__40706),
            .I(N__40688));
    InMux I__8868 (
            .O(N__40705),
            .I(N__40685));
    InMux I__8867 (
            .O(N__40704),
            .I(N__40682));
    InMux I__8866 (
            .O(N__40701),
            .I(N__40677));
    InMux I__8865 (
            .O(N__40700),
            .I(N__40677));
    LocalMux I__8864 (
            .O(N__40695),
            .I(N__40673));
    InMux I__8863 (
            .O(N__40694),
            .I(N__40670));
    InMux I__8862 (
            .O(N__40693),
            .I(N__40663));
    InMux I__8861 (
            .O(N__40692),
            .I(N__40663));
    InMux I__8860 (
            .O(N__40691),
            .I(N__40663));
    LocalMux I__8859 (
            .O(N__40688),
            .I(N__40660));
    LocalMux I__8858 (
            .O(N__40685),
            .I(N__40657));
    LocalMux I__8857 (
            .O(N__40682),
            .I(N__40654));
    LocalMux I__8856 (
            .O(N__40677),
            .I(N__40651));
    CascadeMux I__8855 (
            .O(N__40676),
            .I(N__40647));
    Span4Mux_v I__8854 (
            .O(N__40673),
            .I(N__40644));
    LocalMux I__8853 (
            .O(N__40670),
            .I(N__40638));
    LocalMux I__8852 (
            .O(N__40663),
            .I(N__40638));
    Span4Mux_s2_v I__8851 (
            .O(N__40660),
            .I(N__40635));
    Span4Mux_h I__8850 (
            .O(N__40657),
            .I(N__40630));
    Span4Mux_v I__8849 (
            .O(N__40654),
            .I(N__40630));
    Span4Mux_h I__8848 (
            .O(N__40651),
            .I(N__40627));
    InMux I__8847 (
            .O(N__40650),
            .I(N__40624));
    InMux I__8846 (
            .O(N__40647),
            .I(N__40621));
    Sp12to4 I__8845 (
            .O(N__40644),
            .I(N__40618));
    InMux I__8844 (
            .O(N__40643),
            .I(N__40615));
    Span4Mux_v I__8843 (
            .O(N__40638),
            .I(N__40612));
    Span4Mux_h I__8842 (
            .O(N__40635),
            .I(N__40605));
    Span4Mux_v I__8841 (
            .O(N__40630),
            .I(N__40605));
    Span4Mux_v I__8840 (
            .O(N__40627),
            .I(N__40605));
    LocalMux I__8839 (
            .O(N__40624),
            .I(N__40596));
    LocalMux I__8838 (
            .O(N__40621),
            .I(N__40596));
    Span12Mux_h I__8837 (
            .O(N__40618),
            .I(N__40596));
    LocalMux I__8836 (
            .O(N__40615),
            .I(N__40596));
    Odrv4 I__8835 (
            .O(N__40612),
            .I(debug_CH2_18A_c));
    Odrv4 I__8834 (
            .O(N__40605),
            .I(debug_CH2_18A_c));
    Odrv12 I__8833 (
            .O(N__40596),
            .I(debug_CH2_18A_c));
    InMux I__8832 (
            .O(N__40589),
            .I(N__40586));
    LocalMux I__8831 (
            .O(N__40586),
            .I(N__40582));
    InMux I__8830 (
            .O(N__40585),
            .I(N__40579));
    Span4Mux_h I__8829 (
            .O(N__40582),
            .I(N__40576));
    LocalMux I__8828 (
            .O(N__40579),
            .I(N__40570));
    Span4Mux_h I__8827 (
            .O(N__40576),
            .I(N__40570));
    InMux I__8826 (
            .O(N__40575),
            .I(N__40567));
    Odrv4 I__8825 (
            .O(N__40570),
            .I(\uart_pc.N_152 ));
    LocalMux I__8824 (
            .O(N__40567),
            .I(\uart_pc.N_152 ));
    CascadeMux I__8823 (
            .O(N__40562),
            .I(N__40559));
    InMux I__8822 (
            .O(N__40559),
            .I(N__40556));
    LocalMux I__8821 (
            .O(N__40556),
            .I(N__40553));
    Span4Mux_h I__8820 (
            .O(N__40553),
            .I(N__40550));
    Span4Mux_h I__8819 (
            .O(N__40550),
            .I(N__40547));
    Span4Mux_h I__8818 (
            .O(N__40547),
            .I(N__40544));
    Span4Mux_v I__8817 (
            .O(N__40544),
            .I(N__40540));
    InMux I__8816 (
            .O(N__40543),
            .I(N__40537));
    Odrv4 I__8815 (
            .O(N__40540),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    LocalMux I__8814 (
            .O(N__40537),
            .I(\uart_pc.data_AuxZ0Z_7 ));
    SRMux I__8813 (
            .O(N__40532),
            .I(N__40529));
    LocalMux I__8812 (
            .O(N__40529),
            .I(N__40525));
    SRMux I__8811 (
            .O(N__40528),
            .I(N__40521));
    Span4Mux_h I__8810 (
            .O(N__40525),
            .I(N__40518));
    SRMux I__8809 (
            .O(N__40524),
            .I(N__40515));
    LocalMux I__8808 (
            .O(N__40521),
            .I(N__40512));
    Span4Mux_h I__8807 (
            .O(N__40518),
            .I(N__40509));
    LocalMux I__8806 (
            .O(N__40515),
            .I(N__40506));
    Span4Mux_h I__8805 (
            .O(N__40512),
            .I(N__40503));
    Odrv4 I__8804 (
            .O(N__40509),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv4 I__8803 (
            .O(N__40506),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    Odrv4 I__8802 (
            .O(N__40503),
            .I(\uart_pc.state_RNIEAGSZ0Z_4 ));
    InMux I__8801 (
            .O(N__40496),
            .I(N__40493));
    LocalMux I__8800 (
            .O(N__40493),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ));
    InMux I__8799 (
            .O(N__40490),
            .I(N__40487));
    LocalMux I__8798 (
            .O(N__40487),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ));
    InMux I__8797 (
            .O(N__40484),
            .I(N__40481));
    LocalMux I__8796 (
            .O(N__40481),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ));
    InMux I__8795 (
            .O(N__40478),
            .I(N__40475));
    LocalMux I__8794 (
            .O(N__40475),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_5 ));
    CascadeMux I__8793 (
            .O(N__40472),
            .I(N__40469));
    InMux I__8792 (
            .O(N__40469),
            .I(N__40466));
    LocalMux I__8791 (
            .O(N__40466),
            .I(N__40461));
    InMux I__8790 (
            .O(N__40465),
            .I(N__40456));
    InMux I__8789 (
            .O(N__40464),
            .I(N__40456));
    Odrv4 I__8788 (
            .O(N__40461),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    LocalMux I__8787 (
            .O(N__40456),
            .I(\ppm_encoder_1.init_pulsesZ0Z_13 ));
    CascadeMux I__8786 (
            .O(N__40451),
            .I(N__40448));
    InMux I__8785 (
            .O(N__40448),
            .I(N__40445));
    LocalMux I__8784 (
            .O(N__40445),
            .I(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ));
    CascadeMux I__8783 (
            .O(N__40442),
            .I(N__40439));
    InMux I__8782 (
            .O(N__40439),
            .I(N__40436));
    LocalMux I__8781 (
            .O(N__40436),
            .I(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ));
    InMux I__8780 (
            .O(N__40433),
            .I(N__40430));
    LocalMux I__8779 (
            .O(N__40430),
            .I(N__40427));
    Span4Mux_h I__8778 (
            .O(N__40427),
            .I(N__40422));
    InMux I__8777 (
            .O(N__40426),
            .I(N__40417));
    InMux I__8776 (
            .O(N__40425),
            .I(N__40417));
    Odrv4 I__8775 (
            .O(N__40422),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    LocalMux I__8774 (
            .O(N__40417),
            .I(\ppm_encoder_1.init_pulsesZ0Z_6 ));
    CascadeMux I__8773 (
            .O(N__40412),
            .I(N__40409));
    InMux I__8772 (
            .O(N__40409),
            .I(N__40406));
    LocalMux I__8771 (
            .O(N__40406),
            .I(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ));
    InMux I__8770 (
            .O(N__40403),
            .I(N__40397));
    InMux I__8769 (
            .O(N__40402),
            .I(N__40392));
    InMux I__8768 (
            .O(N__40401),
            .I(N__40389));
    InMux I__8767 (
            .O(N__40400),
            .I(N__40386));
    LocalMux I__8766 (
            .O(N__40397),
            .I(N__40383));
    InMux I__8765 (
            .O(N__40396),
            .I(N__40380));
    InMux I__8764 (
            .O(N__40395),
            .I(N__40375));
    LocalMux I__8763 (
            .O(N__40392),
            .I(N__40370));
    LocalMux I__8762 (
            .O(N__40389),
            .I(N__40370));
    LocalMux I__8761 (
            .O(N__40386),
            .I(N__40366));
    Span4Mux_v I__8760 (
            .O(N__40383),
            .I(N__40363));
    LocalMux I__8759 (
            .O(N__40380),
            .I(N__40360));
    InMux I__8758 (
            .O(N__40379),
            .I(N__40356));
    InMux I__8757 (
            .O(N__40378),
            .I(N__40353));
    LocalMux I__8756 (
            .O(N__40375),
            .I(N__40350));
    Span4Mux_h I__8755 (
            .O(N__40370),
            .I(N__40347));
    InMux I__8754 (
            .O(N__40369),
            .I(N__40344));
    Span4Mux_h I__8753 (
            .O(N__40366),
            .I(N__40341));
    Sp12to4 I__8752 (
            .O(N__40363),
            .I(N__40338));
    Span4Mux_h I__8751 (
            .O(N__40360),
            .I(N__40335));
    InMux I__8750 (
            .O(N__40359),
            .I(N__40332));
    LocalMux I__8749 (
            .O(N__40356),
            .I(N__40329));
    LocalMux I__8748 (
            .O(N__40353),
            .I(N__40324));
    Span4Mux_h I__8747 (
            .O(N__40350),
            .I(N__40324));
    Span4Mux_v I__8746 (
            .O(N__40347),
            .I(N__40317));
    LocalMux I__8745 (
            .O(N__40344),
            .I(N__40317));
    Span4Mux_h I__8744 (
            .O(N__40341),
            .I(N__40317));
    Span12Mux_h I__8743 (
            .O(N__40338),
            .I(N__40312));
    Sp12to4 I__8742 (
            .O(N__40335),
            .I(N__40312));
    LocalMux I__8741 (
            .O(N__40332),
            .I(N__40309));
    Span4Mux_h I__8740 (
            .O(N__40329),
            .I(N__40306));
    Span4Mux_h I__8739 (
            .O(N__40324),
            .I(N__40301));
    Span4Mux_v I__8738 (
            .O(N__40317),
            .I(N__40301));
    Span12Mux_v I__8737 (
            .O(N__40312),
            .I(N__40296));
    Span4Mux_h I__8736 (
            .O(N__40309),
            .I(N__40291));
    Span4Mux_h I__8735 (
            .O(N__40306),
            .I(N__40291));
    Span4Mux_v I__8734 (
            .O(N__40301),
            .I(N__40288));
    InMux I__8733 (
            .O(N__40300),
            .I(N__40283));
    InMux I__8732 (
            .O(N__40299),
            .I(N__40283));
    Odrv12 I__8731 (
            .O(N__40296),
            .I(uart_pc_data_4));
    Odrv4 I__8730 (
            .O(N__40291),
            .I(uart_pc_data_4));
    Odrv4 I__8729 (
            .O(N__40288),
            .I(uart_pc_data_4));
    LocalMux I__8728 (
            .O(N__40283),
            .I(uart_pc_data_4));
    InMux I__8727 (
            .O(N__40274),
            .I(N__40269));
    InMux I__8726 (
            .O(N__40273),
            .I(N__40266));
    InMux I__8725 (
            .O(N__40272),
            .I(N__40263));
    LocalMux I__8724 (
            .O(N__40269),
            .I(N__40258));
    LocalMux I__8723 (
            .O(N__40266),
            .I(N__40251));
    LocalMux I__8722 (
            .O(N__40263),
            .I(N__40247));
    InMux I__8721 (
            .O(N__40262),
            .I(N__40243));
    InMux I__8720 (
            .O(N__40261),
            .I(N__40240));
    Span4Mux_h I__8719 (
            .O(N__40258),
            .I(N__40235));
    InMux I__8718 (
            .O(N__40257),
            .I(N__40232));
    InMux I__8717 (
            .O(N__40256),
            .I(N__40229));
    InMux I__8716 (
            .O(N__40255),
            .I(N__40226));
    InMux I__8715 (
            .O(N__40254),
            .I(N__40223));
    Span4Mux_h I__8714 (
            .O(N__40251),
            .I(N__40220));
    InMux I__8713 (
            .O(N__40250),
            .I(N__40217));
    Span4Mux_v I__8712 (
            .O(N__40247),
            .I(N__40214));
    InMux I__8711 (
            .O(N__40246),
            .I(N__40211));
    LocalMux I__8710 (
            .O(N__40243),
            .I(N__40208));
    LocalMux I__8709 (
            .O(N__40240),
            .I(N__40205));
    InMux I__8708 (
            .O(N__40239),
            .I(N__40200));
    InMux I__8707 (
            .O(N__40238),
            .I(N__40200));
    Span4Mux_v I__8706 (
            .O(N__40235),
            .I(N__40195));
    LocalMux I__8705 (
            .O(N__40232),
            .I(N__40195));
    LocalMux I__8704 (
            .O(N__40229),
            .I(N__40189));
    LocalMux I__8703 (
            .O(N__40226),
            .I(N__40189));
    LocalMux I__8702 (
            .O(N__40223),
            .I(N__40184));
    Span4Mux_h I__8701 (
            .O(N__40220),
            .I(N__40184));
    LocalMux I__8700 (
            .O(N__40217),
            .I(N__40179));
    Sp12to4 I__8699 (
            .O(N__40214),
            .I(N__40179));
    LocalMux I__8698 (
            .O(N__40211),
            .I(N__40170));
    Span4Mux_h I__8697 (
            .O(N__40208),
            .I(N__40170));
    Span4Mux_v I__8696 (
            .O(N__40205),
            .I(N__40170));
    LocalMux I__8695 (
            .O(N__40200),
            .I(N__40170));
    Span4Mux_v I__8694 (
            .O(N__40195),
            .I(N__40167));
    InMux I__8693 (
            .O(N__40194),
            .I(N__40164));
    Span12Mux_v I__8692 (
            .O(N__40189),
            .I(N__40161));
    Sp12to4 I__8691 (
            .O(N__40184),
            .I(N__40156));
    Span12Mux_s8_h I__8690 (
            .O(N__40179),
            .I(N__40156));
    Span4Mux_h I__8689 (
            .O(N__40170),
            .I(N__40151));
    Span4Mux_h I__8688 (
            .O(N__40167),
            .I(N__40151));
    LocalMux I__8687 (
            .O(N__40164),
            .I(uart_pc_data_5));
    Odrv12 I__8686 (
            .O(N__40161),
            .I(uart_pc_data_5));
    Odrv12 I__8685 (
            .O(N__40156),
            .I(uart_pc_data_5));
    Odrv4 I__8684 (
            .O(N__40151),
            .I(uart_pc_data_5));
    InMux I__8683 (
            .O(N__40142),
            .I(N__40135));
    InMux I__8682 (
            .O(N__40141),
            .I(N__40132));
    InMux I__8681 (
            .O(N__40140),
            .I(N__40129));
    InMux I__8680 (
            .O(N__40139),
            .I(N__40126));
    InMux I__8679 (
            .O(N__40138),
            .I(N__40123));
    LocalMux I__8678 (
            .O(N__40135),
            .I(N__40116));
    LocalMux I__8677 (
            .O(N__40132),
            .I(N__40116));
    LocalMux I__8676 (
            .O(N__40129),
            .I(N__40111));
    LocalMux I__8675 (
            .O(N__40126),
            .I(N__40111));
    LocalMux I__8674 (
            .O(N__40123),
            .I(N__40107));
    InMux I__8673 (
            .O(N__40122),
            .I(N__40103));
    InMux I__8672 (
            .O(N__40121),
            .I(N__40100));
    Span4Mux_v I__8671 (
            .O(N__40116),
            .I(N__40097));
    Span4Mux_v I__8670 (
            .O(N__40111),
            .I(N__40094));
    InMux I__8669 (
            .O(N__40110),
            .I(N__40090));
    Span4Mux_h I__8668 (
            .O(N__40107),
            .I(N__40087));
    InMux I__8667 (
            .O(N__40106),
            .I(N__40084));
    LocalMux I__8666 (
            .O(N__40103),
            .I(N__40081));
    LocalMux I__8665 (
            .O(N__40100),
            .I(N__40078));
    Sp12to4 I__8664 (
            .O(N__40097),
            .I(N__40075));
    Sp12to4 I__8663 (
            .O(N__40094),
            .I(N__40072));
    InMux I__8662 (
            .O(N__40093),
            .I(N__40069));
    LocalMux I__8661 (
            .O(N__40090),
            .I(N__40066));
    Span4Mux_h I__8660 (
            .O(N__40087),
            .I(N__40063));
    LocalMux I__8659 (
            .O(N__40084),
            .I(N__40060));
    Span4Mux_v I__8658 (
            .O(N__40081),
            .I(N__40057));
    Span12Mux_s10_v I__8657 (
            .O(N__40078),
            .I(N__40048));
    Span12Mux_s5_h I__8656 (
            .O(N__40075),
            .I(N__40048));
    Span12Mux_h I__8655 (
            .O(N__40072),
            .I(N__40048));
    LocalMux I__8654 (
            .O(N__40069),
            .I(N__40048));
    Span4Mux_h I__8653 (
            .O(N__40066),
            .I(N__40045));
    Span4Mux_v I__8652 (
            .O(N__40063),
            .I(N__40042));
    Span4Mux_h I__8651 (
            .O(N__40060),
            .I(N__40037));
    Sp12to4 I__8650 (
            .O(N__40057),
            .I(N__40032));
    Span12Mux_v I__8649 (
            .O(N__40048),
            .I(N__40032));
    Span4Mux_h I__8648 (
            .O(N__40045),
            .I(N__40027));
    Span4Mux_v I__8647 (
            .O(N__40042),
            .I(N__40027));
    InMux I__8646 (
            .O(N__40041),
            .I(N__40022));
    InMux I__8645 (
            .O(N__40040),
            .I(N__40022));
    Odrv4 I__8644 (
            .O(N__40037),
            .I(uart_pc_data_6));
    Odrv12 I__8643 (
            .O(N__40032),
            .I(uart_pc_data_6));
    Odrv4 I__8642 (
            .O(N__40027),
            .I(uart_pc_data_6));
    LocalMux I__8641 (
            .O(N__40022),
            .I(uart_pc_data_6));
    InMux I__8640 (
            .O(N__40013),
            .I(N__40007));
    InMux I__8639 (
            .O(N__40012),
            .I(N__40002));
    InMux I__8638 (
            .O(N__40011),
            .I(N__39998));
    InMux I__8637 (
            .O(N__40010),
            .I(N__39995));
    LocalMux I__8636 (
            .O(N__40007),
            .I(N__39990));
    InMux I__8635 (
            .O(N__40006),
            .I(N__39987));
    InMux I__8634 (
            .O(N__40005),
            .I(N__39984));
    LocalMux I__8633 (
            .O(N__40002),
            .I(N__39979));
    InMux I__8632 (
            .O(N__40001),
            .I(N__39976));
    LocalMux I__8631 (
            .O(N__39998),
            .I(N__39969));
    LocalMux I__8630 (
            .O(N__39995),
            .I(N__39969));
    InMux I__8629 (
            .O(N__39994),
            .I(N__39966));
    InMux I__8628 (
            .O(N__39993),
            .I(N__39963));
    Span4Mux_v I__8627 (
            .O(N__39990),
            .I(N__39960));
    LocalMux I__8626 (
            .O(N__39987),
            .I(N__39955));
    LocalMux I__8625 (
            .O(N__39984),
            .I(N__39955));
    InMux I__8624 (
            .O(N__39983),
            .I(N__39952));
    InMux I__8623 (
            .O(N__39982),
            .I(N__39949));
    Span4Mux_h I__8622 (
            .O(N__39979),
            .I(N__39944));
    LocalMux I__8621 (
            .O(N__39976),
            .I(N__39944));
    InMux I__8620 (
            .O(N__39975),
            .I(N__39939));
    InMux I__8619 (
            .O(N__39974),
            .I(N__39939));
    Span4Mux_v I__8618 (
            .O(N__39969),
            .I(N__39934));
    LocalMux I__8617 (
            .O(N__39966),
            .I(N__39934));
    LocalMux I__8616 (
            .O(N__39963),
            .I(N__39931));
    Span4Mux_h I__8615 (
            .O(N__39960),
            .I(N__39925));
    Span4Mux_v I__8614 (
            .O(N__39955),
            .I(N__39925));
    LocalMux I__8613 (
            .O(N__39952),
            .I(N__39918));
    LocalMux I__8612 (
            .O(N__39949),
            .I(N__39918));
    Span4Mux_v I__8611 (
            .O(N__39944),
            .I(N__39918));
    LocalMux I__8610 (
            .O(N__39939),
            .I(N__39915));
    Span4Mux_v I__8609 (
            .O(N__39934),
            .I(N__39912));
    Span12Mux_h I__8608 (
            .O(N__39931),
            .I(N__39909));
    InMux I__8607 (
            .O(N__39930),
            .I(N__39906));
    Span4Mux_v I__8606 (
            .O(N__39925),
            .I(N__39901));
    Span4Mux_h I__8605 (
            .O(N__39918),
            .I(N__39901));
    Span4Mux_h I__8604 (
            .O(N__39915),
            .I(N__39898));
    Span4Mux_h I__8603 (
            .O(N__39912),
            .I(N__39895));
    Odrv12 I__8602 (
            .O(N__39909),
            .I(uart_pc_data_7));
    LocalMux I__8601 (
            .O(N__39906),
            .I(uart_pc_data_7));
    Odrv4 I__8600 (
            .O(N__39901),
            .I(uart_pc_data_7));
    Odrv4 I__8599 (
            .O(N__39898),
            .I(uart_pc_data_7));
    Odrv4 I__8598 (
            .O(N__39895),
            .I(uart_pc_data_7));
    CEMux I__8597 (
            .O(N__39884),
            .I(N__39881));
    LocalMux I__8596 (
            .O(N__39881),
            .I(N__39878));
    Span4Mux_v I__8595 (
            .O(N__39878),
            .I(N__39875));
    Sp12to4 I__8594 (
            .O(N__39875),
            .I(N__39872));
    Span12Mux_h I__8593 (
            .O(N__39872),
            .I(N__39869));
    Odrv12 I__8592 (
            .O(N__39869),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ));
    InMux I__8591 (
            .O(N__39866),
            .I(N__39863));
    LocalMux I__8590 (
            .O(N__39863),
            .I(\dron_frame_decoder_1.drone_H_disp_front_10 ));
    InMux I__8589 (
            .O(N__39860),
            .I(N__39857));
    LocalMux I__8588 (
            .O(N__39857),
            .I(\dron_frame_decoder_1.drone_H_disp_front_9 ));
    InMux I__8587 (
            .O(N__39854),
            .I(N__39848));
    InMux I__8586 (
            .O(N__39853),
            .I(N__39848));
    LocalMux I__8585 (
            .O(N__39848),
            .I(front_command_7));
    InMux I__8584 (
            .O(N__39845),
            .I(N__39839));
    InMux I__8583 (
            .O(N__39844),
            .I(N__39839));
    LocalMux I__8582 (
            .O(N__39839),
            .I(drone_H_disp_front_11));
    InMux I__8581 (
            .O(N__39836),
            .I(N__39833));
    LocalMux I__8580 (
            .O(N__39833),
            .I(N__39830));
    Span4Mux_h I__8579 (
            .O(N__39830),
            .I(N__39827));
    Span4Mux_h I__8578 (
            .O(N__39827),
            .I(N__39824));
    Odrv4 I__8577 (
            .O(N__39824),
            .I(\uart_pc.data_Auxce_0_6 ));
    CascadeMux I__8576 (
            .O(N__39821),
            .I(N__39818));
    InMux I__8575 (
            .O(N__39818),
            .I(N__39815));
    LocalMux I__8574 (
            .O(N__39815),
            .I(N__39812));
    Span4Mux_h I__8573 (
            .O(N__39812),
            .I(N__39808));
    CascadeMux I__8572 (
            .O(N__39811),
            .I(N__39805));
    Span4Mux_h I__8571 (
            .O(N__39808),
            .I(N__39802));
    InMux I__8570 (
            .O(N__39805),
            .I(N__39799));
    Odrv4 I__8569 (
            .O(N__39802),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    LocalMux I__8568 (
            .O(N__39799),
            .I(\uart_pc.data_AuxZ0Z_6 ));
    InMux I__8567 (
            .O(N__39794),
            .I(N__39791));
    LocalMux I__8566 (
            .O(N__39791),
            .I(\dron_frame_decoder_1.drone_H_disp_front_4 ));
    InMux I__8565 (
            .O(N__39788),
            .I(N__39785));
    LocalMux I__8564 (
            .O(N__39785),
            .I(\dron_frame_decoder_1.drone_H_disp_front_5 ));
    InMux I__8563 (
            .O(N__39782),
            .I(N__39779));
    LocalMux I__8562 (
            .O(N__39779),
            .I(\dron_frame_decoder_1.drone_H_disp_front_6 ));
    InMux I__8561 (
            .O(N__39776),
            .I(N__39773));
    LocalMux I__8560 (
            .O(N__39773),
            .I(\dron_frame_decoder_1.drone_H_disp_front_7 ));
    InMux I__8559 (
            .O(N__39770),
            .I(N__39765));
    InMux I__8558 (
            .O(N__39769),
            .I(N__39762));
    InMux I__8557 (
            .O(N__39768),
            .I(N__39756));
    LocalMux I__8556 (
            .O(N__39765),
            .I(N__39750));
    LocalMux I__8555 (
            .O(N__39762),
            .I(N__39746));
    InMux I__8554 (
            .O(N__39761),
            .I(N__39743));
    InMux I__8553 (
            .O(N__39760),
            .I(N__39739));
    InMux I__8552 (
            .O(N__39759),
            .I(N__39736));
    LocalMux I__8551 (
            .O(N__39756),
            .I(N__39733));
    InMux I__8550 (
            .O(N__39755),
            .I(N__39730));
    InMux I__8549 (
            .O(N__39754),
            .I(N__39727));
    InMux I__8548 (
            .O(N__39753),
            .I(N__39724));
    Span4Mux_v I__8547 (
            .O(N__39750),
            .I(N__39721));
    InMux I__8546 (
            .O(N__39749),
            .I(N__39718));
    Span4Mux_v I__8545 (
            .O(N__39746),
            .I(N__39713));
    LocalMux I__8544 (
            .O(N__39743),
            .I(N__39713));
    InMux I__8543 (
            .O(N__39742),
            .I(N__39710));
    LocalMux I__8542 (
            .O(N__39739),
            .I(N__39707));
    LocalMux I__8541 (
            .O(N__39736),
            .I(N__39699));
    Sp12to4 I__8540 (
            .O(N__39733),
            .I(N__39699));
    LocalMux I__8539 (
            .O(N__39730),
            .I(N__39699));
    LocalMux I__8538 (
            .O(N__39727),
            .I(N__39692));
    LocalMux I__8537 (
            .O(N__39724),
            .I(N__39692));
    Span4Mux_v I__8536 (
            .O(N__39721),
            .I(N__39683));
    LocalMux I__8535 (
            .O(N__39718),
            .I(N__39683));
    Span4Mux_h I__8534 (
            .O(N__39713),
            .I(N__39683));
    LocalMux I__8533 (
            .O(N__39710),
            .I(N__39683));
    Span12Mux_v I__8532 (
            .O(N__39707),
            .I(N__39680));
    InMux I__8531 (
            .O(N__39706),
            .I(N__39677));
    Span12Mux_v I__8530 (
            .O(N__39699),
            .I(N__39674));
    InMux I__8529 (
            .O(N__39698),
            .I(N__39669));
    InMux I__8528 (
            .O(N__39697),
            .I(N__39669));
    Span4Mux_v I__8527 (
            .O(N__39692),
            .I(N__39664));
    Span4Mux_v I__8526 (
            .O(N__39683),
            .I(N__39664));
    Odrv12 I__8525 (
            .O(N__39680),
            .I(uart_pc_data_0));
    LocalMux I__8524 (
            .O(N__39677),
            .I(uart_pc_data_0));
    Odrv12 I__8523 (
            .O(N__39674),
            .I(uart_pc_data_0));
    LocalMux I__8522 (
            .O(N__39669),
            .I(uart_pc_data_0));
    Odrv4 I__8521 (
            .O(N__39664),
            .I(uart_pc_data_0));
    InMux I__8520 (
            .O(N__39653),
            .I(N__39648));
    InMux I__8519 (
            .O(N__39652),
            .I(N__39645));
    InMux I__8518 (
            .O(N__39651),
            .I(N__39642));
    LocalMux I__8517 (
            .O(N__39648),
            .I(N__39638));
    LocalMux I__8516 (
            .O(N__39645),
            .I(N__39635));
    LocalMux I__8515 (
            .O(N__39642),
            .I(N__39630));
    InMux I__8514 (
            .O(N__39641),
            .I(N__39627));
    Span4Mux_h I__8513 (
            .O(N__39638),
            .I(N__39620));
    Span4Mux_v I__8512 (
            .O(N__39635),
            .I(N__39620));
    InMux I__8511 (
            .O(N__39634),
            .I(N__39615));
    InMux I__8510 (
            .O(N__39633),
            .I(N__39615));
    Span4Mux_v I__8509 (
            .O(N__39630),
            .I(N__39612));
    LocalMux I__8508 (
            .O(N__39627),
            .I(N__39609));
    InMux I__8507 (
            .O(N__39626),
            .I(N__39606));
    InMux I__8506 (
            .O(N__39625),
            .I(N__39603));
    Span4Mux_v I__8505 (
            .O(N__39620),
            .I(N__39598));
    LocalMux I__8504 (
            .O(N__39615),
            .I(N__39598));
    Span4Mux_v I__8503 (
            .O(N__39612),
            .I(N__39595));
    Span4Mux_v I__8502 (
            .O(N__39609),
            .I(N__39591));
    LocalMux I__8501 (
            .O(N__39606),
            .I(N__39588));
    LocalMux I__8500 (
            .O(N__39603),
            .I(N__39585));
    Span4Mux_v I__8499 (
            .O(N__39598),
            .I(N__39582));
    Sp12to4 I__8498 (
            .O(N__39595),
            .I(N__39578));
    InMux I__8497 (
            .O(N__39594),
            .I(N__39573));
    Span4Mux_v I__8496 (
            .O(N__39591),
            .I(N__39570));
    Span4Mux_v I__8495 (
            .O(N__39588),
            .I(N__39565));
    Span4Mux_s3_h I__8494 (
            .O(N__39585),
            .I(N__39565));
    Span4Mux_h I__8493 (
            .O(N__39582),
            .I(N__39562));
    InMux I__8492 (
            .O(N__39581),
            .I(N__39559));
    Span12Mux_h I__8491 (
            .O(N__39578),
            .I(N__39556));
    InMux I__8490 (
            .O(N__39577),
            .I(N__39553));
    InMux I__8489 (
            .O(N__39576),
            .I(N__39550));
    LocalMux I__8488 (
            .O(N__39573),
            .I(N__39541));
    Span4Mux_v I__8487 (
            .O(N__39570),
            .I(N__39541));
    Span4Mux_h I__8486 (
            .O(N__39565),
            .I(N__39541));
    Span4Mux_v I__8485 (
            .O(N__39562),
            .I(N__39541));
    LocalMux I__8484 (
            .O(N__39559),
            .I(N__39538));
    Odrv12 I__8483 (
            .O(N__39556),
            .I(uart_pc_data_1));
    LocalMux I__8482 (
            .O(N__39553),
            .I(uart_pc_data_1));
    LocalMux I__8481 (
            .O(N__39550),
            .I(uart_pc_data_1));
    Odrv4 I__8480 (
            .O(N__39541),
            .I(uart_pc_data_1));
    Odrv4 I__8479 (
            .O(N__39538),
            .I(uart_pc_data_1));
    InMux I__8478 (
            .O(N__39527),
            .I(N__39522));
    InMux I__8477 (
            .O(N__39526),
            .I(N__39519));
    InMux I__8476 (
            .O(N__39525),
            .I(N__39516));
    LocalMux I__8475 (
            .O(N__39522),
            .I(N__39513));
    LocalMux I__8474 (
            .O(N__39519),
            .I(N__39509));
    LocalMux I__8473 (
            .O(N__39516),
            .I(N__39504));
    Span4Mux_v I__8472 (
            .O(N__39513),
            .I(N__39504));
    InMux I__8471 (
            .O(N__39512),
            .I(N__39501));
    Span4Mux_v I__8470 (
            .O(N__39509),
            .I(N__39492));
    Span4Mux_h I__8469 (
            .O(N__39504),
            .I(N__39492));
    LocalMux I__8468 (
            .O(N__39501),
            .I(N__39489));
    InMux I__8467 (
            .O(N__39500),
            .I(N__39484));
    InMux I__8466 (
            .O(N__39499),
            .I(N__39478));
    InMux I__8465 (
            .O(N__39498),
            .I(N__39478));
    CascadeMux I__8464 (
            .O(N__39497),
            .I(N__39475));
    Span4Mux_v I__8463 (
            .O(N__39492),
            .I(N__39471));
    Sp12to4 I__8462 (
            .O(N__39489),
            .I(N__39468));
    InMux I__8461 (
            .O(N__39488),
            .I(N__39463));
    InMux I__8460 (
            .O(N__39487),
            .I(N__39460));
    LocalMux I__8459 (
            .O(N__39484),
            .I(N__39457));
    InMux I__8458 (
            .O(N__39483),
            .I(N__39454));
    LocalMux I__8457 (
            .O(N__39478),
            .I(N__39451));
    InMux I__8456 (
            .O(N__39475),
            .I(N__39448));
    CascadeMux I__8455 (
            .O(N__39474),
            .I(N__39445));
    Sp12to4 I__8454 (
            .O(N__39471),
            .I(N__39440));
    Span12Mux_v I__8453 (
            .O(N__39468),
            .I(N__39440));
    CascadeMux I__8452 (
            .O(N__39467),
            .I(N__39436));
    InMux I__8451 (
            .O(N__39466),
            .I(N__39433));
    LocalMux I__8450 (
            .O(N__39463),
            .I(N__39430));
    LocalMux I__8449 (
            .O(N__39460),
            .I(N__39427));
    Span4Mux_h I__8448 (
            .O(N__39457),
            .I(N__39422));
    LocalMux I__8447 (
            .O(N__39454),
            .I(N__39422));
    Span4Mux_v I__8446 (
            .O(N__39451),
            .I(N__39419));
    LocalMux I__8445 (
            .O(N__39448),
            .I(N__39416));
    InMux I__8444 (
            .O(N__39445),
            .I(N__39413));
    Span12Mux_h I__8443 (
            .O(N__39440),
            .I(N__39410));
    InMux I__8442 (
            .O(N__39439),
            .I(N__39405));
    InMux I__8441 (
            .O(N__39436),
            .I(N__39405));
    LocalMux I__8440 (
            .O(N__39433),
            .I(N__39394));
    Span4Mux_h I__8439 (
            .O(N__39430),
            .I(N__39394));
    Span4Mux_v I__8438 (
            .O(N__39427),
            .I(N__39394));
    Span4Mux_v I__8437 (
            .O(N__39422),
            .I(N__39394));
    Span4Mux_v I__8436 (
            .O(N__39419),
            .I(N__39394));
    Span4Mux_h I__8435 (
            .O(N__39416),
            .I(N__39391));
    LocalMux I__8434 (
            .O(N__39413),
            .I(uart_pc_data_2));
    Odrv12 I__8433 (
            .O(N__39410),
            .I(uart_pc_data_2));
    LocalMux I__8432 (
            .O(N__39405),
            .I(uart_pc_data_2));
    Odrv4 I__8431 (
            .O(N__39394),
            .I(uart_pc_data_2));
    Odrv4 I__8430 (
            .O(N__39391),
            .I(uart_pc_data_2));
    InMux I__8429 (
            .O(N__39380),
            .I(N__39377));
    LocalMux I__8428 (
            .O(N__39377),
            .I(N__39374));
    Span4Mux_v I__8427 (
            .O(N__39374),
            .I(N__39370));
    InMux I__8426 (
            .O(N__39373),
            .I(N__39367));
    Span4Mux_h I__8425 (
            .O(N__39370),
            .I(N__39359));
    LocalMux I__8424 (
            .O(N__39367),
            .I(N__39356));
    InMux I__8423 (
            .O(N__39366),
            .I(N__39353));
    InMux I__8422 (
            .O(N__39365),
            .I(N__39348));
    InMux I__8421 (
            .O(N__39364),
            .I(N__39348));
    InMux I__8420 (
            .O(N__39363),
            .I(N__39345));
    InMux I__8419 (
            .O(N__39362),
            .I(N__39340));
    Span4Mux_h I__8418 (
            .O(N__39359),
            .I(N__39335));
    Span4Mux_v I__8417 (
            .O(N__39356),
            .I(N__39335));
    LocalMux I__8416 (
            .O(N__39353),
            .I(N__39331));
    LocalMux I__8415 (
            .O(N__39348),
            .I(N__39328));
    LocalMux I__8414 (
            .O(N__39345),
            .I(N__39325));
    InMux I__8413 (
            .O(N__39344),
            .I(N__39322));
    InMux I__8412 (
            .O(N__39343),
            .I(N__39319));
    LocalMux I__8411 (
            .O(N__39340),
            .I(N__39316));
    Span4Mux_v I__8410 (
            .O(N__39335),
            .I(N__39313));
    InMux I__8409 (
            .O(N__39334),
            .I(N__39310));
    Span4Mux_v I__8408 (
            .O(N__39331),
            .I(N__39305));
    Span4Mux_h I__8407 (
            .O(N__39328),
            .I(N__39305));
    Span12Mux_s10_v I__8406 (
            .O(N__39325),
            .I(N__39302));
    LocalMux I__8405 (
            .O(N__39322),
            .I(N__39299));
    LocalMux I__8404 (
            .O(N__39319),
            .I(N__39294));
    Span4Mux_h I__8403 (
            .O(N__39316),
            .I(N__39294));
    Sp12to4 I__8402 (
            .O(N__39313),
            .I(N__39291));
    LocalMux I__8401 (
            .O(N__39310),
            .I(N__39288));
    Span4Mux_h I__8400 (
            .O(N__39305),
            .I(N__39285));
    Span12Mux_v I__8399 (
            .O(N__39302),
            .I(N__39280));
    Span4Mux_h I__8398 (
            .O(N__39299),
            .I(N__39277));
    Span4Mux_h I__8397 (
            .O(N__39294),
            .I(N__39274));
    Span12Mux_h I__8396 (
            .O(N__39291),
            .I(N__39267));
    Span12Mux_s9_h I__8395 (
            .O(N__39288),
            .I(N__39267));
    Sp12to4 I__8394 (
            .O(N__39285),
            .I(N__39267));
    InMux I__8393 (
            .O(N__39284),
            .I(N__39262));
    InMux I__8392 (
            .O(N__39283),
            .I(N__39262));
    Odrv12 I__8391 (
            .O(N__39280),
            .I(uart_pc_data_3));
    Odrv4 I__8390 (
            .O(N__39277),
            .I(uart_pc_data_3));
    Odrv4 I__8389 (
            .O(N__39274),
            .I(uart_pc_data_3));
    Odrv12 I__8388 (
            .O(N__39267),
            .I(uart_pc_data_3));
    LocalMux I__8387 (
            .O(N__39262),
            .I(uart_pc_data_3));
    InMux I__8386 (
            .O(N__39251),
            .I(N__39247));
    CascadeMux I__8385 (
            .O(N__39250),
            .I(N__39243));
    LocalMux I__8384 (
            .O(N__39247),
            .I(N__39240));
    InMux I__8383 (
            .O(N__39246),
            .I(N__39237));
    InMux I__8382 (
            .O(N__39243),
            .I(N__39234));
    Span4Mux_h I__8381 (
            .O(N__39240),
            .I(N__39231));
    LocalMux I__8380 (
            .O(N__39237),
            .I(N__39228));
    LocalMux I__8379 (
            .O(N__39234),
            .I(front_order_2));
    Odrv4 I__8378 (
            .O(N__39231),
            .I(front_order_2));
    Odrv4 I__8377 (
            .O(N__39228),
            .I(front_order_2));
    InMux I__8376 (
            .O(N__39221),
            .I(N__39218));
    LocalMux I__8375 (
            .O(N__39218),
            .I(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ));
    CascadeMux I__8374 (
            .O(N__39215),
            .I(N__39211));
    InMux I__8373 (
            .O(N__39214),
            .I(N__39208));
    InMux I__8372 (
            .O(N__39211),
            .I(N__39204));
    LocalMux I__8371 (
            .O(N__39208),
            .I(N__39201));
    InMux I__8370 (
            .O(N__39207),
            .I(N__39198));
    LocalMux I__8369 (
            .O(N__39204),
            .I(N__39193));
    Span4Mux_h I__8368 (
            .O(N__39201),
            .I(N__39193));
    LocalMux I__8367 (
            .O(N__39198),
            .I(N__39190));
    Odrv4 I__8366 (
            .O(N__39193),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    Odrv12 I__8365 (
            .O(N__39190),
            .I(\ppm_encoder_1.elevatorZ0Z_2 ));
    InMux I__8364 (
            .O(N__39185),
            .I(N__39182));
    LocalMux I__8363 (
            .O(N__39182),
            .I(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ));
    CascadeMux I__8362 (
            .O(N__39179),
            .I(N__39176));
    InMux I__8361 (
            .O(N__39176),
            .I(N__39173));
    LocalMux I__8360 (
            .O(N__39173),
            .I(N__39168));
    InMux I__8359 (
            .O(N__39172),
            .I(N__39165));
    InMux I__8358 (
            .O(N__39171),
            .I(N__39162));
    Span4Mux_h I__8357 (
            .O(N__39168),
            .I(N__39157));
    LocalMux I__8356 (
            .O(N__39165),
            .I(N__39157));
    LocalMux I__8355 (
            .O(N__39162),
            .I(front_order_6));
    Odrv4 I__8354 (
            .O(N__39157),
            .I(front_order_6));
    InMux I__8353 (
            .O(N__39152),
            .I(N__39149));
    LocalMux I__8352 (
            .O(N__39149),
            .I(N__39145));
    InMux I__8351 (
            .O(N__39148),
            .I(N__39141));
    Span4Mux_h I__8350 (
            .O(N__39145),
            .I(N__39138));
    InMux I__8349 (
            .O(N__39144),
            .I(N__39135));
    LocalMux I__8348 (
            .O(N__39141),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    Odrv4 I__8347 (
            .O(N__39138),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    LocalMux I__8346 (
            .O(N__39135),
            .I(\ppm_encoder_1.elevatorZ0Z_6 ));
    InMux I__8345 (
            .O(N__39128),
            .I(N__39124));
    InMux I__8344 (
            .O(N__39127),
            .I(N__39121));
    LocalMux I__8343 (
            .O(N__39124),
            .I(N__39118));
    LocalMux I__8342 (
            .O(N__39121),
            .I(N__39115));
    Span4Mux_v I__8341 (
            .O(N__39118),
            .I(N__39112));
    Span4Mux_v I__8340 (
            .O(N__39115),
            .I(N__39109));
    Odrv4 I__8339 (
            .O(N__39112),
            .I(front_order_5));
    Odrv4 I__8338 (
            .O(N__39109),
            .I(front_order_5));
    InMux I__8337 (
            .O(N__39104),
            .I(N__39101));
    LocalMux I__8336 (
            .O(N__39101),
            .I(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ));
    InMux I__8335 (
            .O(N__39098),
            .I(N__39094));
    CascadeMux I__8334 (
            .O(N__39097),
            .I(N__39091));
    LocalMux I__8333 (
            .O(N__39094),
            .I(N__39088));
    InMux I__8332 (
            .O(N__39091),
            .I(N__39084));
    Span4Mux_h I__8331 (
            .O(N__39088),
            .I(N__39081));
    InMux I__8330 (
            .O(N__39087),
            .I(N__39078));
    LocalMux I__8329 (
            .O(N__39084),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    Odrv4 I__8328 (
            .O(N__39081),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    LocalMux I__8327 (
            .O(N__39078),
            .I(\ppm_encoder_1.elevatorZ0Z_5 ));
    InMux I__8326 (
            .O(N__39071),
            .I(N__39068));
    LocalMux I__8325 (
            .O(N__39068),
            .I(N__39064));
    InMux I__8324 (
            .O(N__39067),
            .I(N__39061));
    Span4Mux_v I__8323 (
            .O(N__39064),
            .I(N__39058));
    LocalMux I__8322 (
            .O(N__39061),
            .I(N__39055));
    Span4Mux_h I__8321 (
            .O(N__39058),
            .I(N__39052));
    Span4Mux_v I__8320 (
            .O(N__39055),
            .I(N__39049));
    Span4Mux_h I__8319 (
            .O(N__39052),
            .I(N__39046));
    Span4Mux_h I__8318 (
            .O(N__39049),
            .I(N__39043));
    Span4Mux_h I__8317 (
            .O(N__39046),
            .I(N__39040));
    Span4Mux_h I__8316 (
            .O(N__39043),
            .I(N__39037));
    Odrv4 I__8315 (
            .O(N__39040),
            .I(xy_kp_5));
    Odrv4 I__8314 (
            .O(N__39037),
            .I(xy_kp_5));
    CEMux I__8313 (
            .O(N__39032),
            .I(N__39028));
    CEMux I__8312 (
            .O(N__39031),
            .I(N__39023));
    LocalMux I__8311 (
            .O(N__39028),
            .I(N__39020));
    CEMux I__8310 (
            .O(N__39027),
            .I(N__39017));
    CEMux I__8309 (
            .O(N__39026),
            .I(N__39014));
    LocalMux I__8308 (
            .O(N__39023),
            .I(N__39011));
    Span4Mux_v I__8307 (
            .O(N__39020),
            .I(N__39008));
    LocalMux I__8306 (
            .O(N__39017),
            .I(N__39005));
    LocalMux I__8305 (
            .O(N__39014),
            .I(N__39002));
    Span4Mux_h I__8304 (
            .O(N__39011),
            .I(N__38999));
    Span4Mux_h I__8303 (
            .O(N__39008),
            .I(N__38994));
    Span4Mux_v I__8302 (
            .O(N__39005),
            .I(N__38994));
    Span4Mux_h I__8301 (
            .O(N__39002),
            .I(N__38991));
    Span4Mux_v I__8300 (
            .O(N__38999),
            .I(N__38988));
    Span4Mux_h I__8299 (
            .O(N__38994),
            .I(N__38985));
    Span4Mux_v I__8298 (
            .O(N__38991),
            .I(N__38982));
    Odrv4 I__8297 (
            .O(N__38988),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    Odrv4 I__8296 (
            .O(N__38985),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    Odrv4 I__8295 (
            .O(N__38982),
            .I(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ));
    CascadeMux I__8294 (
            .O(N__38975),
            .I(N__38970));
    InMux I__8293 (
            .O(N__38974),
            .I(N__38967));
    InMux I__8292 (
            .O(N__38973),
            .I(N__38962));
    InMux I__8291 (
            .O(N__38970),
            .I(N__38962));
    LocalMux I__8290 (
            .O(N__38967),
            .I(N__38956));
    LocalMux I__8289 (
            .O(N__38962),
            .I(N__38956));
    InMux I__8288 (
            .O(N__38961),
            .I(N__38952));
    Span4Mux_h I__8287 (
            .O(N__38956),
            .I(N__38949));
    InMux I__8286 (
            .O(N__38955),
            .I(N__38946));
    LocalMux I__8285 (
            .O(N__38952),
            .I(\pid_front.pid_preregZ0Z_4 ));
    Odrv4 I__8284 (
            .O(N__38949),
            .I(\pid_front.pid_preregZ0Z_4 ));
    LocalMux I__8283 (
            .O(N__38946),
            .I(\pid_front.pid_preregZ0Z_4 ));
    InMux I__8282 (
            .O(N__38939),
            .I(N__38931));
    InMux I__8281 (
            .O(N__38938),
            .I(N__38931));
    InMux I__8280 (
            .O(N__38937),
            .I(N__38926));
    InMux I__8279 (
            .O(N__38936),
            .I(N__38926));
    LocalMux I__8278 (
            .O(N__38931),
            .I(N__38919));
    LocalMux I__8277 (
            .O(N__38926),
            .I(N__38919));
    CascadeMux I__8276 (
            .O(N__38925),
            .I(N__38916));
    InMux I__8275 (
            .O(N__38924),
            .I(N__38913));
    Span4Mux_h I__8274 (
            .O(N__38919),
            .I(N__38910));
    InMux I__8273 (
            .O(N__38916),
            .I(N__38907));
    LocalMux I__8272 (
            .O(N__38913),
            .I(\pid_front.pid_preregZ0Z_5 ));
    Odrv4 I__8271 (
            .O(N__38910),
            .I(\pid_front.pid_preregZ0Z_5 ));
    LocalMux I__8270 (
            .O(N__38907),
            .I(\pid_front.pid_preregZ0Z_5 ));
    InMux I__8269 (
            .O(N__38900),
            .I(N__38896));
    InMux I__8268 (
            .O(N__38899),
            .I(N__38893));
    LocalMux I__8267 (
            .O(N__38896),
            .I(N__38887));
    LocalMux I__8266 (
            .O(N__38893),
            .I(N__38887));
    InMux I__8265 (
            .O(N__38892),
            .I(N__38883));
    Span4Mux_v I__8264 (
            .O(N__38887),
            .I(N__38880));
    InMux I__8263 (
            .O(N__38886),
            .I(N__38877));
    LocalMux I__8262 (
            .O(N__38883),
            .I(\pid_front.pid_preregZ0Z_3 ));
    Odrv4 I__8261 (
            .O(N__38880),
            .I(\pid_front.pid_preregZ0Z_3 ));
    LocalMux I__8260 (
            .O(N__38877),
            .I(\pid_front.pid_preregZ0Z_3 ));
    InMux I__8259 (
            .O(N__38870),
            .I(N__38867));
    LocalMux I__8258 (
            .O(N__38867),
            .I(N__38864));
    Span12Mux_v I__8257 (
            .O(N__38864),
            .I(N__38861));
    Span12Mux_h I__8256 (
            .O(N__38861),
            .I(N__38858));
    Odrv12 I__8255 (
            .O(N__38858),
            .I(alt_ki_6));
    CEMux I__8254 (
            .O(N__38855),
            .I(N__38852));
    LocalMux I__8253 (
            .O(N__38852),
            .I(N__38849));
    Span4Mux_h I__8252 (
            .O(N__38849),
            .I(N__38845));
    CEMux I__8251 (
            .O(N__38848),
            .I(N__38842));
    Span4Mux_h I__8250 (
            .O(N__38845),
            .I(N__38836));
    LocalMux I__8249 (
            .O(N__38842),
            .I(N__38836));
    CEMux I__8248 (
            .O(N__38841),
            .I(N__38833));
    Span4Mux_h I__8247 (
            .O(N__38836),
            .I(N__38829));
    LocalMux I__8246 (
            .O(N__38833),
            .I(N__38826));
    CEMux I__8245 (
            .O(N__38832),
            .I(N__38823));
    Span4Mux_v I__8244 (
            .O(N__38829),
            .I(N__38820));
    Span4Mux_v I__8243 (
            .O(N__38826),
            .I(N__38815));
    LocalMux I__8242 (
            .O(N__38823),
            .I(N__38815));
    Span4Mux_v I__8241 (
            .O(N__38820),
            .I(N__38810));
    Span4Mux_h I__8240 (
            .O(N__38815),
            .I(N__38810));
    Odrv4 I__8239 (
            .O(N__38810),
            .I(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ));
    InMux I__8238 (
            .O(N__38807),
            .I(N__38803));
    InMux I__8237 (
            .O(N__38806),
            .I(N__38799));
    LocalMux I__8236 (
            .O(N__38803),
            .I(N__38796));
    InMux I__8235 (
            .O(N__38802),
            .I(N__38793));
    LocalMux I__8234 (
            .O(N__38799),
            .I(N__38790));
    Span4Mux_v I__8233 (
            .O(N__38796),
            .I(N__38787));
    LocalMux I__8232 (
            .O(N__38793),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__8231 (
            .O(N__38790),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    Odrv4 I__8230 (
            .O(N__38787),
            .I(\ppm_encoder_1.throttleZ0Z_6 ));
    InMux I__8229 (
            .O(N__38780),
            .I(N__38777));
    LocalMux I__8228 (
            .O(N__38777),
            .I(N__38772));
    InMux I__8227 (
            .O(N__38776),
            .I(N__38769));
    InMux I__8226 (
            .O(N__38775),
            .I(N__38766));
    Span4Mux_v I__8225 (
            .O(N__38772),
            .I(N__38763));
    LocalMux I__8224 (
            .O(N__38769),
            .I(N__38760));
    LocalMux I__8223 (
            .O(N__38766),
            .I(N__38753));
    Span4Mux_v I__8222 (
            .O(N__38763),
            .I(N__38753));
    Span4Mux_h I__8221 (
            .O(N__38760),
            .I(N__38753));
    Odrv4 I__8220 (
            .O(N__38753),
            .I(\ppm_encoder_1.rudderZ0Z_6 ));
    InMux I__8219 (
            .O(N__38750),
            .I(N__38747));
    LocalMux I__8218 (
            .O(N__38747),
            .I(N__38744));
    Span4Mux_v I__8217 (
            .O(N__38744),
            .I(N__38740));
    InMux I__8216 (
            .O(N__38743),
            .I(N__38737));
    Span4Mux_v I__8215 (
            .O(N__38740),
            .I(N__38734));
    LocalMux I__8214 (
            .O(N__38737),
            .I(N__38731));
    Odrv4 I__8213 (
            .O(N__38734),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    Odrv4 I__8212 (
            .O(N__38731),
            .I(\ppm_encoder_1.un1_init_pulses_0_6 ));
    CascadeMux I__8211 (
            .O(N__38726),
            .I(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ));
    CascadeMux I__8210 (
            .O(N__38723),
            .I(N__38720));
    InMux I__8209 (
            .O(N__38720),
            .I(N__38717));
    LocalMux I__8208 (
            .O(N__38717),
            .I(N__38714));
    Span4Mux_v I__8207 (
            .O(N__38714),
            .I(N__38711));
    Odrv4 I__8206 (
            .O(N__38711),
            .I(\ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ));
    InMux I__8205 (
            .O(N__38708),
            .I(N__38705));
    LocalMux I__8204 (
            .O(N__38705),
            .I(\ppm_encoder_1.un2_throttle_iv_1_6 ));
    CascadeMux I__8203 (
            .O(N__38702),
            .I(N__38699));
    InMux I__8202 (
            .O(N__38699),
            .I(N__38694));
    CascadeMux I__8201 (
            .O(N__38698),
            .I(N__38691));
    CascadeMux I__8200 (
            .O(N__38697),
            .I(N__38688));
    LocalMux I__8199 (
            .O(N__38694),
            .I(N__38685));
    InMux I__8198 (
            .O(N__38691),
            .I(N__38682));
    InMux I__8197 (
            .O(N__38688),
            .I(N__38679));
    Span4Mux_h I__8196 (
            .O(N__38685),
            .I(N__38674));
    LocalMux I__8195 (
            .O(N__38682),
            .I(N__38674));
    LocalMux I__8194 (
            .O(N__38679),
            .I(side_order_6));
    Odrv4 I__8193 (
            .O(N__38674),
            .I(side_order_6));
    InMux I__8192 (
            .O(N__38669),
            .I(N__38666));
    LocalMux I__8191 (
            .O(N__38666),
            .I(N__38663));
    Span4Mux_v I__8190 (
            .O(N__38663),
            .I(N__38660));
    Odrv4 I__8189 (
            .O(N__38660),
            .I(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ));
    InMux I__8188 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__8187 (
            .O(N__38654),
            .I(N__38649));
    CascadeMux I__8186 (
            .O(N__38653),
            .I(N__38646));
    InMux I__8185 (
            .O(N__38652),
            .I(N__38643));
    Span4Mux_h I__8184 (
            .O(N__38649),
            .I(N__38640));
    InMux I__8183 (
            .O(N__38646),
            .I(N__38637));
    LocalMux I__8182 (
            .O(N__38643),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    Odrv4 I__8181 (
            .O(N__38640),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    LocalMux I__8180 (
            .O(N__38637),
            .I(\ppm_encoder_1.aileronZ0Z_6 ));
    InMux I__8179 (
            .O(N__38630),
            .I(N__38627));
    LocalMux I__8178 (
            .O(N__38627),
            .I(N__38624));
    Span4Mux_h I__8177 (
            .O(N__38624),
            .I(N__38621));
    Span4Mux_v I__8176 (
            .O(N__38621),
            .I(N__38618));
    Odrv4 I__8175 (
            .O(N__38618),
            .I(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ));
    InMux I__8174 (
            .O(N__38615),
            .I(N__38610));
    InMux I__8173 (
            .O(N__38614),
            .I(N__38607));
    InMux I__8172 (
            .O(N__38613),
            .I(N__38604));
    LocalMux I__8171 (
            .O(N__38610),
            .I(N__38601));
    LocalMux I__8170 (
            .O(N__38607),
            .I(side_order_3));
    LocalMux I__8169 (
            .O(N__38604),
            .I(side_order_3));
    Odrv4 I__8168 (
            .O(N__38601),
            .I(side_order_3));
    InMux I__8167 (
            .O(N__38594),
            .I(N__38591));
    LocalMux I__8166 (
            .O(N__38591),
            .I(N__38588));
    Span4Mux_h I__8165 (
            .O(N__38588),
            .I(N__38585));
    Span4Mux_v I__8164 (
            .O(N__38585),
            .I(N__38582));
    Odrv4 I__8163 (
            .O(N__38582),
            .I(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ));
    InMux I__8162 (
            .O(N__38579),
            .I(N__38575));
    InMux I__8161 (
            .O(N__38578),
            .I(N__38572));
    LocalMux I__8160 (
            .O(N__38575),
            .I(N__38569));
    LocalMux I__8159 (
            .O(N__38572),
            .I(N__38566));
    Span4Mux_v I__8158 (
            .O(N__38569),
            .I(N__38563));
    Odrv4 I__8157 (
            .O(N__38566),
            .I(side_order_5));
    Odrv4 I__8156 (
            .O(N__38563),
            .I(side_order_5));
    InMux I__8155 (
            .O(N__38558),
            .I(N__38555));
    LocalMux I__8154 (
            .O(N__38555),
            .I(N__38551));
    CascadeMux I__8153 (
            .O(N__38554),
            .I(N__38547));
    Span4Mux_h I__8152 (
            .O(N__38551),
            .I(N__38544));
    CascadeMux I__8151 (
            .O(N__38550),
            .I(N__38541));
    InMux I__8150 (
            .O(N__38547),
            .I(N__38538));
    Span4Mux_h I__8149 (
            .O(N__38544),
            .I(N__38535));
    InMux I__8148 (
            .O(N__38541),
            .I(N__38532));
    LocalMux I__8147 (
            .O(N__38538),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    Odrv4 I__8146 (
            .O(N__38535),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    LocalMux I__8145 (
            .O(N__38532),
            .I(\ppm_encoder_1.aileronZ0Z_5 ));
    InMux I__8144 (
            .O(N__38525),
            .I(N__38521));
    CascadeMux I__8143 (
            .O(N__38524),
            .I(N__38518));
    LocalMux I__8142 (
            .O(N__38521),
            .I(N__38515));
    InMux I__8141 (
            .O(N__38518),
            .I(N__38511));
    Span4Mux_h I__8140 (
            .O(N__38515),
            .I(N__38508));
    InMux I__8139 (
            .O(N__38514),
            .I(N__38505));
    LocalMux I__8138 (
            .O(N__38511),
            .I(side_order_9));
    Odrv4 I__8137 (
            .O(N__38508),
            .I(side_order_9));
    LocalMux I__8136 (
            .O(N__38505),
            .I(side_order_9));
    InMux I__8135 (
            .O(N__38498),
            .I(N__38495));
    LocalMux I__8134 (
            .O(N__38495),
            .I(N__38492));
    Span4Mux_v I__8133 (
            .O(N__38492),
            .I(N__38489));
    Odrv4 I__8132 (
            .O(N__38489),
            .I(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ));
    InMux I__8131 (
            .O(N__38486),
            .I(N__38480));
    InMux I__8130 (
            .O(N__38485),
            .I(N__38480));
    LocalMux I__8129 (
            .O(N__38480),
            .I(N__38476));
    InMux I__8128 (
            .O(N__38479),
            .I(N__38473));
    Span4Mux_h I__8127 (
            .O(N__38476),
            .I(N__38470));
    LocalMux I__8126 (
            .O(N__38473),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    Odrv4 I__8125 (
            .O(N__38470),
            .I(\ppm_encoder_1.aileronZ0Z_9 ));
    CascadeMux I__8124 (
            .O(N__38465),
            .I(N__38461));
    InMux I__8123 (
            .O(N__38464),
            .I(N__38457));
    InMux I__8122 (
            .O(N__38461),
            .I(N__38454));
    InMux I__8121 (
            .O(N__38460),
            .I(N__38451));
    LocalMux I__8120 (
            .O(N__38457),
            .I(N__38448));
    LocalMux I__8119 (
            .O(N__38454),
            .I(N__38443));
    LocalMux I__8118 (
            .O(N__38451),
            .I(N__38443));
    Span4Mux_v I__8117 (
            .O(N__38448),
            .I(N__38440));
    Odrv12 I__8116 (
            .O(N__38443),
            .I(front_order_10));
    Odrv4 I__8115 (
            .O(N__38440),
            .I(front_order_10));
    InMux I__8114 (
            .O(N__38435),
            .I(N__38432));
    LocalMux I__8113 (
            .O(N__38432),
            .I(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ));
    InMux I__8112 (
            .O(N__38429),
            .I(N__38425));
    CascadeMux I__8111 (
            .O(N__38428),
            .I(N__38421));
    LocalMux I__8110 (
            .O(N__38425),
            .I(N__38418));
    InMux I__8109 (
            .O(N__38424),
            .I(N__38415));
    InMux I__8108 (
            .O(N__38421),
            .I(N__38412));
    Span4Mux_v I__8107 (
            .O(N__38418),
            .I(N__38409));
    LocalMux I__8106 (
            .O(N__38415),
            .I(N__38406));
    LocalMux I__8105 (
            .O(N__38412),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__8104 (
            .O(N__38409),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    Odrv4 I__8103 (
            .O(N__38406),
            .I(\ppm_encoder_1.elevatorZ0Z_10 ));
    InMux I__8102 (
            .O(N__38399),
            .I(N__38393));
    InMux I__8101 (
            .O(N__38398),
            .I(N__38393));
    LocalMux I__8100 (
            .O(N__38393),
            .I(N__38390));
    Span4Mux_v I__8099 (
            .O(N__38390),
            .I(N__38385));
    InMux I__8098 (
            .O(N__38389),
            .I(N__38380));
    InMux I__8097 (
            .O(N__38388),
            .I(N__38380));
    Odrv4 I__8096 (
            .O(N__38385),
            .I(\pid_side.N_563 ));
    LocalMux I__8095 (
            .O(N__38380),
            .I(\pid_side.N_563 ));
    CascadeMux I__8094 (
            .O(N__38375),
            .I(N__38372));
    InMux I__8093 (
            .O(N__38372),
            .I(N__38365));
    InMux I__8092 (
            .O(N__38371),
            .I(N__38365));
    CascadeMux I__8091 (
            .O(N__38370),
            .I(N__38362));
    LocalMux I__8090 (
            .O(N__38365),
            .I(N__38357));
    InMux I__8089 (
            .O(N__38362),
            .I(N__38354));
    InMux I__8088 (
            .O(N__38361),
            .I(N__38351));
    InMux I__8087 (
            .O(N__38360),
            .I(N__38348));
    Span4Mux_v I__8086 (
            .O(N__38357),
            .I(N__38345));
    LocalMux I__8085 (
            .O(N__38354),
            .I(N__38340));
    LocalMux I__8084 (
            .O(N__38351),
            .I(N__38340));
    LocalMux I__8083 (
            .O(N__38348),
            .I(N__38337));
    Span4Mux_h I__8082 (
            .O(N__38345),
            .I(N__38332));
    Span4Mux_h I__8081 (
            .O(N__38340),
            .I(N__38332));
    Span4Mux_h I__8080 (
            .O(N__38337),
            .I(N__38329));
    Span4Mux_h I__8079 (
            .O(N__38332),
            .I(N__38326));
    Span4Mux_h I__8078 (
            .O(N__38329),
            .I(N__38323));
    Odrv4 I__8077 (
            .O(N__38326),
            .I(\pid_side.pid_preregZ0Z_21 ));
    Odrv4 I__8076 (
            .O(N__38323),
            .I(\pid_side.pid_preregZ0Z_21 ));
    InMux I__8075 (
            .O(N__38318),
            .I(N__38309));
    InMux I__8074 (
            .O(N__38317),
            .I(N__38309));
    InMux I__8073 (
            .O(N__38316),
            .I(N__38306));
    InMux I__8072 (
            .O(N__38315),
            .I(N__38303));
    CascadeMux I__8071 (
            .O(N__38314),
            .I(N__38299));
    LocalMux I__8070 (
            .O(N__38309),
            .I(N__38296));
    LocalMux I__8069 (
            .O(N__38306),
            .I(N__38293));
    LocalMux I__8068 (
            .O(N__38303),
            .I(N__38290));
    InMux I__8067 (
            .O(N__38302),
            .I(N__38285));
    InMux I__8066 (
            .O(N__38299),
            .I(N__38285));
    Span4Mux_h I__8065 (
            .O(N__38296),
            .I(N__38281));
    Span4Mux_h I__8064 (
            .O(N__38293),
            .I(N__38274));
    Span4Mux_v I__8063 (
            .O(N__38290),
            .I(N__38274));
    LocalMux I__8062 (
            .O(N__38285),
            .I(N__38274));
    InMux I__8061 (
            .O(N__38284),
            .I(N__38271));
    Span4Mux_h I__8060 (
            .O(N__38281),
            .I(N__38268));
    Span4Mux_h I__8059 (
            .O(N__38274),
            .I(N__38265));
    LocalMux I__8058 (
            .O(N__38271),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__8057 (
            .O(N__38268),
            .I(\pid_side.pid_preregZ0Z_13 ));
    Odrv4 I__8056 (
            .O(N__38265),
            .I(\pid_side.pid_preregZ0Z_13 ));
    CascadeMux I__8055 (
            .O(N__38258),
            .I(N__38253));
    InMux I__8054 (
            .O(N__38257),
            .I(N__38250));
    InMux I__8053 (
            .O(N__38256),
            .I(N__38247));
    InMux I__8052 (
            .O(N__38253),
            .I(N__38243));
    LocalMux I__8051 (
            .O(N__38250),
            .I(N__38240));
    LocalMux I__8050 (
            .O(N__38247),
            .I(N__38237));
    InMux I__8049 (
            .O(N__38246),
            .I(N__38234));
    LocalMux I__8048 (
            .O(N__38243),
            .I(N__38231));
    Span4Mux_h I__8047 (
            .O(N__38240),
            .I(N__38227));
    Span4Mux_h I__8046 (
            .O(N__38237),
            .I(N__38224));
    LocalMux I__8045 (
            .O(N__38234),
            .I(N__38219));
    Span4Mux_v I__8044 (
            .O(N__38231),
            .I(N__38219));
    InMux I__8043 (
            .O(N__38230),
            .I(N__38216));
    Span4Mux_h I__8042 (
            .O(N__38227),
            .I(N__38213));
    Span4Mux_h I__8041 (
            .O(N__38224),
            .I(N__38208));
    Span4Mux_h I__8040 (
            .O(N__38219),
            .I(N__38208));
    LocalMux I__8039 (
            .O(N__38216),
            .I(\pid_side.pid_preregZ0Z_4 ));
    Odrv4 I__8038 (
            .O(N__38213),
            .I(\pid_side.pid_preregZ0Z_4 ));
    Odrv4 I__8037 (
            .O(N__38208),
            .I(\pid_side.pid_preregZ0Z_4 ));
    InMux I__8036 (
            .O(N__38201),
            .I(N__38195));
    InMux I__8035 (
            .O(N__38200),
            .I(N__38195));
    LocalMux I__8034 (
            .O(N__38195),
            .I(N__38192));
    Span4Mux_h I__8033 (
            .O(N__38192),
            .I(N__38188));
    InMux I__8032 (
            .O(N__38191),
            .I(N__38185));
    Odrv4 I__8031 (
            .O(N__38188),
            .I(\pid_side.N_534 ));
    LocalMux I__8030 (
            .O(N__38185),
            .I(\pid_side.N_534 ));
    CascadeMux I__8029 (
            .O(N__38180),
            .I(N__38176));
    InMux I__8028 (
            .O(N__38179),
            .I(N__38165));
    InMux I__8027 (
            .O(N__38176),
            .I(N__38165));
    InMux I__8026 (
            .O(N__38175),
            .I(N__38152));
    InMux I__8025 (
            .O(N__38174),
            .I(N__38152));
    InMux I__8024 (
            .O(N__38173),
            .I(N__38152));
    InMux I__8023 (
            .O(N__38172),
            .I(N__38152));
    InMux I__8022 (
            .O(N__38171),
            .I(N__38152));
    InMux I__8021 (
            .O(N__38170),
            .I(N__38152));
    LocalMux I__8020 (
            .O(N__38165),
            .I(\pid_side.N_291 ));
    LocalMux I__8019 (
            .O(N__38152),
            .I(\pid_side.N_291 ));
    CascadeMux I__8018 (
            .O(N__38147),
            .I(N__38144));
    InMux I__8017 (
            .O(N__38144),
            .I(N__38139));
    InMux I__8016 (
            .O(N__38143),
            .I(N__38133));
    InMux I__8015 (
            .O(N__38142),
            .I(N__38133));
    LocalMux I__8014 (
            .O(N__38139),
            .I(N__38130));
    InMux I__8013 (
            .O(N__38138),
            .I(N__38127));
    LocalMux I__8012 (
            .O(N__38133),
            .I(N__38124));
    Span4Mux_v I__8011 (
            .O(N__38130),
            .I(N__38118));
    LocalMux I__8010 (
            .O(N__38127),
            .I(N__38118));
    Span4Mux_v I__8009 (
            .O(N__38124),
            .I(N__38114));
    InMux I__8008 (
            .O(N__38123),
            .I(N__38111));
    Span4Mux_h I__8007 (
            .O(N__38118),
            .I(N__38108));
    InMux I__8006 (
            .O(N__38117),
            .I(N__38105));
    Sp12to4 I__8005 (
            .O(N__38114),
            .I(N__38100));
    LocalMux I__8004 (
            .O(N__38111),
            .I(N__38100));
    Span4Mux_h I__8003 (
            .O(N__38108),
            .I(N__38097));
    LocalMux I__8002 (
            .O(N__38105),
            .I(\pid_side.pid_preregZ0Z_5 ));
    Odrv12 I__8001 (
            .O(N__38100),
            .I(\pid_side.pid_preregZ0Z_5 ));
    Odrv4 I__8000 (
            .O(N__38097),
            .I(\pid_side.pid_preregZ0Z_5 ));
    CEMux I__7999 (
            .O(N__38090),
            .I(N__38087));
    LocalMux I__7998 (
            .O(N__38087),
            .I(N__38084));
    Span4Mux_h I__7997 (
            .O(N__38084),
            .I(N__38081));
    Span4Mux_v I__7996 (
            .O(N__38081),
            .I(N__38078));
    Odrv4 I__7995 (
            .O(N__38078),
            .I(\pid_side.state_0_1 ));
    SRMux I__7994 (
            .O(N__38075),
            .I(N__38070));
    SRMux I__7993 (
            .O(N__38074),
            .I(N__38067));
    SRMux I__7992 (
            .O(N__38073),
            .I(N__38064));
    LocalMux I__7991 (
            .O(N__38070),
            .I(N__38061));
    LocalMux I__7990 (
            .O(N__38067),
            .I(N__38057));
    LocalMux I__7989 (
            .O(N__38064),
            .I(N__38054));
    Span4Mux_h I__7988 (
            .O(N__38061),
            .I(N__38051));
    InMux I__7987 (
            .O(N__38060),
            .I(N__38048));
    Odrv4 I__7986 (
            .O(N__38057),
            .I(\pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ));
    Odrv4 I__7985 (
            .O(N__38054),
            .I(\pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ));
    Odrv4 I__7984 (
            .O(N__38051),
            .I(\pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ));
    LocalMux I__7983 (
            .O(N__38048),
            .I(\pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ));
    CascadeMux I__7982 (
            .O(N__38039),
            .I(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ));
    CascadeMux I__7981 (
            .O(N__38036),
            .I(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ));
    CascadeMux I__7980 (
            .O(N__38033),
            .I(N__38030));
    InMux I__7979 (
            .O(N__38030),
            .I(N__38027));
    LocalMux I__7978 (
            .O(N__38027),
            .I(N__38024));
    Span4Mux_v I__7977 (
            .O(N__38024),
            .I(N__38021));
    Odrv4 I__7976 (
            .O(N__38021),
            .I(\ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ));
    InMux I__7975 (
            .O(N__38018),
            .I(N__38013));
    CascadeMux I__7974 (
            .O(N__38017),
            .I(N__38010));
    InMux I__7973 (
            .O(N__38016),
            .I(N__38007));
    LocalMux I__7972 (
            .O(N__38013),
            .I(N__38004));
    InMux I__7971 (
            .O(N__38010),
            .I(N__38001));
    LocalMux I__7970 (
            .O(N__38007),
            .I(N__37996));
    Span4Mux_h I__7969 (
            .O(N__38004),
            .I(N__37996));
    LocalMux I__7968 (
            .O(N__38001),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    Odrv4 I__7967 (
            .O(N__37996),
            .I(\ppm_encoder_1.throttleZ0Z_5 ));
    CascadeMux I__7966 (
            .O(N__37991),
            .I(\ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ));
    InMux I__7965 (
            .O(N__37988),
            .I(N__37985));
    LocalMux I__7964 (
            .O(N__37985),
            .I(\ppm_encoder_1.un2_throttle_iv_0_5 ));
    CascadeMux I__7963 (
            .O(N__37982),
            .I(N__37979));
    InMux I__7962 (
            .O(N__37979),
            .I(N__37976));
    LocalMux I__7961 (
            .O(N__37976),
            .I(N__37973));
    Span4Mux_v I__7960 (
            .O(N__37973),
            .I(N__37970));
    Odrv4 I__7959 (
            .O(N__37970),
            .I(\ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ));
    InMux I__7958 (
            .O(N__37967),
            .I(N__37960));
    InMux I__7957 (
            .O(N__37966),
            .I(N__37960));
    InMux I__7956 (
            .O(N__37965),
            .I(N__37957));
    LocalMux I__7955 (
            .O(N__37960),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    LocalMux I__7954 (
            .O(N__37957),
            .I(\ppm_encoder_1.aileronZ0Z_1 ));
    CascadeMux I__7953 (
            .O(N__37952),
            .I(N__37948));
    CascadeMux I__7952 (
            .O(N__37951),
            .I(N__37944));
    InMux I__7951 (
            .O(N__37948),
            .I(N__37941));
    InMux I__7950 (
            .O(N__37947),
            .I(N__37938));
    InMux I__7949 (
            .O(N__37944),
            .I(N__37935));
    LocalMux I__7948 (
            .O(N__37941),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    LocalMux I__7947 (
            .O(N__37938),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    LocalMux I__7946 (
            .O(N__37935),
            .I(\ppm_encoder_1.elevatorZ0Z_1 ));
    CascadeMux I__7945 (
            .O(N__37928),
            .I(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ));
    InMux I__7944 (
            .O(N__37925),
            .I(N__37922));
    LocalMux I__7943 (
            .O(N__37922),
            .I(N__37918));
    InMux I__7942 (
            .O(N__37921),
            .I(N__37915));
    Odrv12 I__7941 (
            .O(N__37918),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    LocalMux I__7940 (
            .O(N__37915),
            .I(\ppm_encoder_1.un1_init_pulses_0_1 ));
    CascadeMux I__7939 (
            .O(N__37910),
            .I(N__37907));
    InMux I__7938 (
            .O(N__37907),
            .I(N__37904));
    LocalMux I__7937 (
            .O(N__37904),
            .I(N__37901));
    Span4Mux_h I__7936 (
            .O(N__37901),
            .I(N__37898));
    Odrv4 I__7935 (
            .O(N__37898),
            .I(\ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ));
    InMux I__7934 (
            .O(N__37895),
            .I(N__37890));
    InMux I__7933 (
            .O(N__37894),
            .I(N__37887));
    InMux I__7932 (
            .O(N__37893),
            .I(N__37884));
    LocalMux I__7931 (
            .O(N__37890),
            .I(N__37881));
    LocalMux I__7930 (
            .O(N__37887),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    LocalMux I__7929 (
            .O(N__37884),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    Odrv4 I__7928 (
            .O(N__37881),
            .I(\ppm_encoder_1.throttleZ0Z_1 ));
    CascadeMux I__7927 (
            .O(N__37874),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ));
    InMux I__7926 (
            .O(N__37871),
            .I(N__37868));
    LocalMux I__7925 (
            .O(N__37868),
            .I(\ppm_encoder_1.throttle_m_1 ));
    InMux I__7924 (
            .O(N__37865),
            .I(N__37859));
    InMux I__7923 (
            .O(N__37864),
            .I(N__37859));
    LocalMux I__7922 (
            .O(N__37859),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ));
    InMux I__7921 (
            .O(N__37856),
            .I(N__37852));
    InMux I__7920 (
            .O(N__37855),
            .I(N__37849));
    LocalMux I__7919 (
            .O(N__37852),
            .I(N__37844));
    LocalMux I__7918 (
            .O(N__37849),
            .I(N__37844));
    Span4Mux_v I__7917 (
            .O(N__37844),
            .I(N__37838));
    InMux I__7916 (
            .O(N__37843),
            .I(N__37833));
    InMux I__7915 (
            .O(N__37842),
            .I(N__37833));
    InMux I__7914 (
            .O(N__37841),
            .I(N__37830));
    Sp12to4 I__7913 (
            .O(N__37838),
            .I(N__37825));
    LocalMux I__7912 (
            .O(N__37833),
            .I(N__37825));
    LocalMux I__7911 (
            .O(N__37830),
            .I(\pid_side.pid_preregZ0Z_12 ));
    Odrv12 I__7910 (
            .O(N__37825),
            .I(\pid_side.pid_preregZ0Z_12 ));
    InMux I__7909 (
            .O(N__37820),
            .I(N__37816));
    InMux I__7908 (
            .O(N__37819),
            .I(N__37813));
    LocalMux I__7907 (
            .O(N__37816),
            .I(N__37810));
    LocalMux I__7906 (
            .O(N__37813),
            .I(N__37807));
    Span4Mux_v I__7905 (
            .O(N__37810),
            .I(N__37802));
    Span4Mux_v I__7904 (
            .O(N__37807),
            .I(N__37802));
    Odrv4 I__7903 (
            .O(N__37802),
            .I(side_order_12));
    InMux I__7902 (
            .O(N__37799),
            .I(N__37796));
    LocalMux I__7901 (
            .O(N__37796),
            .I(N__37791));
    InMux I__7900 (
            .O(N__37795),
            .I(N__37788));
    CascadeMux I__7899 (
            .O(N__37794),
            .I(N__37785));
    Span4Mux_h I__7898 (
            .O(N__37791),
            .I(N__37780));
    LocalMux I__7897 (
            .O(N__37788),
            .I(N__37780));
    InMux I__7896 (
            .O(N__37785),
            .I(N__37777));
    Span4Mux_h I__7895 (
            .O(N__37780),
            .I(N__37774));
    LocalMux I__7894 (
            .O(N__37777),
            .I(throttle_order_8));
    Odrv4 I__7893 (
            .O(N__37774),
            .I(throttle_order_8));
    CascadeMux I__7892 (
            .O(N__37769),
            .I(N__37766));
    InMux I__7891 (
            .O(N__37766),
            .I(N__37763));
    LocalMux I__7890 (
            .O(N__37763),
            .I(N__37760));
    Odrv12 I__7889 (
            .O(N__37760),
            .I(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ));
    InMux I__7888 (
            .O(N__37757),
            .I(N__37748));
    InMux I__7887 (
            .O(N__37756),
            .I(N__37748));
    InMux I__7886 (
            .O(N__37755),
            .I(N__37748));
    LocalMux I__7885 (
            .O(N__37748),
            .I(\ppm_encoder_1.throttleZ0Z_8 ));
    CascadeMux I__7884 (
            .O(N__37745),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ));
    InMux I__7883 (
            .O(N__37742),
            .I(N__37738));
    InMux I__7882 (
            .O(N__37741),
            .I(N__37734));
    LocalMux I__7881 (
            .O(N__37738),
            .I(N__37731));
    InMux I__7880 (
            .O(N__37737),
            .I(N__37728));
    LocalMux I__7879 (
            .O(N__37734),
            .I(N__37723));
    Span4Mux_h I__7878 (
            .O(N__37731),
            .I(N__37723));
    LocalMux I__7877 (
            .O(N__37728),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    Odrv4 I__7876 (
            .O(N__37723),
            .I(\ppm_encoder_1.throttleZ0Z_2 ));
    InMux I__7875 (
            .O(N__37718),
            .I(N__37715));
    LocalMux I__7874 (
            .O(N__37715),
            .I(N__37711));
    InMux I__7873 (
            .O(N__37714),
            .I(N__37707));
    Span4Mux_h I__7872 (
            .O(N__37711),
            .I(N__37704));
    InMux I__7871 (
            .O(N__37710),
            .I(N__37701));
    LocalMux I__7870 (
            .O(N__37707),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    Odrv4 I__7869 (
            .O(N__37704),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    LocalMux I__7868 (
            .O(N__37701),
            .I(\ppm_encoder_1.aileronZ0Z_2 ));
    InMux I__7867 (
            .O(N__37694),
            .I(N__37691));
    LocalMux I__7866 (
            .O(N__37691),
            .I(N__37688));
    Span12Mux_v I__7865 (
            .O(N__37688),
            .I(N__37684));
    InMux I__7864 (
            .O(N__37687),
            .I(N__37681));
    Odrv12 I__7863 (
            .O(N__37684),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    LocalMux I__7862 (
            .O(N__37681),
            .I(\ppm_encoder_1.un1_init_pulses_0_2 ));
    CascadeMux I__7861 (
            .O(N__37676),
            .I(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ));
    CascadeMux I__7860 (
            .O(N__37673),
            .I(N__37670));
    InMux I__7859 (
            .O(N__37670),
            .I(N__37667));
    LocalMux I__7858 (
            .O(N__37667),
            .I(N__37664));
    Odrv4 I__7857 (
            .O(N__37664),
            .I(\ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ));
    InMux I__7856 (
            .O(N__37661),
            .I(N__37658));
    LocalMux I__7855 (
            .O(N__37658),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ));
    CascadeMux I__7854 (
            .O(N__37655),
            .I(N__37652));
    InMux I__7853 (
            .O(N__37652),
            .I(N__37649));
    LocalMux I__7852 (
            .O(N__37649),
            .I(N__37646));
    Span4Mux_h I__7851 (
            .O(N__37646),
            .I(N__37643));
    Odrv4 I__7850 (
            .O(N__37643),
            .I(\ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ));
    InMux I__7849 (
            .O(N__37640),
            .I(N__37637));
    LocalMux I__7848 (
            .O(N__37637),
            .I(N__37634));
    Odrv4 I__7847 (
            .O(N__37634),
            .I(\ppm_encoder_1.un1_init_pulses_11_10 ));
    CascadeMux I__7846 (
            .O(N__37631),
            .I(N__37628));
    InMux I__7845 (
            .O(N__37628),
            .I(N__37625));
    LocalMux I__7844 (
            .O(N__37625),
            .I(\ppm_encoder_1.un1_init_pulses_10_10 ));
    InMux I__7843 (
            .O(N__37622),
            .I(N__37619));
    LocalMux I__7842 (
            .O(N__37619),
            .I(N__37616));
    Odrv12 I__7841 (
            .O(N__37616),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_10 ));
    CascadeMux I__7840 (
            .O(N__37613),
            .I(N__37610));
    InMux I__7839 (
            .O(N__37610),
            .I(N__37607));
    LocalMux I__7838 (
            .O(N__37607),
            .I(N__37602));
    InMux I__7837 (
            .O(N__37606),
            .I(N__37599));
    CascadeMux I__7836 (
            .O(N__37605),
            .I(N__37596));
    Span4Mux_h I__7835 (
            .O(N__37602),
            .I(N__37593));
    LocalMux I__7834 (
            .O(N__37599),
            .I(N__37590));
    InMux I__7833 (
            .O(N__37596),
            .I(N__37587));
    Span4Mux_v I__7832 (
            .O(N__37593),
            .I(N__37584));
    Span4Mux_h I__7831 (
            .O(N__37590),
            .I(N__37581));
    LocalMux I__7830 (
            .O(N__37587),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__7829 (
            .O(N__37584),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    Odrv4 I__7828 (
            .O(N__37581),
            .I(\ppm_encoder_1.rudderZ0Z_8 ));
    CascadeMux I__7827 (
            .O(N__37574),
            .I(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ));
    CascadeMux I__7826 (
            .O(N__37571),
            .I(N__37568));
    InMux I__7825 (
            .O(N__37568),
            .I(N__37565));
    LocalMux I__7824 (
            .O(N__37565),
            .I(\ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ));
    InMux I__7823 (
            .O(N__37562),
            .I(N__37559));
    LocalMux I__7822 (
            .O(N__37559),
            .I(\ppm_encoder_1.un2_throttle_iv_1_8 ));
    CascadeMux I__7821 (
            .O(N__37556),
            .I(\ppm_encoder_1.N_294_cascade_ ));
    InMux I__7820 (
            .O(N__37553),
            .I(N__37549));
    CascadeMux I__7819 (
            .O(N__37552),
            .I(N__37546));
    LocalMux I__7818 (
            .O(N__37549),
            .I(N__37543));
    InMux I__7817 (
            .O(N__37546),
            .I(N__37539));
    Span4Mux_v I__7816 (
            .O(N__37543),
            .I(N__37536));
    InMux I__7815 (
            .O(N__37542),
            .I(N__37533));
    LocalMux I__7814 (
            .O(N__37539),
            .I(side_order_8));
    Odrv4 I__7813 (
            .O(N__37536),
            .I(side_order_8));
    LocalMux I__7812 (
            .O(N__37533),
            .I(side_order_8));
    InMux I__7811 (
            .O(N__37526),
            .I(N__37523));
    LocalMux I__7810 (
            .O(N__37523),
            .I(N__37520));
    Span4Mux_h I__7809 (
            .O(N__37520),
            .I(N__37517));
    Odrv4 I__7808 (
            .O(N__37517),
            .I(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ));
    InMux I__7807 (
            .O(N__37514),
            .I(N__37505));
    InMux I__7806 (
            .O(N__37513),
            .I(N__37505));
    InMux I__7805 (
            .O(N__37512),
            .I(N__37505));
    LocalMux I__7804 (
            .O(N__37505),
            .I(\ppm_encoder_1.aileronZ0Z_8 ));
    InMux I__7803 (
            .O(N__37502),
            .I(N__37499));
    LocalMux I__7802 (
            .O(N__37499),
            .I(N__37495));
    InMux I__7801 (
            .O(N__37498),
            .I(N__37492));
    Span4Mux_v I__7800 (
            .O(N__37495),
            .I(N__37488));
    LocalMux I__7799 (
            .O(N__37492),
            .I(N__37485));
    InMux I__7798 (
            .O(N__37491),
            .I(N__37482));
    Span4Mux_h I__7797 (
            .O(N__37488),
            .I(N__37477));
    Span4Mux_h I__7796 (
            .O(N__37485),
            .I(N__37477));
    LocalMux I__7795 (
            .O(N__37482),
            .I(front_order_8));
    Odrv4 I__7794 (
            .O(N__37477),
            .I(front_order_8));
    InMux I__7793 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__7792 (
            .O(N__37469),
            .I(N__37466));
    Span4Mux_v I__7791 (
            .O(N__37466),
            .I(N__37463));
    Odrv4 I__7790 (
            .O(N__37463),
            .I(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ));
    InMux I__7789 (
            .O(N__37460),
            .I(N__37455));
    InMux I__7788 (
            .O(N__37459),
            .I(N__37450));
    InMux I__7787 (
            .O(N__37458),
            .I(N__37450));
    LocalMux I__7786 (
            .O(N__37455),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    LocalMux I__7785 (
            .O(N__37450),
            .I(\ppm_encoder_1.elevatorZ0Z_8 ));
    InMux I__7784 (
            .O(N__37445),
            .I(N__37442));
    LocalMux I__7783 (
            .O(N__37442),
            .I(N__37437));
    InMux I__7782 (
            .O(N__37441),
            .I(N__37432));
    InMux I__7781 (
            .O(N__37440),
            .I(N__37432));
    Span4Mux_v I__7780 (
            .O(N__37437),
            .I(N__37429));
    LocalMux I__7779 (
            .O(N__37432),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    Odrv4 I__7778 (
            .O(N__37429),
            .I(\ppm_encoder_1.init_pulsesZ0Z_14 ));
    InMux I__7777 (
            .O(N__37424),
            .I(N__37421));
    LocalMux I__7776 (
            .O(N__37421),
            .I(N__37418));
    Odrv4 I__7775 (
            .O(N__37418),
            .I(\ppm_encoder_1.un1_init_pulses_11_15 ));
    InMux I__7774 (
            .O(N__37415),
            .I(N__37412));
    LocalMux I__7773 (
            .O(N__37412),
            .I(\ppm_encoder_1.un1_init_pulses_10_15 ));
    InMux I__7772 (
            .O(N__37409),
            .I(N__37406));
    LocalMux I__7771 (
            .O(N__37406),
            .I(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ));
    InMux I__7770 (
            .O(N__37403),
            .I(N__37400));
    LocalMux I__7769 (
            .O(N__37400),
            .I(N__37397));
    Odrv12 I__7768 (
            .O(N__37397),
            .I(\ppm_encoder_1.un1_init_pulses_11_1 ));
    InMux I__7767 (
            .O(N__37394),
            .I(N__37391));
    LocalMux I__7766 (
            .O(N__37391),
            .I(\ppm_encoder_1.un1_init_pulses_10_1 ));
    InMux I__7765 (
            .O(N__37388),
            .I(N__37385));
    LocalMux I__7764 (
            .O(N__37385),
            .I(N__37382));
    Span4Mux_h I__7763 (
            .O(N__37382),
            .I(N__37379));
    Odrv4 I__7762 (
            .O(N__37379),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_1 ));
    InMux I__7761 (
            .O(N__37376),
            .I(N__37373));
    LocalMux I__7760 (
            .O(N__37373),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_8 ));
    CascadeMux I__7759 (
            .O(N__37370),
            .I(N__37367));
    InMux I__7758 (
            .O(N__37367),
            .I(N__37364));
    LocalMux I__7757 (
            .O(N__37364),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_9 ));
    CascadeMux I__7756 (
            .O(N__37361),
            .I(N__37358));
    InMux I__7755 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7754 (
            .O(N__37355),
            .I(N__37352));
    Odrv4 I__7753 (
            .O(N__37352),
            .I(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ));
    CascadeMux I__7752 (
            .O(N__37349),
            .I(\ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ));
    CascadeMux I__7751 (
            .O(N__37346),
            .I(N__37343));
    InMux I__7750 (
            .O(N__37343),
            .I(N__37340));
    LocalMux I__7749 (
            .O(N__37340),
            .I(N__37337));
    Odrv4 I__7748 (
            .O(N__37337),
            .I(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ));
    InMux I__7747 (
            .O(N__37334),
            .I(N__37331));
    LocalMux I__7746 (
            .O(N__37331),
            .I(N__37328));
    Odrv4 I__7745 (
            .O(N__37328),
            .I(\ppm_encoder_1.un1_init_pulses_11_13 ));
    InMux I__7744 (
            .O(N__37325),
            .I(N__37322));
    LocalMux I__7743 (
            .O(N__37322),
            .I(\ppm_encoder_1.un1_init_pulses_10_13 ));
    InMux I__7742 (
            .O(N__37319),
            .I(N__37316));
    LocalMux I__7741 (
            .O(N__37316),
            .I(N__37313));
    Odrv4 I__7740 (
            .O(N__37313),
            .I(\ppm_encoder_1.un1_init_pulses_11_14 ));
    InMux I__7739 (
            .O(N__37310),
            .I(N__37307));
    LocalMux I__7738 (
            .O(N__37307),
            .I(\ppm_encoder_1.un1_init_pulses_10_14 ));
    InMux I__7737 (
            .O(N__37304),
            .I(N__37301));
    LocalMux I__7736 (
            .O(N__37301),
            .I(N__37298));
    Odrv4 I__7735 (
            .O(N__37298),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_14 ));
    InMux I__7734 (
            .O(N__37295),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_9 ));
    InMux I__7733 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__7732 (
            .O(N__37289),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_11 ));
    CascadeMux I__7731 (
            .O(N__37286),
            .I(N__37283));
    InMux I__7730 (
            .O(N__37283),
            .I(N__37280));
    LocalMux I__7729 (
            .O(N__37280),
            .I(\ppm_encoder_1.un1_init_pulses_11_11 ));
    InMux I__7728 (
            .O(N__37277),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_10 ));
    CascadeMux I__7727 (
            .O(N__37274),
            .I(N__37271));
    InMux I__7726 (
            .O(N__37271),
            .I(N__37268));
    LocalMux I__7725 (
            .O(N__37268),
            .I(\ppm_encoder_1.un1_init_pulses_11_12 ));
    InMux I__7724 (
            .O(N__37265),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_11 ));
    InMux I__7723 (
            .O(N__37262),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_12 ));
    InMux I__7722 (
            .O(N__37259),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_13 ));
    InMux I__7721 (
            .O(N__37256),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_14 ));
    InMux I__7720 (
            .O(N__37253),
            .I(N__37250));
    LocalMux I__7719 (
            .O(N__37250),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_16 ));
    InMux I__7718 (
            .O(N__37247),
            .I(N__37244));
    LocalMux I__7717 (
            .O(N__37244),
            .I(\ppm_encoder_1.un1_init_pulses_11_16 ));
    InMux I__7716 (
            .O(N__37241),
            .I(bfn_16_10_0_));
    InMux I__7715 (
            .O(N__37238),
            .I(N__37235));
    LocalMux I__7714 (
            .O(N__37235),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_17 ));
    InMux I__7713 (
            .O(N__37232),
            .I(N__37229));
    LocalMux I__7712 (
            .O(N__37229),
            .I(\ppm_encoder_1.un1_init_pulses_11_17 ));
    InMux I__7711 (
            .O(N__37226),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_16 ));
    InMux I__7710 (
            .O(N__37223),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_17 ));
    InMux I__7709 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7708 (
            .O(N__37217),
            .I(\ppm_encoder_1.un1_init_pulses_11_18 ));
    CascadeMux I__7707 (
            .O(N__37214),
            .I(N__37211));
    InMux I__7706 (
            .O(N__37211),
            .I(N__37208));
    LocalMux I__7705 (
            .O(N__37208),
            .I(N__37205));
    Odrv4 I__7704 (
            .O(N__37205),
            .I(\ppm_encoder_1.un1_init_pulses_11_2 ));
    InMux I__7703 (
            .O(N__37202),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_1 ));
    InMux I__7702 (
            .O(N__37199),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_2 ));
    InMux I__7701 (
            .O(N__37196),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_3 ));
    InMux I__7700 (
            .O(N__37193),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_4 ));
    InMux I__7699 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__7698 (
            .O(N__37187),
            .I(N__37184));
    Span4Mux_h I__7697 (
            .O(N__37184),
            .I(N__37181));
    Odrv4 I__7696 (
            .O(N__37181),
            .I(\ppm_encoder_1.un1_init_pulses_11_6 ));
    InMux I__7695 (
            .O(N__37178),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_5 ));
    InMux I__7694 (
            .O(N__37175),
            .I(N__37172));
    LocalMux I__7693 (
            .O(N__37172),
            .I(N__37169));
    Span4Mux_h I__7692 (
            .O(N__37169),
            .I(N__37166));
    Odrv4 I__7691 (
            .O(N__37166),
            .I(\ppm_encoder_1.un1_init_pulses_3_axb_7 ));
    InMux I__7690 (
            .O(N__37163),
            .I(N__37160));
    LocalMux I__7689 (
            .O(N__37160),
            .I(N__37157));
    Span4Mux_h I__7688 (
            .O(N__37157),
            .I(N__37154));
    Odrv4 I__7687 (
            .O(N__37154),
            .I(\ppm_encoder_1.un1_init_pulses_11_7 ));
    InMux I__7686 (
            .O(N__37151),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_6 ));
    InMux I__7685 (
            .O(N__37148),
            .I(N__37145));
    LocalMux I__7684 (
            .O(N__37145),
            .I(N__37142));
    Span4Mux_h I__7683 (
            .O(N__37142),
            .I(N__37139));
    Odrv4 I__7682 (
            .O(N__37139),
            .I(\ppm_encoder_1.un1_init_pulses_11_8 ));
    InMux I__7681 (
            .O(N__37136),
            .I(bfn_16_9_0_));
    InMux I__7680 (
            .O(N__37133),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_8 ));
    InMux I__7679 (
            .O(N__37130),
            .I(N__37125));
    InMux I__7678 (
            .O(N__37129),
            .I(N__37122));
    InMux I__7677 (
            .O(N__37128),
            .I(N__37119));
    LocalMux I__7676 (
            .O(N__37125),
            .I(N__37115));
    LocalMux I__7675 (
            .O(N__37122),
            .I(N__37109));
    LocalMux I__7674 (
            .O(N__37119),
            .I(N__37106));
    InMux I__7673 (
            .O(N__37118),
            .I(N__37103));
    Span4Mux_h I__7672 (
            .O(N__37115),
            .I(N__37100));
    InMux I__7671 (
            .O(N__37114),
            .I(N__37097));
    InMux I__7670 (
            .O(N__37113),
            .I(N__37094));
    InMux I__7669 (
            .O(N__37112),
            .I(N__37091));
    Span12Mux_h I__7668 (
            .O(N__37109),
            .I(N__37084));
    Sp12to4 I__7667 (
            .O(N__37106),
            .I(N__37084));
    LocalMux I__7666 (
            .O(N__37103),
            .I(N__37084));
    Span4Mux_h I__7665 (
            .O(N__37100),
            .I(N__37081));
    LocalMux I__7664 (
            .O(N__37097),
            .I(N__37078));
    LocalMux I__7663 (
            .O(N__37094),
            .I(N__37075));
    LocalMux I__7662 (
            .O(N__37091),
            .I(N__37072));
    Span12Mux_v I__7661 (
            .O(N__37084),
            .I(N__37069));
    Sp12to4 I__7660 (
            .O(N__37081),
            .I(N__37062));
    Span12Mux_s10_h I__7659 (
            .O(N__37078),
            .I(N__37062));
    Sp12to4 I__7658 (
            .O(N__37075),
            .I(N__37062));
    Span4Mux_h I__7657 (
            .O(N__37072),
            .I(N__37059));
    Odrv12 I__7656 (
            .O(N__37069),
            .I(uart_drone_data_2));
    Odrv12 I__7655 (
            .O(N__37062),
            .I(uart_drone_data_2));
    Odrv4 I__7654 (
            .O(N__37059),
            .I(uart_drone_data_2));
    InMux I__7653 (
            .O(N__37052),
            .I(N__37049));
    LocalMux I__7652 (
            .O(N__37049),
            .I(N__37045));
    InMux I__7651 (
            .O(N__37048),
            .I(N__37041));
    Span4Mux_v I__7650 (
            .O(N__37045),
            .I(N__37038));
    InMux I__7649 (
            .O(N__37044),
            .I(N__37035));
    LocalMux I__7648 (
            .O(N__37041),
            .I(N__37031));
    Span4Mux_h I__7647 (
            .O(N__37038),
            .I(N__37026));
    LocalMux I__7646 (
            .O(N__37035),
            .I(N__37026));
    InMux I__7645 (
            .O(N__37034),
            .I(N__37023));
    Span4Mux_v I__7644 (
            .O(N__37031),
            .I(N__37019));
    Span4Mux_v I__7643 (
            .O(N__37026),
            .I(N__37014));
    LocalMux I__7642 (
            .O(N__37023),
            .I(N__37014));
    InMux I__7641 (
            .O(N__37022),
            .I(N__37011));
    Sp12to4 I__7640 (
            .O(N__37019),
            .I(N__37006));
    Span4Mux_h I__7639 (
            .O(N__37014),
            .I(N__37003));
    LocalMux I__7638 (
            .O(N__37011),
            .I(N__37000));
    InMux I__7637 (
            .O(N__37010),
            .I(N__36997));
    InMux I__7636 (
            .O(N__37009),
            .I(N__36993));
    Span12Mux_h I__7635 (
            .O(N__37006),
            .I(N__36984));
    Sp12to4 I__7634 (
            .O(N__37003),
            .I(N__36984));
    Sp12to4 I__7633 (
            .O(N__37000),
            .I(N__36984));
    LocalMux I__7632 (
            .O(N__36997),
            .I(N__36984));
    InMux I__7631 (
            .O(N__36996),
            .I(N__36981));
    LocalMux I__7630 (
            .O(N__36993),
            .I(N__36978));
    Odrv12 I__7629 (
            .O(N__36984),
            .I(uart_drone_data_3));
    LocalMux I__7628 (
            .O(N__36981),
            .I(uart_drone_data_3));
    Odrv4 I__7627 (
            .O(N__36978),
            .I(uart_drone_data_3));
    InMux I__7626 (
            .O(N__36971),
            .I(N__36966));
    InMux I__7625 (
            .O(N__36970),
            .I(N__36963));
    InMux I__7624 (
            .O(N__36969),
            .I(N__36960));
    LocalMux I__7623 (
            .O(N__36966),
            .I(N__36956));
    LocalMux I__7622 (
            .O(N__36963),
            .I(N__36953));
    LocalMux I__7621 (
            .O(N__36960),
            .I(N__36950));
    InMux I__7620 (
            .O(N__36959),
            .I(N__36947));
    Span4Mux_v I__7619 (
            .O(N__36956),
            .I(N__36943));
    Span4Mux_h I__7618 (
            .O(N__36953),
            .I(N__36940));
    Span4Mux_v I__7617 (
            .O(N__36950),
            .I(N__36935));
    LocalMux I__7616 (
            .O(N__36947),
            .I(N__36935));
    InMux I__7615 (
            .O(N__36946),
            .I(N__36931));
    Sp12to4 I__7614 (
            .O(N__36943),
            .I(N__36928));
    Span4Mux_h I__7613 (
            .O(N__36940),
            .I(N__36923));
    Span4Mux_h I__7612 (
            .O(N__36935),
            .I(N__36923));
    InMux I__7611 (
            .O(N__36934),
            .I(N__36920));
    LocalMux I__7610 (
            .O(N__36931),
            .I(N__36916));
    Span12Mux_h I__7609 (
            .O(N__36928),
            .I(N__36909));
    Sp12to4 I__7608 (
            .O(N__36923),
            .I(N__36909));
    LocalMux I__7607 (
            .O(N__36920),
            .I(N__36909));
    InMux I__7606 (
            .O(N__36919),
            .I(N__36905));
    Span12Mux_v I__7605 (
            .O(N__36916),
            .I(N__36902));
    Span12Mux_v I__7604 (
            .O(N__36909),
            .I(N__36899));
    InMux I__7603 (
            .O(N__36908),
            .I(N__36896));
    LocalMux I__7602 (
            .O(N__36905),
            .I(N__36893));
    Odrv12 I__7601 (
            .O(N__36902),
            .I(uart_drone_data_4));
    Odrv12 I__7600 (
            .O(N__36899),
            .I(uart_drone_data_4));
    LocalMux I__7599 (
            .O(N__36896),
            .I(uart_drone_data_4));
    Odrv4 I__7598 (
            .O(N__36893),
            .I(uart_drone_data_4));
    InMux I__7597 (
            .O(N__36884),
            .I(N__36881));
    LocalMux I__7596 (
            .O(N__36881),
            .I(N__36874));
    InMux I__7595 (
            .O(N__36880),
            .I(N__36871));
    InMux I__7594 (
            .O(N__36879),
            .I(N__36868));
    InMux I__7593 (
            .O(N__36878),
            .I(N__36865));
    InMux I__7592 (
            .O(N__36877),
            .I(N__36862));
    Span4Mux_v I__7591 (
            .O(N__36874),
            .I(N__36857));
    LocalMux I__7590 (
            .O(N__36871),
            .I(N__36857));
    LocalMux I__7589 (
            .O(N__36868),
            .I(N__36852));
    LocalMux I__7588 (
            .O(N__36865),
            .I(N__36852));
    LocalMux I__7587 (
            .O(N__36862),
            .I(N__36849));
    Span4Mux_v I__7586 (
            .O(N__36857),
            .I(N__36845));
    Span4Mux_v I__7585 (
            .O(N__36852),
            .I(N__36841));
    Span4Mux_v I__7584 (
            .O(N__36849),
            .I(N__36838));
    InMux I__7583 (
            .O(N__36848),
            .I(N__36835));
    Sp12to4 I__7582 (
            .O(N__36845),
            .I(N__36832));
    InMux I__7581 (
            .O(N__36844),
            .I(N__36829));
    Span4Mux_h I__7580 (
            .O(N__36841),
            .I(N__36822));
    Span4Mux_v I__7579 (
            .O(N__36838),
            .I(N__36822));
    LocalMux I__7578 (
            .O(N__36835),
            .I(N__36822));
    Span12Mux_h I__7577 (
            .O(N__36832),
            .I(N__36817));
    LocalMux I__7576 (
            .O(N__36829),
            .I(N__36817));
    Span4Mux_v I__7575 (
            .O(N__36822),
            .I(N__36814));
    Odrv12 I__7574 (
            .O(N__36817),
            .I(uart_drone_data_5));
    Odrv4 I__7573 (
            .O(N__36814),
            .I(uart_drone_data_5));
    InMux I__7572 (
            .O(N__36809),
            .I(N__36804));
    InMux I__7571 (
            .O(N__36808),
            .I(N__36800));
    InMux I__7570 (
            .O(N__36807),
            .I(N__36797));
    LocalMux I__7569 (
            .O(N__36804),
            .I(N__36793));
    InMux I__7568 (
            .O(N__36803),
            .I(N__36790));
    LocalMux I__7567 (
            .O(N__36800),
            .I(N__36784));
    LocalMux I__7566 (
            .O(N__36797),
            .I(N__36784));
    InMux I__7565 (
            .O(N__36796),
            .I(N__36781));
    Span4Mux_v I__7564 (
            .O(N__36793),
            .I(N__36778));
    LocalMux I__7563 (
            .O(N__36790),
            .I(N__36775));
    InMux I__7562 (
            .O(N__36789),
            .I(N__36772));
    Span4Mux_h I__7561 (
            .O(N__36784),
            .I(N__36767));
    LocalMux I__7560 (
            .O(N__36781),
            .I(N__36767));
    Span4Mux_h I__7559 (
            .O(N__36778),
            .I(N__36760));
    Span4Mux_h I__7558 (
            .O(N__36775),
            .I(N__36760));
    LocalMux I__7557 (
            .O(N__36772),
            .I(N__36760));
    Span4Mux_v I__7556 (
            .O(N__36767),
            .I(N__36756));
    Span4Mux_v I__7555 (
            .O(N__36760),
            .I(N__36753));
    InMux I__7554 (
            .O(N__36759),
            .I(N__36750));
    Span4Mux_h I__7553 (
            .O(N__36756),
            .I(N__36746));
    Span4Mux_v I__7552 (
            .O(N__36753),
            .I(N__36741));
    LocalMux I__7551 (
            .O(N__36750),
            .I(N__36741));
    InMux I__7550 (
            .O(N__36749),
            .I(N__36738));
    Odrv4 I__7549 (
            .O(N__36746),
            .I(uart_drone_data_1));
    Odrv4 I__7548 (
            .O(N__36741),
            .I(uart_drone_data_1));
    LocalMux I__7547 (
            .O(N__36738),
            .I(uart_drone_data_1));
    InMux I__7546 (
            .O(N__36731),
            .I(N__36727));
    CascadeMux I__7545 (
            .O(N__36730),
            .I(N__36724));
    LocalMux I__7544 (
            .O(N__36727),
            .I(N__36721));
    InMux I__7543 (
            .O(N__36724),
            .I(N__36718));
    Odrv12 I__7542 (
            .O(N__36721),
            .I(scaler_4_data_4));
    LocalMux I__7541 (
            .O(N__36718),
            .I(scaler_4_data_4));
    InMux I__7540 (
            .O(N__36713),
            .I(N__36710));
    LocalMux I__7539 (
            .O(N__36710),
            .I(N__36707));
    Span4Mux_h I__7538 (
            .O(N__36707),
            .I(N__36704));
    Span4Mux_h I__7537 (
            .O(N__36704),
            .I(N__36701));
    Odrv4 I__7536 (
            .O(N__36701),
            .I(scaler_4_data_5));
    CEMux I__7535 (
            .O(N__36698),
            .I(N__36694));
    CEMux I__7534 (
            .O(N__36697),
            .I(N__36689));
    LocalMux I__7533 (
            .O(N__36694),
            .I(N__36685));
    CEMux I__7532 (
            .O(N__36693),
            .I(N__36682));
    CEMux I__7531 (
            .O(N__36692),
            .I(N__36679));
    LocalMux I__7530 (
            .O(N__36689),
            .I(N__36676));
    CEMux I__7529 (
            .O(N__36688),
            .I(N__36673));
    Span4Mux_v I__7528 (
            .O(N__36685),
            .I(N__36670));
    LocalMux I__7527 (
            .O(N__36682),
            .I(N__36667));
    LocalMux I__7526 (
            .O(N__36679),
            .I(N__36664));
    Span4Mux_v I__7525 (
            .O(N__36676),
            .I(N__36661));
    LocalMux I__7524 (
            .O(N__36673),
            .I(N__36658));
    Span4Mux_h I__7523 (
            .O(N__36670),
            .I(N__36653));
    Span4Mux_v I__7522 (
            .O(N__36667),
            .I(N__36653));
    Span4Mux_v I__7521 (
            .O(N__36664),
            .I(N__36650));
    Span4Mux_h I__7520 (
            .O(N__36661),
            .I(N__36647));
    Span12Mux_h I__7519 (
            .O(N__36658),
            .I(N__36644));
    Odrv4 I__7518 (
            .O(N__36653),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__7517 (
            .O(N__36650),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv4 I__7516 (
            .O(N__36647),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    Odrv12 I__7515 (
            .O(N__36644),
            .I(\ppm_encoder_1.pid_altitude_dv_0 ));
    InMux I__7514 (
            .O(N__36635),
            .I(\ppm_encoder_1.un1_init_pulses_3_cry_0 ));
    InMux I__7513 (
            .O(N__36632),
            .I(N__36629));
    LocalMux I__7512 (
            .O(N__36629),
            .I(N__36624));
    InMux I__7511 (
            .O(N__36628),
            .I(N__36621));
    InMux I__7510 (
            .O(N__36627),
            .I(N__36617));
    Span4Mux_h I__7509 (
            .O(N__36624),
            .I(N__36613));
    LocalMux I__7508 (
            .O(N__36621),
            .I(N__36610));
    InMux I__7507 (
            .O(N__36620),
            .I(N__36606));
    LocalMux I__7506 (
            .O(N__36617),
            .I(N__36602));
    InMux I__7505 (
            .O(N__36616),
            .I(N__36599));
    Span4Mux_h I__7504 (
            .O(N__36613),
            .I(N__36594));
    Span4Mux_v I__7503 (
            .O(N__36610),
            .I(N__36594));
    InMux I__7502 (
            .O(N__36609),
            .I(N__36591));
    LocalMux I__7501 (
            .O(N__36606),
            .I(N__36588));
    InMux I__7500 (
            .O(N__36605),
            .I(N__36585));
    Span4Mux_v I__7499 (
            .O(N__36602),
            .I(N__36580));
    LocalMux I__7498 (
            .O(N__36599),
            .I(N__36580));
    Span4Mux_v I__7497 (
            .O(N__36594),
            .I(N__36575));
    LocalMux I__7496 (
            .O(N__36591),
            .I(N__36575));
    Sp12to4 I__7495 (
            .O(N__36588),
            .I(N__36570));
    LocalMux I__7494 (
            .O(N__36585),
            .I(N__36570));
    Span4Mux_h I__7493 (
            .O(N__36580),
            .I(N__36567));
    Span4Mux_v I__7492 (
            .O(N__36575),
            .I(N__36564));
    Span12Mux_v I__7491 (
            .O(N__36570),
            .I(N__36561));
    Span4Mux_v I__7490 (
            .O(N__36567),
            .I(N__36558));
    Span4Mux_h I__7489 (
            .O(N__36564),
            .I(N__36555));
    Odrv12 I__7488 (
            .O(N__36561),
            .I(uart_drone_data_7));
    Odrv4 I__7487 (
            .O(N__36558),
            .I(uart_drone_data_7));
    Odrv4 I__7486 (
            .O(N__36555),
            .I(uart_drone_data_7));
    CascadeMux I__7485 (
            .O(N__36548),
            .I(N__36545));
    InMux I__7484 (
            .O(N__36545),
            .I(N__36541));
    InMux I__7483 (
            .O(N__36544),
            .I(N__36538));
    LocalMux I__7482 (
            .O(N__36541),
            .I(\pid_front.pid_preregZ0Z_17 ));
    LocalMux I__7481 (
            .O(N__36538),
            .I(\pid_front.pid_preregZ0Z_17 ));
    InMux I__7480 (
            .O(N__36533),
            .I(N__36529));
    InMux I__7479 (
            .O(N__36532),
            .I(N__36526));
    LocalMux I__7478 (
            .O(N__36529),
            .I(\pid_front.pid_preregZ0Z_20 ));
    LocalMux I__7477 (
            .O(N__36526),
            .I(\pid_front.pid_preregZ0Z_20 ));
    CascadeMux I__7476 (
            .O(N__36521),
            .I(N__36517));
    InMux I__7475 (
            .O(N__36520),
            .I(N__36511));
    InMux I__7474 (
            .O(N__36517),
            .I(N__36511));
    CascadeMux I__7473 (
            .O(N__36516),
            .I(N__36507));
    LocalMux I__7472 (
            .O(N__36511),
            .I(N__36504));
    InMux I__7471 (
            .O(N__36510),
            .I(N__36501));
    InMux I__7470 (
            .O(N__36507),
            .I(N__36498));
    Span4Mux_h I__7469 (
            .O(N__36504),
            .I(N__36495));
    LocalMux I__7468 (
            .O(N__36501),
            .I(N__36492));
    LocalMux I__7467 (
            .O(N__36498),
            .I(\pid_front.pid_preregZ0Z_7 ));
    Odrv4 I__7466 (
            .O(N__36495),
            .I(\pid_front.pid_preregZ0Z_7 ));
    Odrv4 I__7465 (
            .O(N__36492),
            .I(\pid_front.pid_preregZ0Z_7 ));
    InMux I__7464 (
            .O(N__36485),
            .I(N__36479));
    InMux I__7463 (
            .O(N__36484),
            .I(N__36479));
    LocalMux I__7462 (
            .O(N__36479),
            .I(N__36474));
    InMux I__7461 (
            .O(N__36478),
            .I(N__36471));
    InMux I__7460 (
            .O(N__36477),
            .I(N__36468));
    Span4Mux_h I__7459 (
            .O(N__36474),
            .I(N__36465));
    LocalMux I__7458 (
            .O(N__36471),
            .I(N__36462));
    LocalMux I__7457 (
            .O(N__36468),
            .I(\pid_front.pid_preregZ0Z_6 ));
    Odrv4 I__7456 (
            .O(N__36465),
            .I(\pid_front.pid_preregZ0Z_6 ));
    Odrv4 I__7455 (
            .O(N__36462),
            .I(\pid_front.pid_preregZ0Z_6 ));
    InMux I__7454 (
            .O(N__36455),
            .I(N__36449));
    InMux I__7453 (
            .O(N__36454),
            .I(N__36446));
    InMux I__7452 (
            .O(N__36453),
            .I(N__36441));
    InMux I__7451 (
            .O(N__36452),
            .I(N__36441));
    LocalMux I__7450 (
            .O(N__36449),
            .I(N__36435));
    LocalMux I__7449 (
            .O(N__36446),
            .I(N__36435));
    LocalMux I__7448 (
            .O(N__36441),
            .I(N__36432));
    InMux I__7447 (
            .O(N__36440),
            .I(N__36429));
    Span4Mux_h I__7446 (
            .O(N__36435),
            .I(N__36426));
    Span4Mux_h I__7445 (
            .O(N__36432),
            .I(N__36423));
    LocalMux I__7444 (
            .O(N__36429),
            .I(\pid_front.pid_preregZ0Z_12 ));
    Odrv4 I__7443 (
            .O(N__36426),
            .I(\pid_front.pid_preregZ0Z_12 ));
    Odrv4 I__7442 (
            .O(N__36423),
            .I(\pid_front.pid_preregZ0Z_12 ));
    InMux I__7441 (
            .O(N__36416),
            .I(N__36412));
    InMux I__7440 (
            .O(N__36415),
            .I(N__36409));
    LocalMux I__7439 (
            .O(N__36412),
            .I(N__36406));
    LocalMux I__7438 (
            .O(N__36409),
            .I(\pid_front.pid_preregZ0Z_16 ));
    Odrv4 I__7437 (
            .O(N__36406),
            .I(\pid_front.pid_preregZ0Z_16 ));
    InMux I__7436 (
            .O(N__36401),
            .I(N__36398));
    LocalMux I__7435 (
            .O(N__36398),
            .I(N__36393));
    InMux I__7434 (
            .O(N__36397),
            .I(N__36390));
    InMux I__7433 (
            .O(N__36396),
            .I(N__36387));
    Span4Mux_h I__7432 (
            .O(N__36393),
            .I(N__36383));
    LocalMux I__7431 (
            .O(N__36390),
            .I(N__36380));
    LocalMux I__7430 (
            .O(N__36387),
            .I(N__36377));
    InMux I__7429 (
            .O(N__36386),
            .I(N__36374));
    Span4Mux_v I__7428 (
            .O(N__36383),
            .I(N__36371));
    Span4Mux_h I__7427 (
            .O(N__36380),
            .I(N__36368));
    Span4Mux_h I__7426 (
            .O(N__36377),
            .I(N__36365));
    LocalMux I__7425 (
            .O(N__36374),
            .I(\pid_front.pid_preregZ0Z_2 ));
    Odrv4 I__7424 (
            .O(N__36371),
            .I(\pid_front.pid_preregZ0Z_2 ));
    Odrv4 I__7423 (
            .O(N__36368),
            .I(\pid_front.pid_preregZ0Z_2 ));
    Odrv4 I__7422 (
            .O(N__36365),
            .I(\pid_front.pid_preregZ0Z_2 ));
    InMux I__7421 (
            .O(N__36356),
            .I(N__36352));
    InMux I__7420 (
            .O(N__36355),
            .I(N__36349));
    LocalMux I__7419 (
            .O(N__36352),
            .I(N__36346));
    LocalMux I__7418 (
            .O(N__36349),
            .I(\pid_front.pid_preregZ0Z_15 ));
    Odrv4 I__7417 (
            .O(N__36346),
            .I(\pid_front.pid_preregZ0Z_15 ));
    InMux I__7416 (
            .O(N__36341),
            .I(\ppm_encoder_1.un1_elevator_cry_8 ));
    InMux I__7415 (
            .O(N__36338),
            .I(\ppm_encoder_1.un1_elevator_cry_9 ));
    InMux I__7414 (
            .O(N__36335),
            .I(N__36330));
    InMux I__7413 (
            .O(N__36334),
            .I(N__36327));
    CascadeMux I__7412 (
            .O(N__36333),
            .I(N__36324));
    LocalMux I__7411 (
            .O(N__36330),
            .I(N__36321));
    LocalMux I__7410 (
            .O(N__36327),
            .I(N__36318));
    InMux I__7409 (
            .O(N__36324),
            .I(N__36315));
    Span12Mux_h I__7408 (
            .O(N__36321),
            .I(N__36312));
    Span4Mux_h I__7407 (
            .O(N__36318),
            .I(N__36309));
    LocalMux I__7406 (
            .O(N__36315),
            .I(front_order_11));
    Odrv12 I__7405 (
            .O(N__36312),
            .I(front_order_11));
    Odrv4 I__7404 (
            .O(N__36309),
            .I(front_order_11));
    CascadeMux I__7403 (
            .O(N__36302),
            .I(N__36299));
    InMux I__7402 (
            .O(N__36299),
            .I(N__36296));
    LocalMux I__7401 (
            .O(N__36296),
            .I(N__36293));
    Span4Mux_v I__7400 (
            .O(N__36293),
            .I(N__36290));
    Odrv4 I__7399 (
            .O(N__36290),
            .I(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ));
    InMux I__7398 (
            .O(N__36287),
            .I(\ppm_encoder_1.un1_elevator_cry_10 ));
    CascadeMux I__7397 (
            .O(N__36284),
            .I(N__36281));
    InMux I__7396 (
            .O(N__36281),
            .I(N__36278));
    LocalMux I__7395 (
            .O(N__36278),
            .I(N__36274));
    InMux I__7394 (
            .O(N__36277),
            .I(N__36271));
    Span4Mux_v I__7393 (
            .O(N__36274),
            .I(N__36268));
    LocalMux I__7392 (
            .O(N__36271),
            .I(N__36265));
    Odrv4 I__7391 (
            .O(N__36268),
            .I(front_order_12));
    Odrv4 I__7390 (
            .O(N__36265),
            .I(front_order_12));
    InMux I__7389 (
            .O(N__36260),
            .I(N__36257));
    LocalMux I__7388 (
            .O(N__36257),
            .I(N__36254));
    Span4Mux_h I__7387 (
            .O(N__36254),
            .I(N__36251));
    Span4Mux_v I__7386 (
            .O(N__36251),
            .I(N__36248));
    Odrv4 I__7385 (
            .O(N__36248),
            .I(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ));
    InMux I__7384 (
            .O(N__36245),
            .I(\ppm_encoder_1.un1_elevator_cry_11 ));
    InMux I__7383 (
            .O(N__36242),
            .I(\ppm_encoder_1.un1_elevator_cry_12 ));
    InMux I__7382 (
            .O(N__36239),
            .I(\ppm_encoder_1.un1_elevator_cry_13 ));
    InMux I__7381 (
            .O(N__36236),
            .I(N__36232));
    InMux I__7380 (
            .O(N__36235),
            .I(N__36228));
    LocalMux I__7379 (
            .O(N__36232),
            .I(N__36225));
    InMux I__7378 (
            .O(N__36231),
            .I(N__36222));
    LocalMux I__7377 (
            .O(N__36228),
            .I(N__36219));
    Span4Mux_h I__7376 (
            .O(N__36225),
            .I(N__36216));
    LocalMux I__7375 (
            .O(N__36222),
            .I(N__36213));
    Odrv4 I__7374 (
            .O(N__36219),
            .I(\pid_front.pid_preregZ0Z_0 ));
    Odrv4 I__7373 (
            .O(N__36216),
            .I(\pid_front.pid_preregZ0Z_0 ));
    Odrv4 I__7372 (
            .O(N__36213),
            .I(\pid_front.pid_preregZ0Z_0 ));
    InMux I__7371 (
            .O(N__36206),
            .I(N__36203));
    LocalMux I__7370 (
            .O(N__36203),
            .I(N__36200));
    Odrv4 I__7369 (
            .O(N__36200),
            .I(\pid_front.un1_reset_i_a5_1_7 ));
    InMux I__7368 (
            .O(N__36197),
            .I(N__36193));
    CascadeMux I__7367 (
            .O(N__36196),
            .I(N__36189));
    LocalMux I__7366 (
            .O(N__36193),
            .I(N__36186));
    InMux I__7365 (
            .O(N__36192),
            .I(N__36183));
    InMux I__7364 (
            .O(N__36189),
            .I(N__36180));
    Span4Mux_h I__7363 (
            .O(N__36186),
            .I(N__36177));
    LocalMux I__7362 (
            .O(N__36183),
            .I(N__36174));
    LocalMux I__7361 (
            .O(N__36180),
            .I(front_order_1));
    Odrv4 I__7360 (
            .O(N__36177),
            .I(front_order_1));
    Odrv4 I__7359 (
            .O(N__36174),
            .I(front_order_1));
    InMux I__7358 (
            .O(N__36167),
            .I(N__36164));
    LocalMux I__7357 (
            .O(N__36164),
            .I(N__36161));
    Odrv12 I__7356 (
            .O(N__36161),
            .I(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ));
    InMux I__7355 (
            .O(N__36158),
            .I(\ppm_encoder_1.un1_elevator_cry_0 ));
    InMux I__7354 (
            .O(N__36155),
            .I(\ppm_encoder_1.un1_elevator_cry_1 ));
    InMux I__7353 (
            .O(N__36152),
            .I(N__36149));
    LocalMux I__7352 (
            .O(N__36149),
            .I(N__36144));
    InMux I__7351 (
            .O(N__36148),
            .I(N__36141));
    InMux I__7350 (
            .O(N__36147),
            .I(N__36138));
    Span4Mux_v I__7349 (
            .O(N__36144),
            .I(N__36135));
    LocalMux I__7348 (
            .O(N__36141),
            .I(N__36132));
    LocalMux I__7347 (
            .O(N__36138),
            .I(front_order_3));
    Odrv4 I__7346 (
            .O(N__36135),
            .I(front_order_3));
    Odrv4 I__7345 (
            .O(N__36132),
            .I(front_order_3));
    InMux I__7344 (
            .O(N__36125),
            .I(N__36122));
    LocalMux I__7343 (
            .O(N__36122),
            .I(N__36119));
    Span4Mux_v I__7342 (
            .O(N__36119),
            .I(N__36116));
    Span4Mux_v I__7341 (
            .O(N__36116),
            .I(N__36113));
    Odrv4 I__7340 (
            .O(N__36113),
            .I(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ));
    InMux I__7339 (
            .O(N__36110),
            .I(\ppm_encoder_1.un1_elevator_cry_2 ));
    InMux I__7338 (
            .O(N__36107),
            .I(\ppm_encoder_1.un1_elevator_cry_3 ));
    InMux I__7337 (
            .O(N__36104),
            .I(\ppm_encoder_1.un1_elevator_cry_4 ));
    InMux I__7336 (
            .O(N__36101),
            .I(\ppm_encoder_1.un1_elevator_cry_5 ));
    InMux I__7335 (
            .O(N__36098),
            .I(\ppm_encoder_1.un1_elevator_cry_6 ));
    InMux I__7334 (
            .O(N__36095),
            .I(bfn_15_19_0_));
    InMux I__7333 (
            .O(N__36092),
            .I(N__36087));
    InMux I__7332 (
            .O(N__36091),
            .I(N__36084));
    CascadeMux I__7331 (
            .O(N__36090),
            .I(N__36081));
    LocalMux I__7330 (
            .O(N__36087),
            .I(N__36078));
    LocalMux I__7329 (
            .O(N__36084),
            .I(N__36075));
    InMux I__7328 (
            .O(N__36081),
            .I(N__36072));
    Span4Mux_v I__7327 (
            .O(N__36078),
            .I(N__36067));
    Span4Mux_v I__7326 (
            .O(N__36075),
            .I(N__36067));
    LocalMux I__7325 (
            .O(N__36072),
            .I(front_order_9));
    Odrv4 I__7324 (
            .O(N__36067),
            .I(front_order_9));
    InMux I__7323 (
            .O(N__36062),
            .I(N__36059));
    LocalMux I__7322 (
            .O(N__36059),
            .I(N__36056));
    Span4Mux_v I__7321 (
            .O(N__36056),
            .I(N__36053));
    Odrv4 I__7320 (
            .O(N__36053),
            .I(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ));
    CascadeMux I__7319 (
            .O(N__36050),
            .I(N__36047));
    InMux I__7318 (
            .O(N__36047),
            .I(N__36044));
    LocalMux I__7317 (
            .O(N__36044),
            .I(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ));
    CascadeMux I__7316 (
            .O(N__36041),
            .I(N__36038));
    InMux I__7315 (
            .O(N__36038),
            .I(N__36033));
    InMux I__7314 (
            .O(N__36037),
            .I(N__36030));
    InMux I__7313 (
            .O(N__36036),
            .I(N__36027));
    LocalMux I__7312 (
            .O(N__36033),
            .I(side_order_10));
    LocalMux I__7311 (
            .O(N__36030),
            .I(side_order_10));
    LocalMux I__7310 (
            .O(N__36027),
            .I(side_order_10));
    InMux I__7309 (
            .O(N__36020),
            .I(N__36011));
    InMux I__7308 (
            .O(N__36019),
            .I(N__36011));
    InMux I__7307 (
            .O(N__36018),
            .I(N__36011));
    LocalMux I__7306 (
            .O(N__36011),
            .I(\ppm_encoder_1.aileronZ0Z_10 ));
    InMux I__7305 (
            .O(N__36008),
            .I(N__36004));
    InMux I__7304 (
            .O(N__36007),
            .I(N__36001));
    LocalMux I__7303 (
            .O(N__36004),
            .I(N__35996));
    LocalMux I__7302 (
            .O(N__36001),
            .I(N__35996));
    Odrv12 I__7301 (
            .O(N__35996),
            .I(\pid_side.N_531 ));
    CascadeMux I__7300 (
            .O(N__35993),
            .I(N__35990));
    InMux I__7299 (
            .O(N__35990),
            .I(N__35987));
    LocalMux I__7298 (
            .O(N__35987),
            .I(\pid_side.un1_reset_i_a5_0_5 ));
    InMux I__7297 (
            .O(N__35984),
            .I(N__35981));
    LocalMux I__7296 (
            .O(N__35981),
            .I(\pid_side.un1_reset_i_1 ));
    InMux I__7295 (
            .O(N__35978),
            .I(N__35973));
    InMux I__7294 (
            .O(N__35977),
            .I(N__35970));
    InMux I__7293 (
            .O(N__35976),
            .I(N__35967));
    LocalMux I__7292 (
            .O(N__35973),
            .I(N__35962));
    LocalMux I__7291 (
            .O(N__35970),
            .I(N__35962));
    LocalMux I__7290 (
            .O(N__35967),
            .I(side_order_1));
    Odrv4 I__7289 (
            .O(N__35962),
            .I(side_order_1));
    InMux I__7288 (
            .O(N__35957),
            .I(N__35953));
    InMux I__7287 (
            .O(N__35956),
            .I(N__35950));
    LocalMux I__7286 (
            .O(N__35953),
            .I(N__35945));
    LocalMux I__7285 (
            .O(N__35950),
            .I(N__35942));
    InMux I__7284 (
            .O(N__35949),
            .I(N__35937));
    InMux I__7283 (
            .O(N__35948),
            .I(N__35937));
    Odrv4 I__7282 (
            .O(N__35945),
            .I(\pid_side.pid_preregZ0Z_2 ));
    Odrv4 I__7281 (
            .O(N__35942),
            .I(\pid_side.pid_preregZ0Z_2 ));
    LocalMux I__7280 (
            .O(N__35937),
            .I(\pid_side.pid_preregZ0Z_2 ));
    CascadeMux I__7279 (
            .O(N__35930),
            .I(N__35925));
    InMux I__7278 (
            .O(N__35929),
            .I(N__35922));
    CascadeMux I__7277 (
            .O(N__35928),
            .I(N__35919));
    InMux I__7276 (
            .O(N__35925),
            .I(N__35916));
    LocalMux I__7275 (
            .O(N__35922),
            .I(N__35913));
    InMux I__7274 (
            .O(N__35919),
            .I(N__35910));
    LocalMux I__7273 (
            .O(N__35916),
            .I(N__35907));
    Span4Mux_h I__7272 (
            .O(N__35913),
            .I(N__35904));
    LocalMux I__7271 (
            .O(N__35910),
            .I(side_order_2));
    Odrv12 I__7270 (
            .O(N__35907),
            .I(side_order_2));
    Odrv4 I__7269 (
            .O(N__35904),
            .I(side_order_2));
    InMux I__7268 (
            .O(N__35897),
            .I(N__35882));
    InMux I__7267 (
            .O(N__35896),
            .I(N__35879));
    InMux I__7266 (
            .O(N__35895),
            .I(N__35868));
    InMux I__7265 (
            .O(N__35894),
            .I(N__35868));
    InMux I__7264 (
            .O(N__35893),
            .I(N__35868));
    InMux I__7263 (
            .O(N__35892),
            .I(N__35868));
    InMux I__7262 (
            .O(N__35891),
            .I(N__35852));
    InMux I__7261 (
            .O(N__35890),
            .I(N__35852));
    InMux I__7260 (
            .O(N__35889),
            .I(N__35852));
    InMux I__7259 (
            .O(N__35888),
            .I(N__35852));
    InMux I__7258 (
            .O(N__35887),
            .I(N__35852));
    InMux I__7257 (
            .O(N__35886),
            .I(N__35852));
    InMux I__7256 (
            .O(N__35885),
            .I(N__35852));
    LocalMux I__7255 (
            .O(N__35882),
            .I(N__35849));
    LocalMux I__7254 (
            .O(N__35879),
            .I(N__35846));
    InMux I__7253 (
            .O(N__35878),
            .I(N__35843));
    CascadeMux I__7252 (
            .O(N__35877),
            .I(N__35840));
    LocalMux I__7251 (
            .O(N__35868),
            .I(N__35837));
    InMux I__7250 (
            .O(N__35867),
            .I(N__35834));
    LocalMux I__7249 (
            .O(N__35852),
            .I(N__35831));
    Span4Mux_h I__7248 (
            .O(N__35849),
            .I(N__35828));
    Span4Mux_v I__7247 (
            .O(N__35846),
            .I(N__35823));
    LocalMux I__7246 (
            .O(N__35843),
            .I(N__35823));
    InMux I__7245 (
            .O(N__35840),
            .I(N__35820));
    Span4Mux_h I__7244 (
            .O(N__35837),
            .I(N__35817));
    LocalMux I__7243 (
            .O(N__35834),
            .I(N__35814));
    Span4Mux_v I__7242 (
            .O(N__35831),
            .I(N__35809));
    Span4Mux_v I__7241 (
            .O(N__35828),
            .I(N__35809));
    Span4Mux_h I__7240 (
            .O(N__35823),
            .I(N__35806));
    LocalMux I__7239 (
            .O(N__35820),
            .I(N__35803));
    Odrv4 I__7238 (
            .O(N__35817),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__7237 (
            .O(N__35814),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__7236 (
            .O(N__35809),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv4 I__7235 (
            .O(N__35806),
            .I(\pid_side.stateZ0Z_1 ));
    Odrv12 I__7234 (
            .O(N__35803),
            .I(\pid_side.stateZ0Z_1 ));
    CascadeMux I__7233 (
            .O(N__35792),
            .I(N__35789));
    InMux I__7232 (
            .O(N__35789),
            .I(N__35784));
    InMux I__7231 (
            .O(N__35788),
            .I(N__35780));
    CascadeMux I__7230 (
            .O(N__35787),
            .I(N__35777));
    LocalMux I__7229 (
            .O(N__35784),
            .I(N__35774));
    InMux I__7228 (
            .O(N__35783),
            .I(N__35771));
    LocalMux I__7227 (
            .O(N__35780),
            .I(N__35768));
    InMux I__7226 (
            .O(N__35777),
            .I(N__35765));
    Span4Mux_h I__7225 (
            .O(N__35774),
            .I(N__35758));
    LocalMux I__7224 (
            .O(N__35771),
            .I(N__35758));
    Span4Mux_v I__7223 (
            .O(N__35768),
            .I(N__35758));
    LocalMux I__7222 (
            .O(N__35765),
            .I(\pid_side.pid_preregZ0Z_3 ));
    Odrv4 I__7221 (
            .O(N__35758),
            .I(\pid_side.pid_preregZ0Z_3 ));
    CascadeMux I__7220 (
            .O(N__35753),
            .I(\pid_side.N_291_cascade_ ));
    InMux I__7219 (
            .O(N__35750),
            .I(N__35738));
    InMux I__7218 (
            .O(N__35749),
            .I(N__35738));
    InMux I__7217 (
            .O(N__35748),
            .I(N__35738));
    InMux I__7216 (
            .O(N__35747),
            .I(N__35738));
    LocalMux I__7215 (
            .O(N__35738),
            .I(\pid_side.N_451_1 ));
    InMux I__7214 (
            .O(N__35735),
            .I(N__35732));
    LocalMux I__7213 (
            .O(N__35732),
            .I(N__35728));
    CascadeMux I__7212 (
            .O(N__35731),
            .I(N__35724));
    Span4Mux_h I__7211 (
            .O(N__35728),
            .I(N__35721));
    InMux I__7210 (
            .O(N__35727),
            .I(N__35718));
    InMux I__7209 (
            .O(N__35724),
            .I(N__35715));
    Span4Mux_v I__7208 (
            .O(N__35721),
            .I(N__35712));
    LocalMux I__7207 (
            .O(N__35718),
            .I(N__35709));
    LocalMux I__7206 (
            .O(N__35715),
            .I(front_order_0));
    Odrv4 I__7205 (
            .O(N__35712),
            .I(front_order_0));
    Odrv4 I__7204 (
            .O(N__35709),
            .I(front_order_0));
    InMux I__7203 (
            .O(N__35702),
            .I(N__35696));
    InMux I__7202 (
            .O(N__35701),
            .I(N__35696));
    LocalMux I__7201 (
            .O(N__35696),
            .I(N__35692));
    InMux I__7200 (
            .O(N__35695),
            .I(N__35689));
    Span4Mux_v I__7199 (
            .O(N__35692),
            .I(N__35686));
    LocalMux I__7198 (
            .O(N__35689),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    Odrv4 I__7197 (
            .O(N__35686),
            .I(\ppm_encoder_1.elevatorZ0Z_9 ));
    InMux I__7196 (
            .O(N__35681),
            .I(N__35678));
    LocalMux I__7195 (
            .O(N__35678),
            .I(\ppm_encoder_1.N_295 ));
    CascadeMux I__7194 (
            .O(N__35675),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ));
    InMux I__7193 (
            .O(N__35672),
            .I(N__35669));
    LocalMux I__7192 (
            .O(N__35669),
            .I(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ));
    InMux I__7191 (
            .O(N__35666),
            .I(N__35659));
    InMux I__7190 (
            .O(N__35665),
            .I(N__35659));
    InMux I__7189 (
            .O(N__35664),
            .I(N__35656));
    LocalMux I__7188 (
            .O(N__35659),
            .I(N__35653));
    LocalMux I__7187 (
            .O(N__35656),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    Odrv12 I__7186 (
            .O(N__35653),
            .I(\ppm_encoder_1.rudderZ0Z_9 ));
    InMux I__7185 (
            .O(N__35648),
            .I(N__35642));
    InMux I__7184 (
            .O(N__35647),
            .I(N__35642));
    LocalMux I__7183 (
            .O(N__35642),
            .I(N__35638));
    InMux I__7182 (
            .O(N__35641),
            .I(N__35635));
    Span4Mux_v I__7181 (
            .O(N__35638),
            .I(N__35632));
    LocalMux I__7180 (
            .O(N__35635),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    Odrv4 I__7179 (
            .O(N__35632),
            .I(\ppm_encoder_1.throttleZ0Z_9 ));
    InMux I__7178 (
            .O(N__35627),
            .I(N__35624));
    LocalMux I__7177 (
            .O(N__35624),
            .I(\ppm_encoder_1.un2_throttle_iv_0_9 ));
    InMux I__7176 (
            .O(N__35621),
            .I(N__35616));
    InMux I__7175 (
            .O(N__35620),
            .I(N__35613));
    InMux I__7174 (
            .O(N__35619),
            .I(N__35610));
    LocalMux I__7173 (
            .O(N__35616),
            .I(N__35607));
    LocalMux I__7172 (
            .O(N__35613),
            .I(N__35604));
    LocalMux I__7171 (
            .O(N__35610),
            .I(N__35597));
    Span4Mux_v I__7170 (
            .O(N__35607),
            .I(N__35597));
    Span4Mux_v I__7169 (
            .O(N__35604),
            .I(N__35597));
    Odrv4 I__7168 (
            .O(N__35597),
            .I(\ppm_encoder_1.throttleZ0Z_10 ));
    InMux I__7167 (
            .O(N__35594),
            .I(N__35591));
    LocalMux I__7166 (
            .O(N__35591),
            .I(N__35588));
    Span4Mux_v I__7165 (
            .O(N__35588),
            .I(N__35584));
    InMux I__7164 (
            .O(N__35587),
            .I(N__35581));
    Odrv4 I__7163 (
            .O(N__35584),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    LocalMux I__7162 (
            .O(N__35581),
            .I(\ppm_encoder_1.un1_init_pulses_0_10 ));
    CascadeMux I__7161 (
            .O(N__35576),
            .I(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ));
    CascadeMux I__7160 (
            .O(N__35573),
            .I(N__35570));
    InMux I__7159 (
            .O(N__35570),
            .I(N__35567));
    LocalMux I__7158 (
            .O(N__35567),
            .I(N__35564));
    Odrv12 I__7157 (
            .O(N__35564),
            .I(\ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ));
    InMux I__7156 (
            .O(N__35561),
            .I(N__35558));
    LocalMux I__7155 (
            .O(N__35558),
            .I(\ppm_encoder_1.un2_throttle_iv_1_10 ));
    InMux I__7154 (
            .O(N__35555),
            .I(N__35552));
    LocalMux I__7153 (
            .O(N__35552),
            .I(N__35549));
    Odrv12 I__7152 (
            .O(N__35549),
            .I(\ppm_encoder_1.N_296 ));
    InMux I__7151 (
            .O(N__35546),
            .I(N__35543));
    LocalMux I__7150 (
            .O(N__35543),
            .I(\ppm_encoder_1.N_287 ));
    InMux I__7149 (
            .O(N__35540),
            .I(N__35537));
    LocalMux I__7148 (
            .O(N__35537),
            .I(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ));
    InMux I__7147 (
            .O(N__35534),
            .I(N__35531));
    LocalMux I__7146 (
            .O(N__35531),
            .I(N__35528));
    Span4Mux_h I__7145 (
            .O(N__35528),
            .I(N__35525));
    Odrv4 I__7144 (
            .O(N__35525),
            .I(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ));
    InMux I__7143 (
            .O(N__35522),
            .I(N__35518));
    InMux I__7142 (
            .O(N__35521),
            .I(N__35514));
    LocalMux I__7141 (
            .O(N__35518),
            .I(N__35511));
    InMux I__7140 (
            .O(N__35517),
            .I(N__35508));
    LocalMux I__7139 (
            .O(N__35514),
            .I(N__35503));
    Span4Mux_v I__7138 (
            .O(N__35511),
            .I(N__35503));
    LocalMux I__7137 (
            .O(N__35508),
            .I(N__35500));
    Odrv4 I__7136 (
            .O(N__35503),
            .I(throttle_order_1));
    Odrv4 I__7135 (
            .O(N__35500),
            .I(throttle_order_1));
    InMux I__7134 (
            .O(N__35495),
            .I(N__35492));
    LocalMux I__7133 (
            .O(N__35492),
            .I(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ));
    CascadeMux I__7132 (
            .O(N__35489),
            .I(\ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ));
    CascadeMux I__7131 (
            .O(N__35486),
            .I(N__35483));
    InMux I__7130 (
            .O(N__35483),
            .I(N__35480));
    LocalMux I__7129 (
            .O(N__35480),
            .I(N__35477));
    Odrv4 I__7128 (
            .O(N__35477),
            .I(\ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ));
    InMux I__7127 (
            .O(N__35474),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_14 ));
    InMux I__7126 (
            .O(N__35471),
            .I(N__35468));
    LocalMux I__7125 (
            .O(N__35468),
            .I(N__35465));
    Odrv4 I__7124 (
            .O(N__35465),
            .I(\ppm_encoder_1.un1_init_pulses_10_16 ));
    InMux I__7123 (
            .O(N__35462),
            .I(bfn_15_13_0_));
    CascadeMux I__7122 (
            .O(N__35459),
            .I(N__35456));
    InMux I__7121 (
            .O(N__35456),
            .I(N__35453));
    LocalMux I__7120 (
            .O(N__35453),
            .I(N__35450));
    Odrv4 I__7119 (
            .O(N__35450),
            .I(\ppm_encoder_1.un1_init_pulses_0_axb_17 ));
    InMux I__7118 (
            .O(N__35447),
            .I(N__35444));
    LocalMux I__7117 (
            .O(N__35444),
            .I(N__35441));
    Odrv4 I__7116 (
            .O(N__35441),
            .I(\ppm_encoder_1.un1_init_pulses_10_17 ));
    InMux I__7115 (
            .O(N__35438),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_16 ));
    InMux I__7114 (
            .O(N__35435),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_17 ));
    InMux I__7113 (
            .O(N__35432),
            .I(N__35429));
    LocalMux I__7112 (
            .O(N__35429),
            .I(N__35426));
    Odrv4 I__7111 (
            .O(N__35426),
            .I(\ppm_encoder_1.un1_init_pulses_10_18 ));
    CascadeMux I__7110 (
            .O(N__35423),
            .I(N__35419));
    InMux I__7109 (
            .O(N__35422),
            .I(N__35416));
    InMux I__7108 (
            .O(N__35419),
            .I(N__35413));
    LocalMux I__7107 (
            .O(N__35416),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    LocalMux I__7106 (
            .O(N__35413),
            .I(\ppm_encoder_1.un1_init_pulses_0_12 ));
    InMux I__7105 (
            .O(N__35408),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_5 ));
    InMux I__7104 (
            .O(N__35405),
            .I(N__35402));
    LocalMux I__7103 (
            .O(N__35402),
            .I(\ppm_encoder_1.un1_init_pulses_10_7 ));
    InMux I__7102 (
            .O(N__35399),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_6 ));
    CascadeMux I__7101 (
            .O(N__35396),
            .I(N__35393));
    InMux I__7100 (
            .O(N__35393),
            .I(N__35390));
    LocalMux I__7099 (
            .O(N__35390),
            .I(N__35387));
    Odrv4 I__7098 (
            .O(N__35387),
            .I(\ppm_encoder_1.un1_init_pulses_10_8 ));
    InMux I__7097 (
            .O(N__35384),
            .I(bfn_15_12_0_));
    InMux I__7096 (
            .O(N__35381),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_8 ));
    InMux I__7095 (
            .O(N__35378),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_9 ));
    InMux I__7094 (
            .O(N__35375),
            .I(N__35372));
    LocalMux I__7093 (
            .O(N__35372),
            .I(N__35368));
    InMux I__7092 (
            .O(N__35371),
            .I(N__35365));
    Sp12to4 I__7091 (
            .O(N__35368),
            .I(N__35360));
    LocalMux I__7090 (
            .O(N__35365),
            .I(N__35360));
    Odrv12 I__7089 (
            .O(N__35360),
            .I(\ppm_encoder_1.un1_init_pulses_0_11 ));
    CascadeMux I__7088 (
            .O(N__35357),
            .I(N__35354));
    InMux I__7087 (
            .O(N__35354),
            .I(N__35351));
    LocalMux I__7086 (
            .O(N__35351),
            .I(\ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ));
    InMux I__7085 (
            .O(N__35348),
            .I(N__35345));
    LocalMux I__7084 (
            .O(N__35345),
            .I(N__35342));
    Odrv4 I__7083 (
            .O(N__35342),
            .I(\ppm_encoder_1.un1_init_pulses_10_11 ));
    InMux I__7082 (
            .O(N__35339),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_10 ));
    InMux I__7081 (
            .O(N__35336),
            .I(N__35333));
    LocalMux I__7080 (
            .O(N__35333),
            .I(\ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ));
    InMux I__7079 (
            .O(N__35330),
            .I(N__35327));
    LocalMux I__7078 (
            .O(N__35327),
            .I(N__35324));
    Odrv4 I__7077 (
            .O(N__35324),
            .I(\ppm_encoder_1.un1_init_pulses_10_12 ));
    InMux I__7076 (
            .O(N__35321),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_11 ));
    InMux I__7075 (
            .O(N__35318),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_12 ));
    InMux I__7074 (
            .O(N__35315),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_13 ));
    InMux I__7073 (
            .O(N__35312),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_0 ));
    InMux I__7072 (
            .O(N__35309),
            .I(N__35306));
    LocalMux I__7071 (
            .O(N__35306),
            .I(\ppm_encoder_1.un1_init_pulses_10_2 ));
    InMux I__7070 (
            .O(N__35303),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_1 ));
    InMux I__7069 (
            .O(N__35300),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_2 ));
    InMux I__7068 (
            .O(N__35297),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_3 ));
    InMux I__7067 (
            .O(N__35294),
            .I(\ppm_encoder_1.un1_init_pulses_0_cry_4 ));
    InMux I__7066 (
            .O(N__35291),
            .I(N__35288));
    LocalMux I__7065 (
            .O(N__35288),
            .I(\ppm_encoder_1.un1_init_pulses_10_6 ));
    InMux I__7064 (
            .O(N__35285),
            .I(N__35276));
    InMux I__7063 (
            .O(N__35284),
            .I(N__35276));
    InMux I__7062 (
            .O(N__35283),
            .I(N__35276));
    LocalMux I__7061 (
            .O(N__35276),
            .I(\ppm_encoder_1.init_pulsesZ0Z_11 ));
    InMux I__7060 (
            .O(N__35273),
            .I(N__35270));
    LocalMux I__7059 (
            .O(N__35270),
            .I(N__35265));
    InMux I__7058 (
            .O(N__35269),
            .I(N__35262));
    InMux I__7057 (
            .O(N__35268),
            .I(N__35259));
    Span4Mux_h I__7056 (
            .O(N__35265),
            .I(N__35254));
    LocalMux I__7055 (
            .O(N__35262),
            .I(N__35254));
    LocalMux I__7054 (
            .O(N__35259),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    Odrv4 I__7053 (
            .O(N__35254),
            .I(\ppm_encoder_1.rudderZ0Z_11 ));
    CascadeMux I__7052 (
            .O(N__35249),
            .I(\ppm_encoder_1.N_313_cascade_ ));
    InMux I__7051 (
            .O(N__35246),
            .I(N__35243));
    LocalMux I__7050 (
            .O(N__35243),
            .I(\reset_module_System.count_1_2 ));
    InMux I__7049 (
            .O(N__35240),
            .I(N__35236));
    InMux I__7048 (
            .O(N__35239),
            .I(N__35233));
    LocalMux I__7047 (
            .O(N__35236),
            .I(\reset_module_System.countZ0Z_2 ));
    LocalMux I__7046 (
            .O(N__35233),
            .I(\reset_module_System.countZ0Z_2 ));
    CascadeMux I__7045 (
            .O(N__35228),
            .I(N__35225));
    InMux I__7044 (
            .O(N__35225),
            .I(N__35216));
    InMux I__7043 (
            .O(N__35224),
            .I(N__35216));
    InMux I__7042 (
            .O(N__35223),
            .I(N__35216));
    LocalMux I__7041 (
            .O(N__35216),
            .I(\reset_module_System.reset6_15 ));
    CascadeMux I__7040 (
            .O(N__35213),
            .I(N__35208));
    InMux I__7039 (
            .O(N__35212),
            .I(N__35204));
    InMux I__7038 (
            .O(N__35211),
            .I(N__35201));
    InMux I__7037 (
            .O(N__35208),
            .I(N__35196));
    InMux I__7036 (
            .O(N__35207),
            .I(N__35196));
    LocalMux I__7035 (
            .O(N__35204),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__7034 (
            .O(N__35201),
            .I(\reset_module_System.reset6_14 ));
    LocalMux I__7033 (
            .O(N__35196),
            .I(\reset_module_System.reset6_14 ));
    InMux I__7032 (
            .O(N__35189),
            .I(N__35185));
    InMux I__7031 (
            .O(N__35188),
            .I(N__35182));
    LocalMux I__7030 (
            .O(N__35185),
            .I(\reset_module_System.countZ0Z_8 ));
    LocalMux I__7029 (
            .O(N__35182),
            .I(\reset_module_System.countZ0Z_8 ));
    InMux I__7028 (
            .O(N__35177),
            .I(N__35173));
    InMux I__7027 (
            .O(N__35176),
            .I(N__35170));
    LocalMux I__7026 (
            .O(N__35173),
            .I(\reset_module_System.countZ0Z_7 ));
    LocalMux I__7025 (
            .O(N__35170),
            .I(\reset_module_System.countZ0Z_7 ));
    CascadeMux I__7024 (
            .O(N__35165),
            .I(N__35161));
    InMux I__7023 (
            .O(N__35164),
            .I(N__35158));
    InMux I__7022 (
            .O(N__35161),
            .I(N__35155));
    LocalMux I__7021 (
            .O(N__35158),
            .I(\reset_module_System.countZ0Z_9 ));
    LocalMux I__7020 (
            .O(N__35155),
            .I(\reset_module_System.countZ0Z_9 ));
    InMux I__7019 (
            .O(N__35150),
            .I(N__35146));
    InMux I__7018 (
            .O(N__35149),
            .I(N__35143));
    LocalMux I__7017 (
            .O(N__35146),
            .I(\reset_module_System.countZ0Z_5 ));
    LocalMux I__7016 (
            .O(N__35143),
            .I(\reset_module_System.countZ0Z_5 ));
    InMux I__7015 (
            .O(N__35138),
            .I(N__35134));
    InMux I__7014 (
            .O(N__35137),
            .I(N__35131));
    LocalMux I__7013 (
            .O(N__35134),
            .I(\reset_module_System.countZ0Z_4 ));
    LocalMux I__7012 (
            .O(N__35131),
            .I(\reset_module_System.countZ0Z_4 ));
    InMux I__7011 (
            .O(N__35126),
            .I(N__35121));
    InMux I__7010 (
            .O(N__35125),
            .I(N__35118));
    InMux I__7009 (
            .O(N__35124),
            .I(N__35115));
    LocalMux I__7008 (
            .O(N__35121),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__7007 (
            .O(N__35118),
            .I(\reset_module_System.countZ0Z_1 ));
    LocalMux I__7006 (
            .O(N__35115),
            .I(\reset_module_System.countZ0Z_1 ));
    InMux I__7005 (
            .O(N__35108),
            .I(N__35105));
    LocalMux I__7004 (
            .O(N__35105),
            .I(N__35101));
    InMux I__7003 (
            .O(N__35104),
            .I(N__35098));
    Span4Mux_h I__7002 (
            .O(N__35101),
            .I(N__35095));
    LocalMux I__7001 (
            .O(N__35098),
            .I(\reset_module_System.countZ0Z_18 ));
    Odrv4 I__7000 (
            .O(N__35095),
            .I(\reset_module_System.countZ0Z_18 ));
    InMux I__6999 (
            .O(N__35090),
            .I(N__35086));
    InMux I__6998 (
            .O(N__35089),
            .I(N__35083));
    LocalMux I__6997 (
            .O(N__35086),
            .I(\reset_module_System.countZ0Z_16 ));
    LocalMux I__6996 (
            .O(N__35083),
            .I(\reset_module_System.countZ0Z_16 ));
    CascadeMux I__6995 (
            .O(N__35078),
            .I(\reset_module_System.reset6_3_cascade_ ));
    InMux I__6994 (
            .O(N__35075),
            .I(N__35072));
    LocalMux I__6993 (
            .O(N__35072),
            .I(\reset_module_System.reset6_13 ));
    InMux I__6992 (
            .O(N__35069),
            .I(N__35065));
    InMux I__6991 (
            .O(N__35068),
            .I(N__35062));
    LocalMux I__6990 (
            .O(N__35065),
            .I(\reset_module_System.countZ0Z_12 ));
    LocalMux I__6989 (
            .O(N__35062),
            .I(\reset_module_System.countZ0Z_12 ));
    CascadeMux I__6988 (
            .O(N__35057),
            .I(N__35051));
    InMux I__6987 (
            .O(N__35056),
            .I(N__35048));
    InMux I__6986 (
            .O(N__35055),
            .I(N__35045));
    InMux I__6985 (
            .O(N__35054),
            .I(N__35042));
    InMux I__6984 (
            .O(N__35051),
            .I(N__35039));
    LocalMux I__6983 (
            .O(N__35048),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__6982 (
            .O(N__35045),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__6981 (
            .O(N__35042),
            .I(\reset_module_System.countZ0Z_0 ));
    LocalMux I__6980 (
            .O(N__35039),
            .I(\reset_module_System.countZ0Z_0 ));
    CascadeMux I__6979 (
            .O(N__35030),
            .I(\reset_module_System.reset6_17_cascade_ ));
    InMux I__6978 (
            .O(N__35027),
            .I(N__35024));
    LocalMux I__6977 (
            .O(N__35024),
            .I(N__35021));
    Odrv4 I__6976 (
            .O(N__35021),
            .I(\reset_module_System.reset6_11 ));
    InMux I__6975 (
            .O(N__35018),
            .I(N__35012));
    InMux I__6974 (
            .O(N__35017),
            .I(N__35005));
    InMux I__6973 (
            .O(N__35016),
            .I(N__35005));
    InMux I__6972 (
            .O(N__35015),
            .I(N__35005));
    LocalMux I__6971 (
            .O(N__35012),
            .I(\reset_module_System.reset6_19 ));
    LocalMux I__6970 (
            .O(N__35005),
            .I(\reset_module_System.reset6_19 ));
    InMux I__6969 (
            .O(N__35000),
            .I(N__34997));
    LocalMux I__6968 (
            .O(N__34997),
            .I(N__34994));
    Span4Mux_v I__6967 (
            .O(N__34994),
            .I(N__34991));
    Span4Mux_h I__6966 (
            .O(N__34991),
            .I(N__34988));
    Odrv4 I__6965 (
            .O(N__34988),
            .I(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ));
    InMux I__6964 (
            .O(N__34985),
            .I(N__34982));
    LocalMux I__6963 (
            .O(N__34982),
            .I(N__34979));
    Span4Mux_h I__6962 (
            .O(N__34979),
            .I(N__34975));
    InMux I__6961 (
            .O(N__34978),
            .I(N__34972));
    Span4Mux_h I__6960 (
            .O(N__34975),
            .I(N__34969));
    LocalMux I__6959 (
            .O(N__34972),
            .I(N__34966));
    Odrv4 I__6958 (
            .O(N__34969),
            .I(scaler_4_data_9));
    Odrv4 I__6957 (
            .O(N__34966),
            .I(scaler_4_data_9));
    CascadeMux I__6956 (
            .O(N__34961),
            .I(N__34958));
    InMux I__6955 (
            .O(N__34958),
            .I(N__34955));
    LocalMux I__6954 (
            .O(N__34955),
            .I(\pid_front.m7_e_4 ));
    InMux I__6953 (
            .O(N__34952),
            .I(N__34948));
    InMux I__6952 (
            .O(N__34951),
            .I(N__34945));
    LocalMux I__6951 (
            .O(N__34948),
            .I(\pid_front.pid_preregZ0Z_18 ));
    LocalMux I__6950 (
            .O(N__34945),
            .I(\pid_front.pid_preregZ0Z_18 ));
    CascadeMux I__6949 (
            .O(N__34940),
            .I(N__34936));
    InMux I__6948 (
            .O(N__34939),
            .I(N__34933));
    InMux I__6947 (
            .O(N__34936),
            .I(N__34930));
    LocalMux I__6946 (
            .O(N__34933),
            .I(\pid_front.pid_preregZ0Z_19 ));
    LocalMux I__6945 (
            .O(N__34930),
            .I(\pid_front.pid_preregZ0Z_19 ));
    InMux I__6944 (
            .O(N__34925),
            .I(N__34918));
    InMux I__6943 (
            .O(N__34924),
            .I(N__34918));
    CascadeMux I__6942 (
            .O(N__34923),
            .I(N__34914));
    LocalMux I__6941 (
            .O(N__34918),
            .I(N__34911));
    CascadeMux I__6940 (
            .O(N__34917),
            .I(N__34908));
    InMux I__6939 (
            .O(N__34914),
            .I(N__34905));
    Span4Mux_v I__6938 (
            .O(N__34911),
            .I(N__34902));
    InMux I__6937 (
            .O(N__34908),
            .I(N__34899));
    LocalMux I__6936 (
            .O(N__34905),
            .I(\pid_front.pid_preregZ0Z_9 ));
    Odrv4 I__6935 (
            .O(N__34902),
            .I(\pid_front.pid_preregZ0Z_9 ));
    LocalMux I__6934 (
            .O(N__34899),
            .I(\pid_front.pid_preregZ0Z_9 ));
    InMux I__6933 (
            .O(N__34892),
            .I(N__34888));
    InMux I__6932 (
            .O(N__34891),
            .I(N__34885));
    LocalMux I__6931 (
            .O(N__34888),
            .I(N__34881));
    LocalMux I__6930 (
            .O(N__34885),
            .I(N__34878));
    InMux I__6929 (
            .O(N__34884),
            .I(N__34874));
    Span4Mux_v I__6928 (
            .O(N__34881),
            .I(N__34871));
    Span12Mux_v I__6927 (
            .O(N__34878),
            .I(N__34868));
    InMux I__6926 (
            .O(N__34877),
            .I(N__34865));
    LocalMux I__6925 (
            .O(N__34874),
            .I(\pid_front.pid_preregZ0Z_11 ));
    Odrv4 I__6924 (
            .O(N__34871),
            .I(\pid_front.pid_preregZ0Z_11 ));
    Odrv12 I__6923 (
            .O(N__34868),
            .I(\pid_front.pid_preregZ0Z_11 ));
    LocalMux I__6922 (
            .O(N__34865),
            .I(\pid_front.pid_preregZ0Z_11 ));
    InMux I__6921 (
            .O(N__34856),
            .I(N__34848));
    InMux I__6920 (
            .O(N__34855),
            .I(N__34848));
    InMux I__6919 (
            .O(N__34854),
            .I(N__34842));
    InMux I__6918 (
            .O(N__34853),
            .I(N__34842));
    LocalMux I__6917 (
            .O(N__34848),
            .I(N__34838));
    InMux I__6916 (
            .O(N__34847),
            .I(N__34835));
    LocalMux I__6915 (
            .O(N__34842),
            .I(N__34832));
    CascadeMux I__6914 (
            .O(N__34841),
            .I(N__34829));
    Span4Mux_h I__6913 (
            .O(N__34838),
            .I(N__34822));
    LocalMux I__6912 (
            .O(N__34835),
            .I(N__34822));
    Span4Mux_h I__6911 (
            .O(N__34832),
            .I(N__34822));
    InMux I__6910 (
            .O(N__34829),
            .I(N__34818));
    Span4Mux_v I__6909 (
            .O(N__34822),
            .I(N__34815));
    InMux I__6908 (
            .O(N__34821),
            .I(N__34812));
    LocalMux I__6907 (
            .O(N__34818),
            .I(\pid_front.pid_preregZ0Z_13 ));
    Odrv4 I__6906 (
            .O(N__34815),
            .I(\pid_front.pid_preregZ0Z_13 ));
    LocalMux I__6905 (
            .O(N__34812),
            .I(\pid_front.pid_preregZ0Z_13 ));
    InMux I__6904 (
            .O(N__34805),
            .I(N__34801));
    InMux I__6903 (
            .O(N__34804),
            .I(N__34798));
    LocalMux I__6902 (
            .O(N__34801),
            .I(N__34795));
    LocalMux I__6901 (
            .O(N__34798),
            .I(\pid_side.pid_preregZ0Z_15 ));
    Odrv12 I__6900 (
            .O(N__34795),
            .I(\pid_side.pid_preregZ0Z_15 ));
    CascadeMux I__6899 (
            .O(N__34790),
            .I(N__34786));
    InMux I__6898 (
            .O(N__34789),
            .I(N__34783));
    InMux I__6897 (
            .O(N__34786),
            .I(N__34780));
    LocalMux I__6896 (
            .O(N__34783),
            .I(N__34777));
    LocalMux I__6895 (
            .O(N__34780),
            .I(\pid_side.pid_preregZ0Z_14 ));
    Odrv12 I__6894 (
            .O(N__34777),
            .I(\pid_side.pid_preregZ0Z_14 ));
    CascadeMux I__6893 (
            .O(N__34772),
            .I(N__34769));
    InMux I__6892 (
            .O(N__34769),
            .I(N__34766));
    LocalMux I__6891 (
            .O(N__34766),
            .I(N__34763));
    Span4Mux_h I__6890 (
            .O(N__34763),
            .I(N__34760));
    Odrv4 I__6889 (
            .O(N__34760),
            .I(\pid_side.m7_e_4 ));
    InMux I__6888 (
            .O(N__34757),
            .I(N__34754));
    LocalMux I__6887 (
            .O(N__34754),
            .I(N__34750));
    InMux I__6886 (
            .O(N__34753),
            .I(N__34747));
    Span4Mux_v I__6885 (
            .O(N__34750),
            .I(N__34744));
    LocalMux I__6884 (
            .O(N__34747),
            .I(\pid_side.pid_preregZ0Z_16 ));
    Odrv4 I__6883 (
            .O(N__34744),
            .I(\pid_side.pid_preregZ0Z_16 ));
    InMux I__6882 (
            .O(N__34739),
            .I(N__34736));
    LocalMux I__6881 (
            .O(N__34736),
            .I(\pid_side.un1_reset_i_a5_1_7 ));
    CascadeMux I__6880 (
            .O(N__34733),
            .I(\pid_side.N_563_cascade_ ));
    InMux I__6879 (
            .O(N__34730),
            .I(N__34727));
    LocalMux I__6878 (
            .O(N__34727),
            .I(\pid_side.un1_reset_i_a5_1_8 ));
    CascadeMux I__6877 (
            .O(N__34724),
            .I(\pid_side.N_311_cascade_ ));
    InMux I__6876 (
            .O(N__34721),
            .I(N__34718));
    LocalMux I__6875 (
            .O(N__34718),
            .I(\pid_side.un1_reset_i_a5_1_6 ));
    InMux I__6874 (
            .O(N__34715),
            .I(N__34712));
    LocalMux I__6873 (
            .O(N__34712),
            .I(N__34709));
    Span4Mux_v I__6872 (
            .O(N__34709),
            .I(N__34705));
    InMux I__6871 (
            .O(N__34708),
            .I(N__34702));
    Span4Mux_h I__6870 (
            .O(N__34705),
            .I(N__34698));
    LocalMux I__6869 (
            .O(N__34702),
            .I(N__34695));
    InMux I__6868 (
            .O(N__34701),
            .I(N__34692));
    Sp12to4 I__6867 (
            .O(N__34698),
            .I(N__34687));
    Span12Mux_v I__6866 (
            .O(N__34695),
            .I(N__34687));
    LocalMux I__6865 (
            .O(N__34692),
            .I(\pid_side.error_p_regZ0Z_2 ));
    Odrv12 I__6864 (
            .O(N__34687),
            .I(\pid_side.error_p_regZ0Z_2 ));
    CascadeMux I__6863 (
            .O(N__34682),
            .I(N__34679));
    InMux I__6862 (
            .O(N__34679),
            .I(N__34676));
    LocalMux I__6861 (
            .O(N__34676),
            .I(N__34673));
    Span4Mux_h I__6860 (
            .O(N__34673),
            .I(N__34670));
    Span4Mux_h I__6859 (
            .O(N__34670),
            .I(N__34667));
    Odrv4 I__6858 (
            .O(N__34667),
            .I(\pid_side.un1_pid_prereg_cry_1_THRU_CO ));
    InMux I__6857 (
            .O(N__34664),
            .I(N__34661));
    LocalMux I__6856 (
            .O(N__34661),
            .I(N__34658));
    Odrv12 I__6855 (
            .O(N__34658),
            .I(\pid_side.un1_reset_i_a5_0_2 ));
    CascadeMux I__6854 (
            .O(N__34655),
            .I(N__34652));
    InMux I__6853 (
            .O(N__34652),
            .I(N__34649));
    LocalMux I__6852 (
            .O(N__34649),
            .I(N__34646));
    Odrv4 I__6851 (
            .O(N__34646),
            .I(\pid_side.un1_reset_i_a5_0_3 ));
    InMux I__6850 (
            .O(N__34643),
            .I(N__34637));
    InMux I__6849 (
            .O(N__34642),
            .I(N__34634));
    InMux I__6848 (
            .O(N__34641),
            .I(N__34628));
    InMux I__6847 (
            .O(N__34640),
            .I(N__34628));
    LocalMux I__6846 (
            .O(N__34637),
            .I(N__34625));
    LocalMux I__6845 (
            .O(N__34634),
            .I(N__34622));
    InMux I__6844 (
            .O(N__34633),
            .I(N__34619));
    LocalMux I__6843 (
            .O(N__34628),
            .I(\pid_front.N_569 ));
    Odrv4 I__6842 (
            .O(N__34625),
            .I(\pid_front.N_569 ));
    Odrv4 I__6841 (
            .O(N__34622),
            .I(\pid_front.N_569 ));
    LocalMux I__6840 (
            .O(N__34619),
            .I(\pid_front.N_569 ));
    InMux I__6839 (
            .O(N__34610),
            .I(N__34604));
    InMux I__6838 (
            .O(N__34609),
            .I(N__34604));
    LocalMux I__6837 (
            .O(N__34604),
            .I(\pid_front.pid_preregZ0Z_14 ));
    InMux I__6836 (
            .O(N__34601),
            .I(N__34598));
    LocalMux I__6835 (
            .O(N__34598),
            .I(N__34595));
    Span4Mux_v I__6834 (
            .O(N__34595),
            .I(N__34590));
    CascadeMux I__6833 (
            .O(N__34594),
            .I(N__34587));
    InMux I__6832 (
            .O(N__34593),
            .I(N__34583));
    Span4Mux_h I__6831 (
            .O(N__34590),
            .I(N__34580));
    InMux I__6830 (
            .O(N__34587),
            .I(N__34575));
    InMux I__6829 (
            .O(N__34586),
            .I(N__34575));
    LocalMux I__6828 (
            .O(N__34583),
            .I(\pid_side.pid_preregZ0Z_8 ));
    Odrv4 I__6827 (
            .O(N__34580),
            .I(\pid_side.pid_preregZ0Z_8 ));
    LocalMux I__6826 (
            .O(N__34575),
            .I(\pid_side.pid_preregZ0Z_8 ));
    InMux I__6825 (
            .O(N__34568),
            .I(N__34565));
    LocalMux I__6824 (
            .O(N__34565),
            .I(N__34562));
    Span4Mux_v I__6823 (
            .O(N__34562),
            .I(N__34556));
    InMux I__6822 (
            .O(N__34561),
            .I(N__34551));
    InMux I__6821 (
            .O(N__34560),
            .I(N__34551));
    InMux I__6820 (
            .O(N__34559),
            .I(N__34548));
    Span4Mux_h I__6819 (
            .O(N__34556),
            .I(N__34543));
    LocalMux I__6818 (
            .O(N__34551),
            .I(N__34543));
    LocalMux I__6817 (
            .O(N__34548),
            .I(\pid_side.pid_preregZ0Z_9 ));
    Odrv4 I__6816 (
            .O(N__34543),
            .I(\pid_side.pid_preregZ0Z_9 ));
    InMux I__6815 (
            .O(N__34538),
            .I(N__34526));
    InMux I__6814 (
            .O(N__34537),
            .I(N__34526));
    InMux I__6813 (
            .O(N__34536),
            .I(N__34526));
    InMux I__6812 (
            .O(N__34535),
            .I(N__34526));
    LocalMux I__6811 (
            .O(N__34526),
            .I(N__34521));
    InMux I__6810 (
            .O(N__34525),
            .I(N__34518));
    InMux I__6809 (
            .O(N__34524),
            .I(N__34511));
    Span4Mux_h I__6808 (
            .O(N__34521),
            .I(N__34506));
    LocalMux I__6807 (
            .O(N__34518),
            .I(N__34506));
    InMux I__6806 (
            .O(N__34517),
            .I(N__34503));
    InMux I__6805 (
            .O(N__34516),
            .I(N__34497));
    InMux I__6804 (
            .O(N__34515),
            .I(N__34497));
    InMux I__6803 (
            .O(N__34514),
            .I(N__34494));
    LocalMux I__6802 (
            .O(N__34511),
            .I(N__34489));
    Span4Mux_v I__6801 (
            .O(N__34506),
            .I(N__34489));
    LocalMux I__6800 (
            .O(N__34503),
            .I(N__34486));
    InMux I__6799 (
            .O(N__34502),
            .I(N__34483));
    LocalMux I__6798 (
            .O(N__34497),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__6797 (
            .O(N__34494),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__6796 (
            .O(N__34489),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    Odrv4 I__6795 (
            .O(N__34486),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    LocalMux I__6794 (
            .O(N__34483),
            .I(\uart_drone.bit_CountZ0Z_0 ));
    InMux I__6793 (
            .O(N__34472),
            .I(N__34469));
    LocalMux I__6792 (
            .O(N__34469),
            .I(N__34463));
    InMux I__6791 (
            .O(N__34468),
            .I(N__34456));
    InMux I__6790 (
            .O(N__34467),
            .I(N__34456));
    InMux I__6789 (
            .O(N__34466),
            .I(N__34456));
    Span4Mux_h I__6788 (
            .O(N__34463),
            .I(N__34453));
    LocalMux I__6787 (
            .O(N__34456),
            .I(\uart_drone.un1_state_4_0 ));
    Odrv4 I__6786 (
            .O(N__34453),
            .I(\uart_drone.un1_state_4_0 ));
    InMux I__6785 (
            .O(N__34448),
            .I(N__34445));
    LocalMux I__6784 (
            .O(N__34445),
            .I(N__34442));
    Odrv4 I__6783 (
            .O(N__34442),
            .I(\uart_drone.CO0 ));
    InMux I__6782 (
            .O(N__34439),
            .I(N__34436));
    LocalMux I__6781 (
            .O(N__34436),
            .I(N__34433));
    Span4Mux_v I__6780 (
            .O(N__34433),
            .I(N__34427));
    InMux I__6779 (
            .O(N__34432),
            .I(N__34424));
    InMux I__6778 (
            .O(N__34431),
            .I(N__34421));
    InMux I__6777 (
            .O(N__34430),
            .I(N__34418));
    Sp12to4 I__6776 (
            .O(N__34427),
            .I(N__34413));
    LocalMux I__6775 (
            .O(N__34424),
            .I(N__34413));
    LocalMux I__6774 (
            .O(N__34421),
            .I(\pid_side.pid_preregZ0Z_11 ));
    LocalMux I__6773 (
            .O(N__34418),
            .I(\pid_side.pid_preregZ0Z_11 ));
    Odrv12 I__6772 (
            .O(N__34413),
            .I(\pid_side.pid_preregZ0Z_11 ));
    InMux I__6771 (
            .O(N__34406),
            .I(N__34403));
    LocalMux I__6770 (
            .O(N__34403),
            .I(N__34397));
    InMux I__6769 (
            .O(N__34402),
            .I(N__34394));
    InMux I__6768 (
            .O(N__34401),
            .I(N__34391));
    InMux I__6767 (
            .O(N__34400),
            .I(N__34388));
    Span4Mux_v I__6766 (
            .O(N__34397),
            .I(N__34383));
    LocalMux I__6765 (
            .O(N__34394),
            .I(N__34383));
    LocalMux I__6764 (
            .O(N__34391),
            .I(\pid_side.pid_preregZ0Z_7 ));
    LocalMux I__6763 (
            .O(N__34388),
            .I(\pid_side.pid_preregZ0Z_7 ));
    Odrv4 I__6762 (
            .O(N__34383),
            .I(\pid_side.pid_preregZ0Z_7 ));
    InMux I__6761 (
            .O(N__34376),
            .I(N__34373));
    LocalMux I__6760 (
            .O(N__34373),
            .I(N__34370));
    Span4Mux_h I__6759 (
            .O(N__34370),
            .I(N__34367));
    Odrv4 I__6758 (
            .O(N__34367),
            .I(\pid_side.un1_reset_i_a5_1_5 ));
    InMux I__6757 (
            .O(N__34364),
            .I(N__34361));
    LocalMux I__6756 (
            .O(N__34361),
            .I(N__34358));
    Odrv12 I__6755 (
            .O(N__34358),
            .I(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ));
    InMux I__6754 (
            .O(N__34355),
            .I(\ppm_encoder_1.un1_aileron_cry_10 ));
    InMux I__6753 (
            .O(N__34352),
            .I(N__34349));
    LocalMux I__6752 (
            .O(N__34349),
            .I(N__34346));
    Odrv4 I__6751 (
            .O(N__34346),
            .I(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ));
    InMux I__6750 (
            .O(N__34343),
            .I(\ppm_encoder_1.un1_aileron_cry_11 ));
    InMux I__6749 (
            .O(N__34340),
            .I(\ppm_encoder_1.un1_aileron_cry_12 ));
    InMux I__6748 (
            .O(N__34337),
            .I(\ppm_encoder_1.un1_aileron_cry_13 ));
    InMux I__6747 (
            .O(N__34334),
            .I(N__34331));
    LocalMux I__6746 (
            .O(N__34331),
            .I(N__34328));
    Span4Mux_v I__6745 (
            .O(N__34328),
            .I(N__34323));
    InMux I__6744 (
            .O(N__34327),
            .I(N__34320));
    InMux I__6743 (
            .O(N__34326),
            .I(N__34317));
    Span4Mux_v I__6742 (
            .O(N__34323),
            .I(N__34314));
    LocalMux I__6741 (
            .O(N__34320),
            .I(N__34311));
    LocalMux I__6740 (
            .O(N__34317),
            .I(N__34308));
    Span4Mux_v I__6739 (
            .O(N__34314),
            .I(N__34303));
    Span4Mux_v I__6738 (
            .O(N__34311),
            .I(N__34303));
    Span12Mux_s1_h I__6737 (
            .O(N__34308),
            .I(N__34300));
    Sp12to4 I__6736 (
            .O(N__34303),
            .I(N__34297));
    Span12Mux_h I__6735 (
            .O(N__34300),
            .I(N__34293));
    Span12Mux_h I__6734 (
            .O(N__34297),
            .I(N__34290));
    InMux I__6733 (
            .O(N__34296),
            .I(N__34287));
    Odrv12 I__6732 (
            .O(N__34293),
            .I(drone_altitude_0));
    Odrv12 I__6731 (
            .O(N__34290),
            .I(drone_altitude_0));
    LocalMux I__6730 (
            .O(N__34287),
            .I(drone_altitude_0));
    CascadeMux I__6729 (
            .O(N__34280),
            .I(N__34277));
    InMux I__6728 (
            .O(N__34277),
            .I(N__34274));
    LocalMux I__6727 (
            .O(N__34274),
            .I(N__34270));
    InMux I__6726 (
            .O(N__34273),
            .I(N__34267));
    Span12Mux_v I__6725 (
            .O(N__34270),
            .I(N__34264));
    LocalMux I__6724 (
            .O(N__34267),
            .I(\pid_alt.drone_altitude_i_0 ));
    Odrv12 I__6723 (
            .O(N__34264),
            .I(\pid_alt.drone_altitude_i_0 ));
    InMux I__6722 (
            .O(N__34259),
            .I(N__34256));
    LocalMux I__6721 (
            .O(N__34256),
            .I(N__34253));
    Span4Mux_v I__6720 (
            .O(N__34253),
            .I(N__34250));
    Span4Mux_h I__6719 (
            .O(N__34250),
            .I(N__34244));
    InMux I__6718 (
            .O(N__34249),
            .I(N__34237));
    InMux I__6717 (
            .O(N__34248),
            .I(N__34237));
    InMux I__6716 (
            .O(N__34247),
            .I(N__34237));
    Odrv4 I__6715 (
            .O(N__34244),
            .I(\pid_side.pid_preregZ0Z_10 ));
    LocalMux I__6714 (
            .O(N__34237),
            .I(\pid_side.pid_preregZ0Z_10 ));
    CascadeMux I__6713 (
            .O(N__34232),
            .I(N__34228));
    InMux I__6712 (
            .O(N__34231),
            .I(N__34225));
    InMux I__6711 (
            .O(N__34228),
            .I(N__34221));
    LocalMux I__6710 (
            .O(N__34225),
            .I(N__34218));
    InMux I__6709 (
            .O(N__34224),
            .I(N__34215));
    LocalMux I__6708 (
            .O(N__34221),
            .I(side_order_11));
    Odrv12 I__6707 (
            .O(N__34218),
            .I(side_order_11));
    LocalMux I__6706 (
            .O(N__34215),
            .I(side_order_11));
    InMux I__6705 (
            .O(N__34208),
            .I(N__34205));
    LocalMux I__6704 (
            .O(N__34205),
            .I(N__34201));
    CascadeMux I__6703 (
            .O(N__34204),
            .I(N__34197));
    Span4Mux_h I__6702 (
            .O(N__34201),
            .I(N__34194));
    CascadeMux I__6701 (
            .O(N__34200),
            .I(N__34190));
    InMux I__6700 (
            .O(N__34197),
            .I(N__34187));
    Span4Mux_h I__6699 (
            .O(N__34194),
            .I(N__34184));
    InMux I__6698 (
            .O(N__34193),
            .I(N__34181));
    InMux I__6697 (
            .O(N__34190),
            .I(N__34178));
    LocalMux I__6696 (
            .O(N__34187),
            .I(\pid_side.pid_preregZ0Z_6 ));
    Odrv4 I__6695 (
            .O(N__34184),
            .I(\pid_side.pid_preregZ0Z_6 ));
    LocalMux I__6694 (
            .O(N__34181),
            .I(\pid_side.pid_preregZ0Z_6 ));
    LocalMux I__6693 (
            .O(N__34178),
            .I(\pid_side.pid_preregZ0Z_6 ));
    InMux I__6692 (
            .O(N__34169),
            .I(\ppm_encoder_1.un1_aileron_cry_1 ));
    InMux I__6691 (
            .O(N__34166),
            .I(\ppm_encoder_1.un1_aileron_cry_2 ));
    InMux I__6690 (
            .O(N__34163),
            .I(\ppm_encoder_1.un1_aileron_cry_3 ));
    InMux I__6689 (
            .O(N__34160),
            .I(\ppm_encoder_1.un1_aileron_cry_4 ));
    InMux I__6688 (
            .O(N__34157),
            .I(\ppm_encoder_1.un1_aileron_cry_5 ));
    InMux I__6687 (
            .O(N__34154),
            .I(\ppm_encoder_1.un1_aileron_cry_6 ));
    InMux I__6686 (
            .O(N__34151),
            .I(bfn_14_15_0_));
    InMux I__6685 (
            .O(N__34148),
            .I(\ppm_encoder_1.un1_aileron_cry_8 ));
    InMux I__6684 (
            .O(N__34145),
            .I(\ppm_encoder_1.un1_aileron_cry_9 ));
    InMux I__6683 (
            .O(N__34142),
            .I(N__34137));
    InMux I__6682 (
            .O(N__34141),
            .I(N__34134));
    InMux I__6681 (
            .O(N__34140),
            .I(N__34131));
    LocalMux I__6680 (
            .O(N__34137),
            .I(N__34128));
    LocalMux I__6679 (
            .O(N__34134),
            .I(N__34125));
    LocalMux I__6678 (
            .O(N__34131),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv12 I__6677 (
            .O(N__34128),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    Odrv4 I__6676 (
            .O(N__34125),
            .I(\ppm_encoder_1.rudderZ0Z_12 ));
    CascadeMux I__6675 (
            .O(N__34118),
            .I(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ));
    InMux I__6674 (
            .O(N__34115),
            .I(N__34112));
    LocalMux I__6673 (
            .O(N__34112),
            .I(\ppm_encoder_1.un2_throttle_iv_1_12 ));
    CascadeMux I__6672 (
            .O(N__34109),
            .I(N__34104));
    InMux I__6671 (
            .O(N__34108),
            .I(N__34099));
    InMux I__6670 (
            .O(N__34107),
            .I(N__34099));
    InMux I__6669 (
            .O(N__34104),
            .I(N__34096));
    LocalMux I__6668 (
            .O(N__34099),
            .I(N__34093));
    LocalMux I__6667 (
            .O(N__34096),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    Odrv4 I__6666 (
            .O(N__34093),
            .I(\ppm_encoder_1.throttleZ0Z_12 ));
    CascadeMux I__6665 (
            .O(N__34088),
            .I(\ppm_encoder_1.N_298_cascade_ ));
    CascadeMux I__6664 (
            .O(N__34085),
            .I(N__34080));
    InMux I__6663 (
            .O(N__34084),
            .I(N__34075));
    InMux I__6662 (
            .O(N__34083),
            .I(N__34075));
    InMux I__6661 (
            .O(N__34080),
            .I(N__34072));
    LocalMux I__6660 (
            .O(N__34075),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    LocalMux I__6659 (
            .O(N__34072),
            .I(\ppm_encoder_1.aileronZ0Z_12 ));
    InMux I__6658 (
            .O(N__34067),
            .I(N__34062));
    InMux I__6657 (
            .O(N__34066),
            .I(N__34057));
    InMux I__6656 (
            .O(N__34065),
            .I(N__34057));
    LocalMux I__6655 (
            .O(N__34062),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    LocalMux I__6654 (
            .O(N__34057),
            .I(\ppm_encoder_1.elevatorZ0Z_12 ));
    InMux I__6653 (
            .O(N__34052),
            .I(\ppm_encoder_1.un1_aileron_cry_0 ));
    InMux I__6652 (
            .O(N__34049),
            .I(N__34046));
    LocalMux I__6651 (
            .O(N__34046),
            .I(N__34042));
    CascadeMux I__6650 (
            .O(N__34045),
            .I(N__34039));
    Span4Mux_v I__6649 (
            .O(N__34042),
            .I(N__34036));
    InMux I__6648 (
            .O(N__34039),
            .I(N__34033));
    Span4Mux_h I__6647 (
            .O(N__34036),
            .I(N__34030));
    LocalMux I__6646 (
            .O(N__34033),
            .I(N__34027));
    Odrv4 I__6645 (
            .O(N__34030),
            .I(scaler_4_data_10));
    Odrv4 I__6644 (
            .O(N__34027),
            .I(scaler_4_data_10));
    InMux I__6643 (
            .O(N__34022),
            .I(N__34019));
    LocalMux I__6642 (
            .O(N__34019),
            .I(N__34016));
    Span4Mux_v I__6641 (
            .O(N__34016),
            .I(N__34013));
    Odrv4 I__6640 (
            .O(N__34013),
            .I(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ));
    CascadeMux I__6639 (
            .O(N__34010),
            .I(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ));
    InMux I__6638 (
            .O(N__34007),
            .I(N__34004));
    LocalMux I__6637 (
            .O(N__34004),
            .I(\ppm_encoder_1.un2_throttle_iv_1_11 ));
    InMux I__6636 (
            .O(N__34001),
            .I(N__33996));
    InMux I__6635 (
            .O(N__34000),
            .I(N__33991));
    InMux I__6634 (
            .O(N__33999),
            .I(N__33991));
    LocalMux I__6633 (
            .O(N__33996),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    LocalMux I__6632 (
            .O(N__33991),
            .I(\ppm_encoder_1.throttleZ0Z_11 ));
    CascadeMux I__6631 (
            .O(N__33986),
            .I(\ppm_encoder_1.N_297_cascade_ ));
    InMux I__6630 (
            .O(N__33983),
            .I(N__33974));
    InMux I__6629 (
            .O(N__33982),
            .I(N__33974));
    InMux I__6628 (
            .O(N__33981),
            .I(N__33974));
    LocalMux I__6627 (
            .O(N__33974),
            .I(\ppm_encoder_1.aileronZ0Z_11 ));
    InMux I__6626 (
            .O(N__33971),
            .I(N__33962));
    InMux I__6625 (
            .O(N__33970),
            .I(N__33962));
    InMux I__6624 (
            .O(N__33969),
            .I(N__33962));
    LocalMux I__6623 (
            .O(N__33962),
            .I(\ppm_encoder_1.elevatorZ0Z_11 ));
    CascadeMux I__6622 (
            .O(N__33959),
            .I(N__33956));
    InMux I__6621 (
            .O(N__33956),
            .I(N__33952));
    InMux I__6620 (
            .O(N__33955),
            .I(N__33949));
    LocalMux I__6619 (
            .O(N__33952),
            .I(N__33946));
    LocalMux I__6618 (
            .O(N__33949),
            .I(\reset_module_System.countZ0Z_20 ));
    Odrv4 I__6617 (
            .O(N__33946),
            .I(\reset_module_System.countZ0Z_20 ));
    InMux I__6616 (
            .O(N__33941),
            .I(\reset_module_System.count_1_cry_19 ));
    InMux I__6615 (
            .O(N__33938),
            .I(\reset_module_System.count_1_cry_20 ));
    CascadeMux I__6614 (
            .O(N__33935),
            .I(N__33932));
    InMux I__6613 (
            .O(N__33932),
            .I(N__33926));
    InMux I__6612 (
            .O(N__33931),
            .I(N__33926));
    LocalMux I__6611 (
            .O(N__33926),
            .I(\reset_module_System.countZ0Z_19 ));
    InMux I__6610 (
            .O(N__33923),
            .I(N__33919));
    InMux I__6609 (
            .O(N__33922),
            .I(N__33916));
    LocalMux I__6608 (
            .O(N__33919),
            .I(\reset_module_System.countZ0Z_15 ));
    LocalMux I__6607 (
            .O(N__33916),
            .I(\reset_module_System.countZ0Z_15 ));
    CascadeMux I__6606 (
            .O(N__33911),
            .I(N__33907));
    InMux I__6605 (
            .O(N__33910),
            .I(N__33902));
    InMux I__6604 (
            .O(N__33907),
            .I(N__33902));
    LocalMux I__6603 (
            .O(N__33902),
            .I(\reset_module_System.countZ0Z_21 ));
    InMux I__6602 (
            .O(N__33899),
            .I(N__33895));
    InMux I__6601 (
            .O(N__33898),
            .I(N__33892));
    LocalMux I__6600 (
            .O(N__33895),
            .I(\reset_module_System.countZ0Z_13 ));
    LocalMux I__6599 (
            .O(N__33892),
            .I(\reset_module_System.countZ0Z_13 ));
    InMux I__6598 (
            .O(N__33887),
            .I(N__33884));
    LocalMux I__6597 (
            .O(N__33884),
            .I(N__33880));
    InMux I__6596 (
            .O(N__33883),
            .I(N__33877));
    Odrv4 I__6595 (
            .O(N__33880),
            .I(\reset_module_System.countZ0Z_11 ));
    LocalMux I__6594 (
            .O(N__33877),
            .I(\reset_module_System.countZ0Z_11 ));
    InMux I__6593 (
            .O(N__33872),
            .I(\reset_module_System.count_1_cry_10 ));
    InMux I__6592 (
            .O(N__33869),
            .I(\reset_module_System.count_1_cry_11 ));
    InMux I__6591 (
            .O(N__33866),
            .I(\reset_module_System.count_1_cry_12 ));
    InMux I__6590 (
            .O(N__33863),
            .I(N__33860));
    LocalMux I__6589 (
            .O(N__33860),
            .I(N__33856));
    InMux I__6588 (
            .O(N__33859),
            .I(N__33853));
    Odrv4 I__6587 (
            .O(N__33856),
            .I(\reset_module_System.countZ0Z_14 ));
    LocalMux I__6586 (
            .O(N__33853),
            .I(\reset_module_System.countZ0Z_14 ));
    InMux I__6585 (
            .O(N__33848),
            .I(\reset_module_System.count_1_cry_13 ));
    InMux I__6584 (
            .O(N__33845),
            .I(\reset_module_System.count_1_cry_14 ));
    InMux I__6583 (
            .O(N__33842),
            .I(\reset_module_System.count_1_cry_15 ));
    CascadeMux I__6582 (
            .O(N__33839),
            .I(N__33836));
    InMux I__6581 (
            .O(N__33836),
            .I(N__33833));
    LocalMux I__6580 (
            .O(N__33833),
            .I(N__33829));
    InMux I__6579 (
            .O(N__33832),
            .I(N__33826));
    Odrv12 I__6578 (
            .O(N__33829),
            .I(\reset_module_System.countZ0Z_17 ));
    LocalMux I__6577 (
            .O(N__33826),
            .I(\reset_module_System.countZ0Z_17 ));
    InMux I__6576 (
            .O(N__33821),
            .I(bfn_14_9_0_));
    InMux I__6575 (
            .O(N__33818),
            .I(\reset_module_System.count_1_cry_17 ));
    InMux I__6574 (
            .O(N__33815),
            .I(\reset_module_System.count_1_cry_18 ));
    InMux I__6573 (
            .O(N__33812),
            .I(\reset_module_System.count_1_cry_1 ));
    InMux I__6572 (
            .O(N__33809),
            .I(N__33805));
    InMux I__6571 (
            .O(N__33808),
            .I(N__33802));
    LocalMux I__6570 (
            .O(N__33805),
            .I(\reset_module_System.countZ0Z_3 ));
    LocalMux I__6569 (
            .O(N__33802),
            .I(\reset_module_System.countZ0Z_3 ));
    InMux I__6568 (
            .O(N__33797),
            .I(\reset_module_System.count_1_cry_2 ));
    InMux I__6567 (
            .O(N__33794),
            .I(\reset_module_System.count_1_cry_3 ));
    InMux I__6566 (
            .O(N__33791),
            .I(\reset_module_System.count_1_cry_4 ));
    InMux I__6565 (
            .O(N__33788),
            .I(N__33784));
    InMux I__6564 (
            .O(N__33787),
            .I(N__33781));
    LocalMux I__6563 (
            .O(N__33784),
            .I(\reset_module_System.countZ0Z_6 ));
    LocalMux I__6562 (
            .O(N__33781),
            .I(\reset_module_System.countZ0Z_6 ));
    InMux I__6561 (
            .O(N__33776),
            .I(\reset_module_System.count_1_cry_5 ));
    InMux I__6560 (
            .O(N__33773),
            .I(\reset_module_System.count_1_cry_6 ));
    InMux I__6559 (
            .O(N__33770),
            .I(\reset_module_System.count_1_cry_7 ));
    InMux I__6558 (
            .O(N__33767),
            .I(bfn_14_8_0_));
    InMux I__6557 (
            .O(N__33764),
            .I(N__33761));
    LocalMux I__6556 (
            .O(N__33761),
            .I(N__33757));
    InMux I__6555 (
            .O(N__33760),
            .I(N__33754));
    Odrv4 I__6554 (
            .O(N__33757),
            .I(\reset_module_System.countZ0Z_10 ));
    LocalMux I__6553 (
            .O(N__33754),
            .I(\reset_module_System.countZ0Z_10 ));
    InMux I__6552 (
            .O(N__33749),
            .I(\reset_module_System.count_1_cry_9 ));
    CascadeMux I__6551 (
            .O(N__33746),
            .I(\pid_front.un1_reset_i_a5_1_5_cascade_ ));
    CascadeMux I__6550 (
            .O(N__33743),
            .I(N__33740));
    InMux I__6549 (
            .O(N__33740),
            .I(N__33737));
    LocalMux I__6548 (
            .O(N__33737),
            .I(N__33734));
    Odrv4 I__6547 (
            .O(N__33734),
            .I(\pid_front.un1_reset_i_a5_1_8 ));
    InMux I__6546 (
            .O(N__33731),
            .I(N__33727));
    InMux I__6545 (
            .O(N__33730),
            .I(N__33724));
    LocalMux I__6544 (
            .O(N__33727),
            .I(N__33718));
    LocalMux I__6543 (
            .O(N__33724),
            .I(N__33718));
    InMux I__6542 (
            .O(N__33723),
            .I(N__33714));
    Span4Mux_v I__6541 (
            .O(N__33718),
            .I(N__33711));
    InMux I__6540 (
            .O(N__33717),
            .I(N__33708));
    LocalMux I__6539 (
            .O(N__33714),
            .I(\pid_front.pid_preregZ0Z_10 ));
    Odrv4 I__6538 (
            .O(N__33711),
            .I(\pid_front.pid_preregZ0Z_10 ));
    LocalMux I__6537 (
            .O(N__33708),
            .I(\pid_front.pid_preregZ0Z_10 ));
    InMux I__6536 (
            .O(N__33701),
            .I(N__33698));
    LocalMux I__6535 (
            .O(N__33698),
            .I(\dron_frame_decoder_1.drone_H_disp_front_8 ));
    CascadeMux I__6534 (
            .O(N__33695),
            .I(\reset_module_System.reset6_15_cascade_ ));
    InMux I__6533 (
            .O(N__33692),
            .I(N__33689));
    LocalMux I__6532 (
            .O(N__33689),
            .I(\reset_module_System.count_1_1 ));
    CascadeMux I__6531 (
            .O(N__33686),
            .I(N__33682));
    CascadeMux I__6530 (
            .O(N__33685),
            .I(N__33675));
    InMux I__6529 (
            .O(N__33682),
            .I(N__33666));
    InMux I__6528 (
            .O(N__33681),
            .I(N__33666));
    InMux I__6527 (
            .O(N__33680),
            .I(N__33666));
    InMux I__6526 (
            .O(N__33679),
            .I(N__33666));
    InMux I__6525 (
            .O(N__33678),
            .I(N__33653));
    InMux I__6524 (
            .O(N__33675),
            .I(N__33650));
    LocalMux I__6523 (
            .O(N__33666),
            .I(N__33647));
    InMux I__6522 (
            .O(N__33665),
            .I(N__33642));
    InMux I__6521 (
            .O(N__33664),
            .I(N__33642));
    InMux I__6520 (
            .O(N__33663),
            .I(N__33639));
    InMux I__6519 (
            .O(N__33662),
            .I(N__33628));
    InMux I__6518 (
            .O(N__33661),
            .I(N__33628));
    InMux I__6517 (
            .O(N__33660),
            .I(N__33628));
    InMux I__6516 (
            .O(N__33659),
            .I(N__33628));
    InMux I__6515 (
            .O(N__33658),
            .I(N__33628));
    InMux I__6514 (
            .O(N__33657),
            .I(N__33625));
    InMux I__6513 (
            .O(N__33656),
            .I(N__33622));
    LocalMux I__6512 (
            .O(N__33653),
            .I(N__33617));
    LocalMux I__6511 (
            .O(N__33650),
            .I(N__33617));
    Sp12to4 I__6510 (
            .O(N__33647),
            .I(N__33602));
    LocalMux I__6509 (
            .O(N__33642),
            .I(N__33602));
    LocalMux I__6508 (
            .O(N__33639),
            .I(N__33602));
    LocalMux I__6507 (
            .O(N__33628),
            .I(N__33602));
    LocalMux I__6506 (
            .O(N__33625),
            .I(N__33602));
    LocalMux I__6505 (
            .O(N__33622),
            .I(N__33602));
    Sp12to4 I__6504 (
            .O(N__33617),
            .I(N__33602));
    Odrv12 I__6503 (
            .O(N__33602),
            .I(\pid_front.stateZ0Z_1 ));
    CascadeMux I__6502 (
            .O(N__33599),
            .I(N__33594));
    CascadeMux I__6501 (
            .O(N__33598),
            .I(N__33590));
    InMux I__6500 (
            .O(N__33597),
            .I(N__33575));
    InMux I__6499 (
            .O(N__33594),
            .I(N__33575));
    InMux I__6498 (
            .O(N__33593),
            .I(N__33575));
    InMux I__6497 (
            .O(N__33590),
            .I(N__33575));
    InMux I__6496 (
            .O(N__33589),
            .I(N__33575));
    InMux I__6495 (
            .O(N__33588),
            .I(N__33575));
    LocalMux I__6494 (
            .O(N__33575),
            .I(N__33569));
    InMux I__6493 (
            .O(N__33574),
            .I(N__33564));
    InMux I__6492 (
            .O(N__33573),
            .I(N__33564));
    InMux I__6491 (
            .O(N__33572),
            .I(N__33561));
    Odrv4 I__6490 (
            .O(N__33569),
            .I(\pid_front.N_287 ));
    LocalMux I__6489 (
            .O(N__33564),
            .I(\pid_front.N_287 ));
    LocalMux I__6488 (
            .O(N__33561),
            .I(\pid_front.N_287 ));
    CascadeMux I__6487 (
            .O(N__33554),
            .I(N__33550));
    InMux I__6486 (
            .O(N__33553),
            .I(N__33545));
    InMux I__6485 (
            .O(N__33550),
            .I(N__33545));
    LocalMux I__6484 (
            .O(N__33545),
            .I(\pid_front.N_533 ));
    CEMux I__6483 (
            .O(N__33542),
            .I(N__33539));
    LocalMux I__6482 (
            .O(N__33539),
            .I(N__33536));
    Odrv4 I__6481 (
            .O(N__33536),
            .I(\pid_front.state_0_1 ));
    SRMux I__6480 (
            .O(N__33533),
            .I(N__33530));
    LocalMux I__6479 (
            .O(N__33530),
            .I(N__33527));
    Span4Mux_h I__6478 (
            .O(N__33527),
            .I(N__33523));
    SRMux I__6477 (
            .O(N__33526),
            .I(N__33520));
    Span4Mux_h I__6476 (
            .O(N__33523),
            .I(N__33514));
    LocalMux I__6475 (
            .O(N__33520),
            .I(N__33514));
    SRMux I__6474 (
            .O(N__33519),
            .I(N__33511));
    Span4Mux_v I__6473 (
            .O(N__33514),
            .I(N__33507));
    LocalMux I__6472 (
            .O(N__33511),
            .I(N__33504));
    InMux I__6471 (
            .O(N__33510),
            .I(N__33501));
    Odrv4 I__6470 (
            .O(N__33507),
            .I(\pid_front.pid_prereg_RNI2A6A6Z0Z_2 ));
    Odrv12 I__6469 (
            .O(N__33504),
            .I(\pid_front.pid_prereg_RNI2A6A6Z0Z_2 ));
    LocalMux I__6468 (
            .O(N__33501),
            .I(\pid_front.pid_prereg_RNI2A6A6Z0Z_2 ));
    InMux I__6467 (
            .O(N__33494),
            .I(N__33491));
    LocalMux I__6466 (
            .O(N__33491),
            .I(\pid_front.un1_reset_i_a5_1_6 ));
    InMux I__6465 (
            .O(N__33488),
            .I(N__33485));
    LocalMux I__6464 (
            .O(N__33485),
            .I(N__33482));
    Odrv4 I__6463 (
            .O(N__33482),
            .I(\pid_front.N_315 ));
    InMux I__6462 (
            .O(N__33479),
            .I(N__33476));
    LocalMux I__6461 (
            .O(N__33476),
            .I(drone_H_disp_front_1));
    CascadeMux I__6460 (
            .O(N__33473),
            .I(\pid_side.state_ns_0_cascade_ ));
    CEMux I__6459 (
            .O(N__33470),
            .I(N__33466));
    CEMux I__6458 (
            .O(N__33469),
            .I(N__33463));
    LocalMux I__6457 (
            .O(N__33466),
            .I(N__33459));
    LocalMux I__6456 (
            .O(N__33463),
            .I(N__33456));
    CEMux I__6455 (
            .O(N__33462),
            .I(N__33453));
    Span4Mux_h I__6454 (
            .O(N__33459),
            .I(N__33450));
    Span4Mux_v I__6453 (
            .O(N__33456),
            .I(N__33447));
    LocalMux I__6452 (
            .O(N__33453),
            .I(N__33444));
    Span4Mux_v I__6451 (
            .O(N__33450),
            .I(N__33439));
    Span4Mux_h I__6450 (
            .O(N__33447),
            .I(N__33439));
    Span4Mux_v I__6449 (
            .O(N__33444),
            .I(N__33436));
    Span4Mux_h I__6448 (
            .O(N__33439),
            .I(N__33433));
    Span4Mux_v I__6447 (
            .O(N__33436),
            .I(N__33430));
    Odrv4 I__6446 (
            .O(N__33433),
            .I(\dron_frame_decoder_1.N_763_0 ));
    Odrv4 I__6445 (
            .O(N__33430),
            .I(\dron_frame_decoder_1.N_763_0 ));
    InMux I__6444 (
            .O(N__33425),
            .I(N__33422));
    LocalMux I__6443 (
            .O(N__33422),
            .I(N__33419));
    Odrv4 I__6442 (
            .O(N__33419),
            .I(\pid_front.un1_reset_i_a5_0_5 ));
    CascadeMux I__6441 (
            .O(N__33416),
            .I(\pid_front.un1_reset_i_1_cascade_ ));
    InMux I__6440 (
            .O(N__33413),
            .I(N__33409));
    InMux I__6439 (
            .O(N__33412),
            .I(N__33406));
    LocalMux I__6438 (
            .O(N__33409),
            .I(\pid_front.N_532 ));
    LocalMux I__6437 (
            .O(N__33406),
            .I(\pid_front.N_532 ));
    InMux I__6436 (
            .O(N__33401),
            .I(N__33398));
    LocalMux I__6435 (
            .O(N__33398),
            .I(\pid_front.un1_reset_i_a2_3 ));
    InMux I__6434 (
            .O(N__33395),
            .I(N__33390));
    InMux I__6433 (
            .O(N__33394),
            .I(N__33387));
    CascadeMux I__6432 (
            .O(N__33393),
            .I(N__33383));
    LocalMux I__6431 (
            .O(N__33390),
            .I(N__33378));
    LocalMux I__6430 (
            .O(N__33387),
            .I(N__33378));
    InMux I__6429 (
            .O(N__33386),
            .I(N__33374));
    InMux I__6428 (
            .O(N__33383),
            .I(N__33371));
    Span4Mux_v I__6427 (
            .O(N__33378),
            .I(N__33368));
    CascadeMux I__6426 (
            .O(N__33377),
            .I(N__33365));
    LocalMux I__6425 (
            .O(N__33374),
            .I(N__33360));
    LocalMux I__6424 (
            .O(N__33371),
            .I(N__33360));
    Span4Mux_h I__6423 (
            .O(N__33368),
            .I(N__33357));
    InMux I__6422 (
            .O(N__33365),
            .I(N__33354));
    Odrv12 I__6421 (
            .O(N__33360),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    Odrv4 I__6420 (
            .O(N__33357),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    LocalMux I__6419 (
            .O(N__33354),
            .I(\pid_alt.error_i_acumm_preregZ0Z_21 ));
    InMux I__6418 (
            .O(N__33347),
            .I(N__33343));
    CascadeMux I__6417 (
            .O(N__33346),
            .I(N__33340));
    LocalMux I__6416 (
            .O(N__33343),
            .I(N__33337));
    InMux I__6415 (
            .O(N__33340),
            .I(N__33333));
    Span12Mux_h I__6414 (
            .O(N__33337),
            .I(N__33330));
    InMux I__6413 (
            .O(N__33336),
            .I(N__33327));
    LocalMux I__6412 (
            .O(N__33333),
            .I(\pid_alt.N_557 ));
    Odrv12 I__6411 (
            .O(N__33330),
            .I(\pid_alt.N_557 ));
    LocalMux I__6410 (
            .O(N__33327),
            .I(\pid_alt.N_557 ));
    InMux I__6409 (
            .O(N__33320),
            .I(N__33315));
    InMux I__6408 (
            .O(N__33319),
            .I(N__33308));
    InMux I__6407 (
            .O(N__33318),
            .I(N__33308));
    LocalMux I__6406 (
            .O(N__33315),
            .I(N__33305));
    InMux I__6405 (
            .O(N__33314),
            .I(N__33302));
    InMux I__6404 (
            .O(N__33313),
            .I(N__33299));
    LocalMux I__6403 (
            .O(N__33308),
            .I(N__33296));
    Span12Mux_h I__6402 (
            .O(N__33305),
            .I(N__33293));
    LocalMux I__6401 (
            .O(N__33302),
            .I(N__33286));
    LocalMux I__6400 (
            .O(N__33299),
            .I(N__33286));
    Span4Mux_v I__6399 (
            .O(N__33296),
            .I(N__33286));
    Odrv12 I__6398 (
            .O(N__33293),
            .I(\pid_alt.error_i_acumm7lto13 ));
    Odrv4 I__6397 (
            .O(N__33286),
            .I(\pid_alt.error_i_acumm7lto13 ));
    InMux I__6396 (
            .O(N__33281),
            .I(N__33278));
    LocalMux I__6395 (
            .O(N__33278),
            .I(N__33275));
    Span4Mux_h I__6394 (
            .O(N__33275),
            .I(N__33272));
    Span4Mux_h I__6393 (
            .O(N__33272),
            .I(N__33269));
    Span4Mux_h I__6392 (
            .O(N__33269),
            .I(N__33266));
    Odrv4 I__6391 (
            .O(N__33266),
            .I(\pid_alt.error_i_acummZ0Z_13 ));
    CEMux I__6390 (
            .O(N__33263),
            .I(N__33260));
    LocalMux I__6389 (
            .O(N__33260),
            .I(N__33257));
    Span4Mux_h I__6388 (
            .O(N__33257),
            .I(N__33252));
    CEMux I__6387 (
            .O(N__33256),
            .I(N__33249));
    CEMux I__6386 (
            .O(N__33255),
            .I(N__33246));
    Span4Mux_h I__6385 (
            .O(N__33252),
            .I(N__33241));
    LocalMux I__6384 (
            .O(N__33249),
            .I(N__33241));
    LocalMux I__6383 (
            .O(N__33246),
            .I(N__33238));
    Span4Mux_h I__6382 (
            .O(N__33241),
            .I(N__33235));
    Span4Mux_v I__6381 (
            .O(N__33238),
            .I(N__33232));
    Odrv4 I__6380 (
            .O(N__33235),
            .I(\pid_alt.N_72_i_0 ));
    Odrv4 I__6379 (
            .O(N__33232),
            .I(\pid_alt.N_72_i_0 ));
    SRMux I__6378 (
            .O(N__33227),
            .I(N__33222));
    SRMux I__6377 (
            .O(N__33226),
            .I(N__33219));
    SRMux I__6376 (
            .O(N__33225),
            .I(N__33216));
    LocalMux I__6375 (
            .O(N__33222),
            .I(N__33213));
    LocalMux I__6374 (
            .O(N__33219),
            .I(N__33210));
    LocalMux I__6373 (
            .O(N__33216),
            .I(N__33207));
    Span4Mux_h I__6372 (
            .O(N__33213),
            .I(N__33204));
    Span4Mux_h I__6371 (
            .O(N__33210),
            .I(N__33201));
    Span4Mux_v I__6370 (
            .O(N__33207),
            .I(N__33198));
    Span4Mux_v I__6369 (
            .O(N__33204),
            .I(N__33191));
    Span4Mux_h I__6368 (
            .O(N__33201),
            .I(N__33191));
    Span4Mux_s3_h I__6367 (
            .O(N__33198),
            .I(N__33188));
    SRMux I__6366 (
            .O(N__33197),
            .I(N__33185));
    SRMux I__6365 (
            .O(N__33196),
            .I(N__33182));
    Odrv4 I__6364 (
            .O(N__33191),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ));
    Odrv4 I__6363 (
            .O(N__33188),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ));
    LocalMux I__6362 (
            .O(N__33185),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ));
    LocalMux I__6361 (
            .O(N__33182),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ));
    InMux I__6360 (
            .O(N__33173),
            .I(N__33168));
    InMux I__6359 (
            .O(N__33172),
            .I(N__33165));
    InMux I__6358 (
            .O(N__33171),
            .I(N__33162));
    LocalMux I__6357 (
            .O(N__33168),
            .I(N__33159));
    LocalMux I__6356 (
            .O(N__33165),
            .I(N__33154));
    LocalMux I__6355 (
            .O(N__33162),
            .I(N__33150));
    Span4Mux_v I__6354 (
            .O(N__33159),
            .I(N__33147));
    InMux I__6353 (
            .O(N__33158),
            .I(N__33144));
    InMux I__6352 (
            .O(N__33157),
            .I(N__33141));
    Span4Mux_v I__6351 (
            .O(N__33154),
            .I(N__33138));
    InMux I__6350 (
            .O(N__33153),
            .I(N__33135));
    Odrv4 I__6349 (
            .O(N__33150),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__6348 (
            .O(N__33147),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6347 (
            .O(N__33144),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6346 (
            .O(N__33141),
            .I(\uart_drone.stateZ0Z_4 ));
    Odrv4 I__6345 (
            .O(N__33138),
            .I(\uart_drone.stateZ0Z_4 ));
    LocalMux I__6344 (
            .O(N__33135),
            .I(\uart_drone.stateZ0Z_4 ));
    SRMux I__6343 (
            .O(N__33122),
            .I(N__33119));
    LocalMux I__6342 (
            .O(N__33119),
            .I(N__33116));
    Span4Mux_v I__6341 (
            .O(N__33116),
            .I(N__33113));
    Odrv4 I__6340 (
            .O(N__33113),
            .I(\uart_drone.state_RNIOU0NZ0Z_4 ));
    InMux I__6339 (
            .O(N__33110),
            .I(N__33107));
    LocalMux I__6338 (
            .O(N__33107),
            .I(\ppm_encoder_1.N_291 ));
    InMux I__6337 (
            .O(N__33104),
            .I(N__33101));
    LocalMux I__6336 (
            .O(N__33101),
            .I(N__33097));
    InMux I__6335 (
            .O(N__33100),
            .I(N__33092));
    Span4Mux_h I__6334 (
            .O(N__33097),
            .I(N__33088));
    InMux I__6333 (
            .O(N__33096),
            .I(N__33085));
    InMux I__6332 (
            .O(N__33095),
            .I(N__33082));
    LocalMux I__6331 (
            .O(N__33092),
            .I(N__33078));
    CascadeMux I__6330 (
            .O(N__33091),
            .I(N__33072));
    Sp12to4 I__6329 (
            .O(N__33088),
            .I(N__33065));
    LocalMux I__6328 (
            .O(N__33085),
            .I(N__33065));
    LocalMux I__6327 (
            .O(N__33082),
            .I(N__33065));
    InMux I__6326 (
            .O(N__33081),
            .I(N__33062));
    Span4Mux_h I__6325 (
            .O(N__33078),
            .I(N__33059));
    InMux I__6324 (
            .O(N__33077),
            .I(N__33054));
    InMux I__6323 (
            .O(N__33076),
            .I(N__33054));
    InMux I__6322 (
            .O(N__33075),
            .I(N__33049));
    InMux I__6321 (
            .O(N__33072),
            .I(N__33049));
    Span12Mux_v I__6320 (
            .O(N__33065),
            .I(N__33046));
    LocalMux I__6319 (
            .O(N__33062),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv4 I__6318 (
            .O(N__33059),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__6317 (
            .O(N__33054),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    LocalMux I__6316 (
            .O(N__33049),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    Odrv12 I__6315 (
            .O(N__33046),
            .I(\uart_drone.timer_CountZ0Z_4 ));
    CascadeMux I__6314 (
            .O(N__33035),
            .I(N__33032));
    InMux I__6313 (
            .O(N__33032),
            .I(N__33029));
    LocalMux I__6312 (
            .O(N__33029),
            .I(N__33024));
    InMux I__6311 (
            .O(N__33028),
            .I(N__33019));
    InMux I__6310 (
            .O(N__33027),
            .I(N__33016));
    Span4Mux_h I__6309 (
            .O(N__33024),
            .I(N__33013));
    InMux I__6308 (
            .O(N__33023),
            .I(N__33010));
    InMux I__6307 (
            .O(N__33022),
            .I(N__33007));
    LocalMux I__6306 (
            .O(N__33019),
            .I(N__32999));
    LocalMux I__6305 (
            .O(N__33016),
            .I(N__32999));
    Span4Mux_v I__6304 (
            .O(N__33013),
            .I(N__32996));
    LocalMux I__6303 (
            .O(N__33010),
            .I(N__32991));
    LocalMux I__6302 (
            .O(N__33007),
            .I(N__32991));
    InMux I__6301 (
            .O(N__33006),
            .I(N__32988));
    InMux I__6300 (
            .O(N__33005),
            .I(N__32983));
    InMux I__6299 (
            .O(N__33004),
            .I(N__32983));
    Span12Mux_v I__6298 (
            .O(N__32999),
            .I(N__32980));
    Odrv4 I__6297 (
            .O(N__32996),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv4 I__6296 (
            .O(N__32991),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__6295 (
            .O(N__32988),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    LocalMux I__6294 (
            .O(N__32983),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    Odrv12 I__6293 (
            .O(N__32980),
            .I(\uart_drone.timer_CountZ1Z_3 ));
    InMux I__6292 (
            .O(N__32969),
            .I(N__32962));
    InMux I__6291 (
            .O(N__32968),
            .I(N__32962));
    CascadeMux I__6290 (
            .O(N__32967),
            .I(N__32959));
    LocalMux I__6289 (
            .O(N__32962),
            .I(N__32955));
    InMux I__6288 (
            .O(N__32959),
            .I(N__32952));
    InMux I__6287 (
            .O(N__32958),
            .I(N__32949));
    Span12Mux_h I__6286 (
            .O(N__32955),
            .I(N__32946));
    LocalMux I__6285 (
            .O(N__32952),
            .I(N__32943));
    LocalMux I__6284 (
            .O(N__32949),
            .I(\uart_drone.stateZ0Z_2 ));
    Odrv12 I__6283 (
            .O(N__32946),
            .I(\uart_drone.stateZ0Z_2 ));
    Odrv12 I__6282 (
            .O(N__32943),
            .I(\uart_drone.stateZ0Z_2 ));
    InMux I__6281 (
            .O(N__32936),
            .I(N__32933));
    LocalMux I__6280 (
            .O(N__32933),
            .I(N__32929));
    InMux I__6279 (
            .O(N__32932),
            .I(N__32926));
    Span12Mux_s11_v I__6278 (
            .O(N__32929),
            .I(N__32923));
    LocalMux I__6277 (
            .O(N__32926),
            .I(N__32920));
    Odrv12 I__6276 (
            .O(N__32923),
            .I(\uart_drone.N_144_1 ));
    Odrv4 I__6275 (
            .O(N__32920),
            .I(\uart_drone.N_144_1 ));
    CascadeMux I__6274 (
            .O(N__32915),
            .I(\uart_drone.N_145_cascade_ ));
    InMux I__6273 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__6272 (
            .O(N__32909),
            .I(N__32904));
    InMux I__6271 (
            .O(N__32908),
            .I(N__32899));
    InMux I__6270 (
            .O(N__32907),
            .I(N__32899));
    Span4Mux_v I__6269 (
            .O(N__32904),
            .I(N__32891));
    LocalMux I__6268 (
            .O(N__32899),
            .I(N__32888));
    InMux I__6267 (
            .O(N__32898),
            .I(N__32883));
    InMux I__6266 (
            .O(N__32897),
            .I(N__32883));
    CascadeMux I__6265 (
            .O(N__32896),
            .I(N__32880));
    InMux I__6264 (
            .O(N__32895),
            .I(N__32877));
    InMux I__6263 (
            .O(N__32894),
            .I(N__32874));
    Span4Mux_v I__6262 (
            .O(N__32891),
            .I(N__32871));
    Span4Mux_v I__6261 (
            .O(N__32888),
            .I(N__32868));
    LocalMux I__6260 (
            .O(N__32883),
            .I(N__32865));
    InMux I__6259 (
            .O(N__32880),
            .I(N__32862));
    LocalMux I__6258 (
            .O(N__32877),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__6257 (
            .O(N__32874),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__6256 (
            .O(N__32871),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__6255 (
            .O(N__32868),
            .I(\uart_drone.stateZ0Z_3 ));
    Odrv4 I__6254 (
            .O(N__32865),
            .I(\uart_drone.stateZ0Z_3 ));
    LocalMux I__6253 (
            .O(N__32862),
            .I(\uart_drone.stateZ0Z_3 ));
    IoInMux I__6252 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__6251 (
            .O(N__32846),
            .I(N__32843));
    Span4Mux_s0_v I__6250 (
            .O(N__32843),
            .I(N__32838));
    InMux I__6249 (
            .O(N__32842),
            .I(N__32835));
    InMux I__6248 (
            .O(N__32841),
            .I(N__32828));
    Span4Mux_v I__6247 (
            .O(N__32838),
            .I(N__32823));
    LocalMux I__6246 (
            .O(N__32835),
            .I(N__32823));
    InMux I__6245 (
            .O(N__32834),
            .I(N__32820));
    InMux I__6244 (
            .O(N__32833),
            .I(N__32815));
    InMux I__6243 (
            .O(N__32832),
            .I(N__32815));
    InMux I__6242 (
            .O(N__32831),
            .I(N__32812));
    LocalMux I__6241 (
            .O(N__32828),
            .I(N__32809));
    Span4Mux_v I__6240 (
            .O(N__32823),
            .I(N__32806));
    LocalMux I__6239 (
            .O(N__32820),
            .I(N__32803));
    LocalMux I__6238 (
            .O(N__32815),
            .I(N__32799));
    LocalMux I__6237 (
            .O(N__32812),
            .I(N__32796));
    Span4Mux_v I__6236 (
            .O(N__32809),
            .I(N__32793));
    Span4Mux_h I__6235 (
            .O(N__32806),
            .I(N__32790));
    Span4Mux_v I__6234 (
            .O(N__32803),
            .I(N__32787));
    InMux I__6233 (
            .O(N__32802),
            .I(N__32784));
    Span4Mux_h I__6232 (
            .O(N__32799),
            .I(N__32781));
    Span4Mux_v I__6231 (
            .O(N__32796),
            .I(N__32776));
    Span4Mux_v I__6230 (
            .O(N__32793),
            .I(N__32776));
    Odrv4 I__6229 (
            .O(N__32790),
            .I(debug_CH1_0A_c));
    Odrv4 I__6228 (
            .O(N__32787),
            .I(debug_CH1_0A_c));
    LocalMux I__6227 (
            .O(N__32784),
            .I(debug_CH1_0A_c));
    Odrv4 I__6226 (
            .O(N__32781),
            .I(debug_CH1_0A_c));
    Odrv4 I__6225 (
            .O(N__32776),
            .I(debug_CH1_0A_c));
    InMux I__6224 (
            .O(N__32765),
            .I(N__32762));
    LocalMux I__6223 (
            .O(N__32762),
            .I(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ));
    InMux I__6222 (
            .O(N__32759),
            .I(N__32756));
    LocalMux I__6221 (
            .O(N__32756),
            .I(N__32753));
    Span4Mux_h I__6220 (
            .O(N__32753),
            .I(N__32749));
    InMux I__6219 (
            .O(N__32752),
            .I(N__32746));
    Odrv4 I__6218 (
            .O(N__32749),
            .I(throttle_order_12));
    LocalMux I__6217 (
            .O(N__32746),
            .I(throttle_order_12));
    InMux I__6216 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__6215 (
            .O(N__32738),
            .I(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ));
    CascadeMux I__6214 (
            .O(N__32735),
            .I(N__32730));
    InMux I__6213 (
            .O(N__32734),
            .I(N__32727));
    InMux I__6212 (
            .O(N__32733),
            .I(N__32724));
    InMux I__6211 (
            .O(N__32730),
            .I(N__32721));
    LocalMux I__6210 (
            .O(N__32727),
            .I(N__32718));
    LocalMux I__6209 (
            .O(N__32724),
            .I(N__32715));
    LocalMux I__6208 (
            .O(N__32721),
            .I(throttle_order_3));
    Odrv4 I__6207 (
            .O(N__32718),
            .I(throttle_order_3));
    Odrv4 I__6206 (
            .O(N__32715),
            .I(throttle_order_3));
    InMux I__6205 (
            .O(N__32708),
            .I(N__32705));
    LocalMux I__6204 (
            .O(N__32705),
            .I(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ));
    InMux I__6203 (
            .O(N__32702),
            .I(N__32698));
    CascadeMux I__6202 (
            .O(N__32701),
            .I(N__32695));
    LocalMux I__6201 (
            .O(N__32698),
            .I(N__32692));
    InMux I__6200 (
            .O(N__32695),
            .I(N__32689));
    Span4Mux_h I__6199 (
            .O(N__32692),
            .I(N__32686));
    LocalMux I__6198 (
            .O(N__32689),
            .I(N__32683));
    Odrv4 I__6197 (
            .O(N__32686),
            .I(throttle_order_5));
    Odrv4 I__6196 (
            .O(N__32683),
            .I(throttle_order_5));
    InMux I__6195 (
            .O(N__32678),
            .I(N__32675));
    LocalMux I__6194 (
            .O(N__32675),
            .I(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ));
    CascadeMux I__6193 (
            .O(N__32672),
            .I(N__32667));
    InMux I__6192 (
            .O(N__32671),
            .I(N__32664));
    InMux I__6191 (
            .O(N__32670),
            .I(N__32661));
    InMux I__6190 (
            .O(N__32667),
            .I(N__32658));
    LocalMux I__6189 (
            .O(N__32664),
            .I(N__32653));
    LocalMux I__6188 (
            .O(N__32661),
            .I(N__32653));
    LocalMux I__6187 (
            .O(N__32658),
            .I(N__32648));
    Span4Mux_v I__6186 (
            .O(N__32653),
            .I(N__32648));
    Odrv4 I__6185 (
            .O(N__32648),
            .I(throttle_order_6));
    CascadeMux I__6184 (
            .O(N__32645),
            .I(\ppm_encoder_1.N_314_cascade_ ));
    CascadeMux I__6183 (
            .O(N__32642),
            .I(\ppm_encoder_1.N_288_cascade_ ));
    InMux I__6182 (
            .O(N__32639),
            .I(N__32635));
    InMux I__6181 (
            .O(N__32638),
            .I(N__32632));
    LocalMux I__6180 (
            .O(N__32635),
            .I(N__32627));
    LocalMux I__6179 (
            .O(N__32632),
            .I(N__32627));
    Odrv12 I__6178 (
            .O(N__32627),
            .I(scaler_4_data_11));
    InMux I__6177 (
            .O(N__32624),
            .I(N__32621));
    LocalMux I__6176 (
            .O(N__32621),
            .I(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ));
    CascadeMux I__6175 (
            .O(N__32618),
            .I(N__32613));
    InMux I__6174 (
            .O(N__32617),
            .I(N__32610));
    InMux I__6173 (
            .O(N__32616),
            .I(N__32607));
    InMux I__6172 (
            .O(N__32613),
            .I(N__32604));
    LocalMux I__6171 (
            .O(N__32610),
            .I(N__32601));
    LocalMux I__6170 (
            .O(N__32607),
            .I(N__32598));
    LocalMux I__6169 (
            .O(N__32604),
            .I(throttle_order_11));
    Odrv4 I__6168 (
            .O(N__32601),
            .I(throttle_order_11));
    Odrv4 I__6167 (
            .O(N__32598),
            .I(throttle_order_11));
    InMux I__6166 (
            .O(N__32591),
            .I(N__32588));
    LocalMux I__6165 (
            .O(N__32588),
            .I(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ));
    InMux I__6164 (
            .O(N__32585),
            .I(N__32581));
    InMux I__6163 (
            .O(N__32584),
            .I(N__32578));
    LocalMux I__6162 (
            .O(N__32581),
            .I(N__32575));
    LocalMux I__6161 (
            .O(N__32578),
            .I(N__32572));
    Span4Mux_h I__6160 (
            .O(N__32575),
            .I(N__32569));
    Span4Mux_v I__6159 (
            .O(N__32572),
            .I(N__32566));
    Odrv4 I__6158 (
            .O(N__32569),
            .I(scaler_4_data_13));
    Odrv4 I__6157 (
            .O(N__32566),
            .I(scaler_4_data_13));
    InMux I__6156 (
            .O(N__32561),
            .I(N__32558));
    LocalMux I__6155 (
            .O(N__32558),
            .I(N__32555));
    Odrv4 I__6154 (
            .O(N__32555),
            .I(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ));
    InMux I__6153 (
            .O(N__32552),
            .I(N__32549));
    LocalMux I__6152 (
            .O(N__32549),
            .I(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ));
    CascadeMux I__6151 (
            .O(N__32546),
            .I(N__32541));
    InMux I__6150 (
            .O(N__32545),
            .I(N__32538));
    InMux I__6149 (
            .O(N__32544),
            .I(N__32535));
    InMux I__6148 (
            .O(N__32541),
            .I(N__32532));
    LocalMux I__6147 (
            .O(N__32538),
            .I(N__32529));
    LocalMux I__6146 (
            .O(N__32535),
            .I(N__32526));
    LocalMux I__6145 (
            .O(N__32532),
            .I(throttle_order_2));
    Odrv4 I__6144 (
            .O(N__32529),
            .I(throttle_order_2));
    Odrv4 I__6143 (
            .O(N__32526),
            .I(throttle_order_2));
    IoInMux I__6142 (
            .O(N__32519),
            .I(N__32516));
    LocalMux I__6141 (
            .O(N__32516),
            .I(N__32512));
    CascadeMux I__6140 (
            .O(N__32515),
            .I(N__32509));
    Span12Mux_s8_v I__6139 (
            .O(N__32512),
            .I(N__32506));
    InMux I__6138 (
            .O(N__32509),
            .I(N__32503));
    Odrv12 I__6137 (
            .O(N__32506),
            .I(ppm_output_c));
    LocalMux I__6136 (
            .O(N__32503),
            .I(ppm_output_c));
    InMux I__6135 (
            .O(N__32498),
            .I(N__32495));
    LocalMux I__6134 (
            .O(N__32495),
            .I(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ));
    CascadeMux I__6133 (
            .O(N__32492),
            .I(N__32487));
    InMux I__6132 (
            .O(N__32491),
            .I(N__32484));
    InMux I__6131 (
            .O(N__32490),
            .I(N__32481));
    InMux I__6130 (
            .O(N__32487),
            .I(N__32478));
    LocalMux I__6129 (
            .O(N__32484),
            .I(N__32473));
    LocalMux I__6128 (
            .O(N__32481),
            .I(N__32473));
    LocalMux I__6127 (
            .O(N__32478),
            .I(N__32468));
    Span4Mux_v I__6126 (
            .O(N__32473),
            .I(N__32468));
    Odrv4 I__6125 (
            .O(N__32468),
            .I(throttle_order_10));
    InMux I__6124 (
            .O(N__32465),
            .I(N__32460));
    InMux I__6123 (
            .O(N__32464),
            .I(N__32457));
    InMux I__6122 (
            .O(N__32463),
            .I(N__32454));
    LocalMux I__6121 (
            .O(N__32460),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__6120 (
            .O(N__32457),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    LocalMux I__6119 (
            .O(N__32454),
            .I(\uart_drone.timer_CountZ1Z_2 ));
    InMux I__6118 (
            .O(N__32447),
            .I(N__32444));
    LocalMux I__6117 (
            .O(N__32444),
            .I(\uart_drone.timer_Count_RNO_0_0_2 ));
    InMux I__6116 (
            .O(N__32441),
            .I(\uart_drone.un4_timer_Count_1_cry_1 ));
    InMux I__6115 (
            .O(N__32438),
            .I(N__32435));
    LocalMux I__6114 (
            .O(N__32435),
            .I(N__32432));
    Odrv4 I__6113 (
            .O(N__32432),
            .I(\uart_drone.timer_Count_RNO_0_0_3 ));
    InMux I__6112 (
            .O(N__32429),
            .I(\uart_drone.un4_timer_Count_1_cry_2 ));
    InMux I__6111 (
            .O(N__32426),
            .I(\uart_drone.un4_timer_Count_1_cry_3 ));
    InMux I__6110 (
            .O(N__32423),
            .I(N__32420));
    LocalMux I__6109 (
            .O(N__32420),
            .I(\uart_drone.timer_Count_RNO_0_0_4 ));
    CascadeMux I__6108 (
            .O(N__32417),
            .I(N__32412));
    InMux I__6107 (
            .O(N__32416),
            .I(N__32409));
    CascadeMux I__6106 (
            .O(N__32415),
            .I(N__32406));
    InMux I__6105 (
            .O(N__32412),
            .I(N__32402));
    LocalMux I__6104 (
            .O(N__32409),
            .I(N__32399));
    InMux I__6103 (
            .O(N__32406),
            .I(N__32394));
    InMux I__6102 (
            .O(N__32405),
            .I(N__32394));
    LocalMux I__6101 (
            .O(N__32402),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    Odrv12 I__6100 (
            .O(N__32399),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    LocalMux I__6099 (
            .O(N__32394),
            .I(\uart_drone.timer_Count_0_sqmuxa ));
    CascadeMux I__6098 (
            .O(N__32387),
            .I(N__32381));
    InMux I__6097 (
            .O(N__32386),
            .I(N__32378));
    InMux I__6096 (
            .O(N__32385),
            .I(N__32375));
    InMux I__6095 (
            .O(N__32384),
            .I(N__32370));
    InMux I__6094 (
            .O(N__32381),
            .I(N__32370));
    LocalMux I__6093 (
            .O(N__32378),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__6092 (
            .O(N__32375),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    LocalMux I__6091 (
            .O(N__32370),
            .I(\uart_drone.timer_CountZ0Z_0 ));
    CascadeMux I__6090 (
            .O(N__32363),
            .I(N__32358));
    InMux I__6089 (
            .O(N__32362),
            .I(N__32355));
    InMux I__6088 (
            .O(N__32361),
            .I(N__32352));
    InMux I__6087 (
            .O(N__32358),
            .I(N__32349));
    LocalMux I__6086 (
            .O(N__32355),
            .I(\uart_drone.N_126_li ));
    LocalMux I__6085 (
            .O(N__32352),
            .I(\uart_drone.N_126_li ));
    LocalMux I__6084 (
            .O(N__32349),
            .I(\uart_drone.N_126_li ));
    InMux I__6083 (
            .O(N__32342),
            .I(N__32336));
    CascadeMux I__6082 (
            .O(N__32341),
            .I(N__32331));
    CascadeMux I__6081 (
            .O(N__32340),
            .I(N__32328));
    InMux I__6080 (
            .O(N__32339),
            .I(N__32325));
    LocalMux I__6079 (
            .O(N__32336),
            .I(N__32322));
    InMux I__6078 (
            .O(N__32335),
            .I(N__32317));
    InMux I__6077 (
            .O(N__32334),
            .I(N__32317));
    InMux I__6076 (
            .O(N__32331),
            .I(N__32314));
    InMux I__6075 (
            .O(N__32328),
            .I(N__32311));
    LocalMux I__6074 (
            .O(N__32325),
            .I(\uart_drone.N_143 ));
    Odrv4 I__6073 (
            .O(N__32322),
            .I(\uart_drone.N_143 ));
    LocalMux I__6072 (
            .O(N__32317),
            .I(\uart_drone.N_143 ));
    LocalMux I__6071 (
            .O(N__32314),
            .I(\uart_drone.N_143 ));
    LocalMux I__6070 (
            .O(N__32311),
            .I(\uart_drone.N_143 ));
    InMux I__6069 (
            .O(N__32300),
            .I(N__32296));
    InMux I__6068 (
            .O(N__32299),
            .I(N__32293));
    LocalMux I__6067 (
            .O(N__32296),
            .I(N__32288));
    LocalMux I__6066 (
            .O(N__32293),
            .I(N__32288));
    Odrv12 I__6065 (
            .O(N__32288),
            .I(scaler_4_data_12));
    InMux I__6064 (
            .O(N__32285),
            .I(N__32282));
    LocalMux I__6063 (
            .O(N__32282),
            .I(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ));
    InMux I__6062 (
            .O(N__32279),
            .I(N__32276));
    LocalMux I__6061 (
            .O(N__32276),
            .I(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ));
    InMux I__6060 (
            .O(N__32273),
            .I(N__32270));
    LocalMux I__6059 (
            .O(N__32270),
            .I(N__32266));
    InMux I__6058 (
            .O(N__32269),
            .I(N__32263));
    Span4Mux_v I__6057 (
            .O(N__32266),
            .I(N__32258));
    LocalMux I__6056 (
            .O(N__32263),
            .I(N__32258));
    Odrv4 I__6055 (
            .O(N__32258),
            .I(scaler_4_data_8));
    InMux I__6054 (
            .O(N__32255),
            .I(N__32252));
    LocalMux I__6053 (
            .O(N__32252),
            .I(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ));
    InMux I__6052 (
            .O(N__32249),
            .I(N__32246));
    LocalMux I__6051 (
            .O(N__32246),
            .I(N__32242));
    InMux I__6050 (
            .O(N__32245),
            .I(N__32239));
    Span4Mux_h I__6049 (
            .O(N__32242),
            .I(N__32234));
    LocalMux I__6048 (
            .O(N__32239),
            .I(N__32234));
    Odrv4 I__6047 (
            .O(N__32234),
            .I(scaler_4_data_7));
    CascadeMux I__6046 (
            .O(N__32231),
            .I(\pid_front.un1_reset_i_a5_0_2_cascade_ ));
    InMux I__6045 (
            .O(N__32228),
            .I(N__32225));
    LocalMux I__6044 (
            .O(N__32225),
            .I(\pid_front.un1_reset_i_a5_0_3 ));
    InMux I__6043 (
            .O(N__32222),
            .I(N__32218));
    InMux I__6042 (
            .O(N__32221),
            .I(N__32213));
    LocalMux I__6041 (
            .O(N__32218),
            .I(N__32210));
    InMux I__6040 (
            .O(N__32217),
            .I(N__32207));
    InMux I__6039 (
            .O(N__32216),
            .I(N__32204));
    LocalMux I__6038 (
            .O(N__32213),
            .I(N__32201));
    Span4Mux_v I__6037 (
            .O(N__32210),
            .I(N__32196));
    LocalMux I__6036 (
            .O(N__32207),
            .I(N__32196));
    LocalMux I__6035 (
            .O(N__32204),
            .I(\pid_front.pid_preregZ0Z_1 ));
    Odrv4 I__6034 (
            .O(N__32201),
            .I(\pid_front.pid_preregZ0Z_1 ));
    Odrv4 I__6033 (
            .O(N__32196),
            .I(\pid_front.pid_preregZ0Z_1 ));
    CascadeMux I__6032 (
            .O(N__32189),
            .I(N__32185));
    InMux I__6031 (
            .O(N__32188),
            .I(N__32180));
    InMux I__6030 (
            .O(N__32185),
            .I(N__32180));
    LocalMux I__6029 (
            .O(N__32180),
            .I(N__32176));
    CascadeMux I__6028 (
            .O(N__32179),
            .I(N__32173));
    Span4Mux_h I__6027 (
            .O(N__32176),
            .I(N__32169));
    InMux I__6026 (
            .O(N__32173),
            .I(N__32166));
    InMux I__6025 (
            .O(N__32172),
            .I(N__32163));
    Odrv4 I__6024 (
            .O(N__32169),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__6023 (
            .O(N__32166),
            .I(\uart_pc.stateZ0Z_2 ));
    LocalMux I__6022 (
            .O(N__32163),
            .I(\uart_pc.stateZ0Z_2 ));
    InMux I__6021 (
            .O(N__32156),
            .I(N__32153));
    LocalMux I__6020 (
            .O(N__32153),
            .I(\uart_pc.state_srsts_i_0_2 ));
    InMux I__6019 (
            .O(N__32150),
            .I(N__32147));
    LocalMux I__6018 (
            .O(N__32147),
            .I(N__32143));
    InMux I__6017 (
            .O(N__32146),
            .I(N__32140));
    Odrv4 I__6016 (
            .O(N__32143),
            .I(\uart_pc.stateZ0Z_0 ));
    LocalMux I__6015 (
            .O(N__32140),
            .I(\uart_pc.stateZ0Z_0 ));
    CascadeMux I__6014 (
            .O(N__32135),
            .I(N__32132));
    InMux I__6013 (
            .O(N__32132),
            .I(N__32127));
    InMux I__6012 (
            .O(N__32131),
            .I(N__32122));
    InMux I__6011 (
            .O(N__32130),
            .I(N__32122));
    LocalMux I__6010 (
            .O(N__32127),
            .I(\uart_pc.stateZ0Z_1 ));
    LocalMux I__6009 (
            .O(N__32122),
            .I(\uart_pc.stateZ0Z_1 ));
    InMux I__6008 (
            .O(N__32117),
            .I(N__32113));
    InMux I__6007 (
            .O(N__32116),
            .I(N__32110));
    LocalMux I__6006 (
            .O(N__32113),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    LocalMux I__6005 (
            .O(N__32110),
            .I(\uart_drone.timer_CountZ1Z_1 ));
    CascadeMux I__6004 (
            .O(N__32105),
            .I(N__32102));
    InMux I__6003 (
            .O(N__32102),
            .I(N__32099));
    LocalMux I__6002 (
            .O(N__32099),
            .I(\uart_drone.un1_state_2_0_a3_0 ));
    InMux I__6001 (
            .O(N__32096),
            .I(N__32093));
    LocalMux I__6000 (
            .O(N__32093),
            .I(N__32089));
    CascadeMux I__5999 (
            .O(N__32092),
            .I(N__32086));
    Span4Mux_v I__5998 (
            .O(N__32089),
            .I(N__32082));
    InMux I__5997 (
            .O(N__32086),
            .I(N__32077));
    InMux I__5996 (
            .O(N__32085),
            .I(N__32077));
    Odrv4 I__5995 (
            .O(N__32082),
            .I(\uart_drone.N_152 ));
    LocalMux I__5994 (
            .O(N__32077),
            .I(\uart_drone.N_152 ));
    CascadeMux I__5993 (
            .O(N__32072),
            .I(\pid_front.N_533_cascade_ ));
    InMux I__5992 (
            .O(N__32069),
            .I(N__32057));
    InMux I__5991 (
            .O(N__32068),
            .I(N__32057));
    InMux I__5990 (
            .O(N__32067),
            .I(N__32057));
    InMux I__5989 (
            .O(N__32066),
            .I(N__32057));
    LocalMux I__5988 (
            .O(N__32057),
            .I(\pid_front.N_10_1 ));
    InMux I__5987 (
            .O(N__32054),
            .I(N__32051));
    LocalMux I__5986 (
            .O(N__32051),
            .I(N__32048));
    Span4Mux_v I__5985 (
            .O(N__32048),
            .I(N__32043));
    InMux I__5984 (
            .O(N__32047),
            .I(N__32038));
    InMux I__5983 (
            .O(N__32046),
            .I(N__32038));
    Sp12to4 I__5982 (
            .O(N__32043),
            .I(N__32033));
    LocalMux I__5981 (
            .O(N__32038),
            .I(N__32033));
    Odrv12 I__5980 (
            .O(N__32033),
            .I(\pid_alt.pid_preregZ0Z_11 ));
    InMux I__5979 (
            .O(N__32030),
            .I(N__32019));
    InMux I__5978 (
            .O(N__32029),
            .I(N__32001));
    InMux I__5977 (
            .O(N__32028),
            .I(N__32001));
    InMux I__5976 (
            .O(N__32027),
            .I(N__32001));
    InMux I__5975 (
            .O(N__32026),
            .I(N__32001));
    InMux I__5974 (
            .O(N__32025),
            .I(N__32001));
    InMux I__5973 (
            .O(N__32024),
            .I(N__32001));
    InMux I__5972 (
            .O(N__32023),
            .I(N__31998));
    InMux I__5971 (
            .O(N__32022),
            .I(N__31995));
    LocalMux I__5970 (
            .O(N__32019),
            .I(N__31992));
    InMux I__5969 (
            .O(N__32018),
            .I(N__31989));
    InMux I__5968 (
            .O(N__32017),
            .I(N__31979));
    InMux I__5967 (
            .O(N__32016),
            .I(N__31979));
    InMux I__5966 (
            .O(N__32015),
            .I(N__31979));
    InMux I__5965 (
            .O(N__32014),
            .I(N__31976));
    LocalMux I__5964 (
            .O(N__32001),
            .I(N__31971));
    LocalMux I__5963 (
            .O(N__31998),
            .I(N__31971));
    LocalMux I__5962 (
            .O(N__31995),
            .I(N__31965));
    Span4Mux_v I__5961 (
            .O(N__31992),
            .I(N__31962));
    LocalMux I__5960 (
            .O(N__31989),
            .I(N__31959));
    InMux I__5959 (
            .O(N__31988),
            .I(N__31954));
    InMux I__5958 (
            .O(N__31987),
            .I(N__31954));
    InMux I__5957 (
            .O(N__31986),
            .I(N__31951));
    LocalMux I__5956 (
            .O(N__31979),
            .I(N__31943));
    LocalMux I__5955 (
            .O(N__31976),
            .I(N__31943));
    Span4Mux_h I__5954 (
            .O(N__31971),
            .I(N__31940));
    InMux I__5953 (
            .O(N__31970),
            .I(N__31933));
    InMux I__5952 (
            .O(N__31969),
            .I(N__31933));
    InMux I__5951 (
            .O(N__31968),
            .I(N__31933));
    Span4Mux_h I__5950 (
            .O(N__31965),
            .I(N__31926));
    Span4Mux_h I__5949 (
            .O(N__31962),
            .I(N__31926));
    Span4Mux_h I__5948 (
            .O(N__31959),
            .I(N__31926));
    LocalMux I__5947 (
            .O(N__31954),
            .I(N__31923));
    LocalMux I__5946 (
            .O(N__31951),
            .I(N__31920));
    CascadeMux I__5945 (
            .O(N__31950),
            .I(N__31917));
    CascadeMux I__5944 (
            .O(N__31949),
            .I(N__31914));
    CascadeMux I__5943 (
            .O(N__31948),
            .I(N__31911));
    Span4Mux_h I__5942 (
            .O(N__31943),
            .I(N__31907));
    Span4Mux_h I__5941 (
            .O(N__31940),
            .I(N__31902));
    LocalMux I__5940 (
            .O(N__31933),
            .I(N__31902));
    Span4Mux_v I__5939 (
            .O(N__31926),
            .I(N__31899));
    Span4Mux_v I__5938 (
            .O(N__31923),
            .I(N__31896));
    Span4Mux_h I__5937 (
            .O(N__31920),
            .I(N__31893));
    InMux I__5936 (
            .O(N__31917),
            .I(N__31883));
    InMux I__5935 (
            .O(N__31914),
            .I(N__31883));
    InMux I__5934 (
            .O(N__31911),
            .I(N__31883));
    InMux I__5933 (
            .O(N__31910),
            .I(N__31883));
    Span4Mux_h I__5932 (
            .O(N__31907),
            .I(N__31880));
    Span4Mux_v I__5931 (
            .O(N__31902),
            .I(N__31877));
    Span4Mux_h I__5930 (
            .O(N__31899),
            .I(N__31870));
    Span4Mux_v I__5929 (
            .O(N__31896),
            .I(N__31870));
    Span4Mux_v I__5928 (
            .O(N__31893),
            .I(N__31870));
    InMux I__5927 (
            .O(N__31892),
            .I(N__31867));
    LocalMux I__5926 (
            .O(N__31883),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__5925 (
            .O(N__31880),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__5924 (
            .O(N__31877),
            .I(\pid_alt.N_72_i ));
    Odrv4 I__5923 (
            .O(N__31870),
            .I(\pid_alt.N_72_i ));
    LocalMux I__5922 (
            .O(N__31867),
            .I(\pid_alt.N_72_i ));
    InMux I__5921 (
            .O(N__31856),
            .I(N__31844));
    InMux I__5920 (
            .O(N__31855),
            .I(N__31844));
    InMux I__5919 (
            .O(N__31854),
            .I(N__31844));
    InMux I__5918 (
            .O(N__31853),
            .I(N__31839));
    InMux I__5917 (
            .O(N__31852),
            .I(N__31834));
    InMux I__5916 (
            .O(N__31851),
            .I(N__31834));
    LocalMux I__5915 (
            .O(N__31844),
            .I(N__31830));
    InMux I__5914 (
            .O(N__31843),
            .I(N__31825));
    InMux I__5913 (
            .O(N__31842),
            .I(N__31825));
    LocalMux I__5912 (
            .O(N__31839),
            .I(N__31820));
    LocalMux I__5911 (
            .O(N__31834),
            .I(N__31820));
    InMux I__5910 (
            .O(N__31833),
            .I(N__31817));
    Odrv4 I__5909 (
            .O(N__31830),
            .I(\pid_alt.N_299 ));
    LocalMux I__5908 (
            .O(N__31825),
            .I(\pid_alt.N_299 ));
    Odrv4 I__5907 (
            .O(N__31820),
            .I(\pid_alt.N_299 ));
    LocalMux I__5906 (
            .O(N__31817),
            .I(\pid_alt.N_299 ));
    InMux I__5905 (
            .O(N__31808),
            .I(N__31804));
    CascadeMux I__5904 (
            .O(N__31807),
            .I(N__31800));
    LocalMux I__5903 (
            .O(N__31804),
            .I(N__31797));
    InMux I__5902 (
            .O(N__31803),
            .I(N__31794));
    InMux I__5901 (
            .O(N__31800),
            .I(N__31791));
    Span4Mux_v I__5900 (
            .O(N__31797),
            .I(N__31784));
    LocalMux I__5899 (
            .O(N__31794),
            .I(N__31784));
    LocalMux I__5898 (
            .O(N__31791),
            .I(N__31784));
    Span4Mux_h I__5897 (
            .O(N__31784),
            .I(N__31781));
    Odrv4 I__5896 (
            .O(N__31781),
            .I(\pid_alt.pid_preregZ0Z_7 ));
    SRMux I__5895 (
            .O(N__31778),
            .I(N__31775));
    LocalMux I__5894 (
            .O(N__31775),
            .I(N__31771));
    SRMux I__5893 (
            .O(N__31774),
            .I(N__31765));
    Span4Mux_h I__5892 (
            .O(N__31771),
            .I(N__31762));
    SRMux I__5891 (
            .O(N__31770),
            .I(N__31759));
    SRMux I__5890 (
            .O(N__31769),
            .I(N__31756));
    InMux I__5889 (
            .O(N__31768),
            .I(N__31753));
    LocalMux I__5888 (
            .O(N__31765),
            .I(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ));
    Odrv4 I__5887 (
            .O(N__31762),
            .I(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ));
    LocalMux I__5886 (
            .O(N__31759),
            .I(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ));
    LocalMux I__5885 (
            .O(N__31756),
            .I(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ));
    LocalMux I__5884 (
            .O(N__31753),
            .I(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ));
    InMux I__5883 (
            .O(N__31742),
            .I(N__31739));
    LocalMux I__5882 (
            .O(N__31739),
            .I(N__31736));
    Odrv4 I__5881 (
            .O(N__31736),
            .I(\ppm_encoder_1.N_292 ));
    CascadeMux I__5880 (
            .O(N__31733),
            .I(\uart_drone.un1_state_7_0_cascade_ ));
    CascadeMux I__5879 (
            .O(N__31730),
            .I(\uart_drone.N_152_cascade_ ));
    InMux I__5878 (
            .O(N__31727),
            .I(N__31715));
    InMux I__5877 (
            .O(N__31726),
            .I(N__31715));
    InMux I__5876 (
            .O(N__31725),
            .I(N__31715));
    InMux I__5875 (
            .O(N__31724),
            .I(N__31715));
    LocalMux I__5874 (
            .O(N__31715),
            .I(N__31710));
    InMux I__5873 (
            .O(N__31714),
            .I(N__31707));
    InMux I__5872 (
            .O(N__31713),
            .I(N__31704));
    Span4Mux_v I__5871 (
            .O(N__31710),
            .I(N__31695));
    LocalMux I__5870 (
            .O(N__31707),
            .I(N__31695));
    LocalMux I__5869 (
            .O(N__31704),
            .I(N__31692));
    InMux I__5868 (
            .O(N__31703),
            .I(N__31689));
    InMux I__5867 (
            .O(N__31702),
            .I(N__31682));
    InMux I__5866 (
            .O(N__31701),
            .I(N__31682));
    InMux I__5865 (
            .O(N__31700),
            .I(N__31682));
    Odrv4 I__5864 (
            .O(N__31695),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    Odrv4 I__5863 (
            .O(N__31692),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__5862 (
            .O(N__31689),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    LocalMux I__5861 (
            .O(N__31682),
            .I(\uart_drone.bit_CountZ0Z_1 ));
    CascadeMux I__5860 (
            .O(N__31673),
            .I(N__31670));
    InMux I__5859 (
            .O(N__31670),
            .I(N__31667));
    LocalMux I__5858 (
            .O(N__31667),
            .I(\uart_drone.un1_state_7_0 ));
    CascadeMux I__5857 (
            .O(N__31664),
            .I(N__31658));
    CascadeMux I__5856 (
            .O(N__31663),
            .I(N__31655));
    InMux I__5855 (
            .O(N__31662),
            .I(N__31651));
    InMux I__5854 (
            .O(N__31661),
            .I(N__31642));
    InMux I__5853 (
            .O(N__31658),
            .I(N__31642));
    InMux I__5852 (
            .O(N__31655),
            .I(N__31642));
    InMux I__5851 (
            .O(N__31654),
            .I(N__31642));
    LocalMux I__5850 (
            .O(N__31651),
            .I(N__31637));
    LocalMux I__5849 (
            .O(N__31642),
            .I(N__31634));
    InMux I__5848 (
            .O(N__31641),
            .I(N__31631));
    InMux I__5847 (
            .O(N__31640),
            .I(N__31628));
    Span12Mux_v I__5846 (
            .O(N__31637),
            .I(N__31623));
    Span4Mux_h I__5845 (
            .O(N__31634),
            .I(N__31616));
    LocalMux I__5844 (
            .O(N__31631),
            .I(N__31616));
    LocalMux I__5843 (
            .O(N__31628),
            .I(N__31616));
    InMux I__5842 (
            .O(N__31627),
            .I(N__31611));
    InMux I__5841 (
            .O(N__31626),
            .I(N__31611));
    Odrv12 I__5840 (
            .O(N__31623),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    Odrv4 I__5839 (
            .O(N__31616),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    LocalMux I__5838 (
            .O(N__31611),
            .I(\uart_drone.bit_CountZ0Z_2 ));
    InMux I__5837 (
            .O(N__31604),
            .I(\ppm_encoder_1.un1_throttle_cry_12 ));
    InMux I__5836 (
            .O(N__31601),
            .I(\ppm_encoder_1.un1_throttle_cry_13 ));
    CEMux I__5835 (
            .O(N__31598),
            .I(N__31595));
    LocalMux I__5834 (
            .O(N__31595),
            .I(N__31592));
    Span4Mux_h I__5833 (
            .O(N__31592),
            .I(N__31589));
    Odrv4 I__5832 (
            .O(N__31589),
            .I(\pid_alt.N_72_i_1 ));
    InMux I__5831 (
            .O(N__31586),
            .I(N__31583));
    LocalMux I__5830 (
            .O(N__31583),
            .I(N__31580));
    Span4Mux_v I__5829 (
            .O(N__31580),
            .I(N__31577));
    Odrv4 I__5828 (
            .O(N__31577),
            .I(\uart_drone.data_Auxce_0_0_2 ));
    CascadeMux I__5827 (
            .O(N__31574),
            .I(N__31571));
    InMux I__5826 (
            .O(N__31571),
            .I(N__31567));
    InMux I__5825 (
            .O(N__31570),
            .I(N__31564));
    LocalMux I__5824 (
            .O(N__31567),
            .I(N__31560));
    LocalMux I__5823 (
            .O(N__31564),
            .I(N__31557));
    InMux I__5822 (
            .O(N__31563),
            .I(N__31554));
    Span4Mux_h I__5821 (
            .O(N__31560),
            .I(N__31551));
    Span4Mux_h I__5820 (
            .O(N__31557),
            .I(N__31546));
    LocalMux I__5819 (
            .O(N__31554),
            .I(N__31546));
    Span4Mux_h I__5818 (
            .O(N__31551),
            .I(N__31543));
    Span4Mux_h I__5817 (
            .O(N__31546),
            .I(N__31540));
    Odrv4 I__5816 (
            .O(N__31543),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    Odrv4 I__5815 (
            .O(N__31540),
            .I(\pid_alt.pid_preregZ0Z_0 ));
    CascadeMux I__5814 (
            .O(N__31535),
            .I(N__31532));
    InMux I__5813 (
            .O(N__31532),
            .I(N__31529));
    LocalMux I__5812 (
            .O(N__31529),
            .I(N__31525));
    InMux I__5811 (
            .O(N__31528),
            .I(N__31522));
    Span4Mux_v I__5810 (
            .O(N__31525),
            .I(N__31517));
    LocalMux I__5809 (
            .O(N__31522),
            .I(N__31517));
    Span4Mux_h I__5808 (
            .O(N__31517),
            .I(N__31513));
    InMux I__5807 (
            .O(N__31516),
            .I(N__31510));
    Span4Mux_h I__5806 (
            .O(N__31513),
            .I(N__31507));
    LocalMux I__5805 (
            .O(N__31510),
            .I(N__31504));
    Odrv4 I__5804 (
            .O(N__31507),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    Odrv4 I__5803 (
            .O(N__31504),
            .I(\pid_alt.pid_preregZ0Z_1 ));
    InMux I__5802 (
            .O(N__31499),
            .I(N__31496));
    LocalMux I__5801 (
            .O(N__31496),
            .I(N__31492));
    InMux I__5800 (
            .O(N__31495),
            .I(N__31489));
    Span4Mux_v I__5799 (
            .O(N__31492),
            .I(N__31484));
    LocalMux I__5798 (
            .O(N__31489),
            .I(N__31484));
    Span4Mux_h I__5797 (
            .O(N__31484),
            .I(N__31480));
    InMux I__5796 (
            .O(N__31483),
            .I(N__31477));
    Span4Mux_h I__5795 (
            .O(N__31480),
            .I(N__31474));
    LocalMux I__5794 (
            .O(N__31477),
            .I(N__31471));
    Odrv4 I__5793 (
            .O(N__31474),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    Odrv4 I__5792 (
            .O(N__31471),
            .I(\pid_alt.pid_preregZ0Z_2 ));
    InMux I__5791 (
            .O(N__31466),
            .I(N__31462));
    InMux I__5790 (
            .O(N__31465),
            .I(N__31459));
    LocalMux I__5789 (
            .O(N__31462),
            .I(N__31456));
    LocalMux I__5788 (
            .O(N__31459),
            .I(N__31453));
    Span4Mux_v I__5787 (
            .O(N__31456),
            .I(N__31450));
    Odrv12 I__5786 (
            .O(N__31453),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    Odrv4 I__5785 (
            .O(N__31450),
            .I(\pid_alt.pid_preregZ0Z_3 ));
    InMux I__5784 (
            .O(N__31445),
            .I(N__31433));
    InMux I__5783 (
            .O(N__31444),
            .I(N__31433));
    InMux I__5782 (
            .O(N__31443),
            .I(N__31433));
    InMux I__5781 (
            .O(N__31442),
            .I(N__31433));
    LocalMux I__5780 (
            .O(N__31433),
            .I(\pid_alt.N_472_1 ));
    InMux I__5779 (
            .O(N__31430),
            .I(\ppm_encoder_1.un1_throttle_cry_3 ));
    InMux I__5778 (
            .O(N__31427),
            .I(\ppm_encoder_1.un1_throttle_cry_4 ));
    InMux I__5777 (
            .O(N__31424),
            .I(\ppm_encoder_1.un1_throttle_cry_5 ));
    InMux I__5776 (
            .O(N__31421),
            .I(\ppm_encoder_1.un1_throttle_cry_6 ));
    InMux I__5775 (
            .O(N__31418),
            .I(bfn_12_13_0_));
    CascadeMux I__5774 (
            .O(N__31415),
            .I(N__31411));
    InMux I__5773 (
            .O(N__31414),
            .I(N__31408));
    InMux I__5772 (
            .O(N__31411),
            .I(N__31404));
    LocalMux I__5771 (
            .O(N__31408),
            .I(N__31401));
    InMux I__5770 (
            .O(N__31407),
            .I(N__31398));
    LocalMux I__5769 (
            .O(N__31404),
            .I(throttle_order_9));
    Odrv4 I__5768 (
            .O(N__31401),
            .I(throttle_order_9));
    LocalMux I__5767 (
            .O(N__31398),
            .I(throttle_order_9));
    InMux I__5766 (
            .O(N__31391),
            .I(N__31388));
    LocalMux I__5765 (
            .O(N__31388),
            .I(N__31385));
    Odrv4 I__5764 (
            .O(N__31385),
            .I(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ));
    InMux I__5763 (
            .O(N__31382),
            .I(\ppm_encoder_1.un1_throttle_cry_8 ));
    InMux I__5762 (
            .O(N__31379),
            .I(\ppm_encoder_1.un1_throttle_cry_9 ));
    InMux I__5761 (
            .O(N__31376),
            .I(\ppm_encoder_1.un1_throttle_cry_10 ));
    InMux I__5760 (
            .O(N__31373),
            .I(\ppm_encoder_1.un1_throttle_cry_11 ));
    InMux I__5759 (
            .O(N__31370),
            .I(\ppm_encoder_1.un1_rudder_cry_9 ));
    InMux I__5758 (
            .O(N__31367),
            .I(\ppm_encoder_1.un1_rudder_cry_10 ));
    InMux I__5757 (
            .O(N__31364),
            .I(\ppm_encoder_1.un1_rudder_cry_11 ));
    InMux I__5756 (
            .O(N__31361),
            .I(\ppm_encoder_1.un1_rudder_cry_12 ));
    InMux I__5755 (
            .O(N__31358),
            .I(N__31355));
    LocalMux I__5754 (
            .O(N__31355),
            .I(N__31352));
    Odrv4 I__5753 (
            .O(N__31352),
            .I(scaler_4_data_14));
    InMux I__5752 (
            .O(N__31349),
            .I(bfn_12_11_0_));
    InMux I__5751 (
            .O(N__31346),
            .I(\ppm_encoder_1.un1_throttle_cry_0 ));
    InMux I__5750 (
            .O(N__31343),
            .I(\ppm_encoder_1.un1_throttle_cry_1 ));
    InMux I__5749 (
            .O(N__31340),
            .I(\ppm_encoder_1.un1_throttle_cry_2 ));
    CascadeMux I__5748 (
            .O(N__31337),
            .I(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ));
    InMux I__5747 (
            .O(N__31334),
            .I(N__31329));
    InMux I__5746 (
            .O(N__31333),
            .I(N__31326));
    InMux I__5745 (
            .O(N__31332),
            .I(N__31323));
    LocalMux I__5744 (
            .O(N__31329),
            .I(N__31320));
    LocalMux I__5743 (
            .O(N__31326),
            .I(N__31317));
    LocalMux I__5742 (
            .O(N__31323),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    Odrv4 I__5741 (
            .O(N__31320),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    Odrv4 I__5740 (
            .O(N__31317),
            .I(\uart_pc.timer_CountZ1Z_2 ));
    InMux I__5739 (
            .O(N__31310),
            .I(N__31307));
    LocalMux I__5738 (
            .O(N__31307),
            .I(N__31300));
    InMux I__5737 (
            .O(N__31306),
            .I(N__31297));
    InMux I__5736 (
            .O(N__31305),
            .I(N__31294));
    InMux I__5735 (
            .O(N__31304),
            .I(N__31286));
    InMux I__5734 (
            .O(N__31303),
            .I(N__31286));
    Span4Mux_v I__5733 (
            .O(N__31300),
            .I(N__31279));
    LocalMux I__5732 (
            .O(N__31297),
            .I(N__31279));
    LocalMux I__5731 (
            .O(N__31294),
            .I(N__31279));
    InMux I__5730 (
            .O(N__31293),
            .I(N__31272));
    InMux I__5729 (
            .O(N__31292),
            .I(N__31272));
    InMux I__5728 (
            .O(N__31291),
            .I(N__31272));
    LocalMux I__5727 (
            .O(N__31286),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    Odrv4 I__5726 (
            .O(N__31279),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    LocalMux I__5725 (
            .O(N__31272),
            .I(\uart_pc.timer_CountZ1Z_3 ));
    InMux I__5724 (
            .O(N__31265),
            .I(N__31262));
    LocalMux I__5723 (
            .O(N__31262),
            .I(N__31257));
    InMux I__5722 (
            .O(N__31261),
            .I(N__31254));
    InMux I__5721 (
            .O(N__31260),
            .I(N__31251));
    Span4Mux_v I__5720 (
            .O(N__31257),
            .I(N__31246));
    LocalMux I__5719 (
            .O(N__31254),
            .I(N__31246));
    LocalMux I__5718 (
            .O(N__31251),
            .I(\uart_pc.N_126_li ));
    Odrv4 I__5717 (
            .O(N__31246),
            .I(\uart_pc.N_126_li ));
    InMux I__5716 (
            .O(N__31241),
            .I(N__31217));
    InMux I__5715 (
            .O(N__31240),
            .I(N__31217));
    InMux I__5714 (
            .O(N__31239),
            .I(N__31217));
    InMux I__5713 (
            .O(N__31238),
            .I(N__31217));
    InMux I__5712 (
            .O(N__31237),
            .I(N__31217));
    InMux I__5711 (
            .O(N__31236),
            .I(N__31217));
    InMux I__5710 (
            .O(N__31235),
            .I(N__31217));
    InMux I__5709 (
            .O(N__31234),
            .I(N__31217));
    LocalMux I__5708 (
            .O(N__31217),
            .I(N__31214));
    Odrv4 I__5707 (
            .O(N__31214),
            .I(\uart_drone.un1_state_2_0 ));
    InMux I__5706 (
            .O(N__31211),
            .I(N__31208));
    LocalMux I__5705 (
            .O(N__31208),
            .I(N__31205));
    Span4Mux_v I__5704 (
            .O(N__31205),
            .I(N__31201));
    InMux I__5703 (
            .O(N__31204),
            .I(N__31198));
    Span4Mux_v I__5702 (
            .O(N__31201),
            .I(N__31195));
    LocalMux I__5701 (
            .O(N__31198),
            .I(N__31192));
    Odrv4 I__5700 (
            .O(N__31195),
            .I(scaler_4_data_6));
    Odrv4 I__5699 (
            .O(N__31192),
            .I(scaler_4_data_6));
    InMux I__5698 (
            .O(N__31187),
            .I(\ppm_encoder_1.un1_rudder_cry_6 ));
    InMux I__5697 (
            .O(N__31184),
            .I(\ppm_encoder_1.un1_rudder_cry_7 ));
    InMux I__5696 (
            .O(N__31181),
            .I(\ppm_encoder_1.un1_rudder_cry_8 ));
    CascadeMux I__5695 (
            .O(N__31178),
            .I(N__31174));
    InMux I__5694 (
            .O(N__31177),
            .I(N__31171));
    InMux I__5693 (
            .O(N__31174),
            .I(N__31168));
    LocalMux I__5692 (
            .O(N__31171),
            .I(N__31164));
    LocalMux I__5691 (
            .O(N__31168),
            .I(N__31160));
    InMux I__5690 (
            .O(N__31167),
            .I(N__31157));
    Span4Mux_v I__5689 (
            .O(N__31164),
            .I(N__31154));
    InMux I__5688 (
            .O(N__31163),
            .I(N__31151));
    Span4Mux_v I__5687 (
            .O(N__31160),
            .I(N__31148));
    LocalMux I__5686 (
            .O(N__31157),
            .I(N__31144));
    Sp12to4 I__5685 (
            .O(N__31154),
            .I(N__31139));
    LocalMux I__5684 (
            .O(N__31151),
            .I(N__31139));
    Span4Mux_v I__5683 (
            .O(N__31148),
            .I(N__31136));
    InMux I__5682 (
            .O(N__31147),
            .I(N__31133));
    Sp12to4 I__5681 (
            .O(N__31144),
            .I(N__31128));
    Span12Mux_h I__5680 (
            .O(N__31139),
            .I(N__31128));
    Span4Mux_v I__5679 (
            .O(N__31136),
            .I(N__31125));
    LocalMux I__5678 (
            .O(N__31133),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv12 I__5677 (
            .O(N__31128),
            .I(\pid_alt.stateZ0Z_0 ));
    Odrv4 I__5676 (
            .O(N__31125),
            .I(\pid_alt.stateZ0Z_0 ));
    IoInMux I__5675 (
            .O(N__31118),
            .I(N__31115));
    LocalMux I__5674 (
            .O(N__31115),
            .I(\pid_alt.state_0_0 ));
    CascadeMux I__5673 (
            .O(N__31112),
            .I(N__31105));
    CascadeMux I__5672 (
            .O(N__31111),
            .I(N__31102));
    CascadeMux I__5671 (
            .O(N__31110),
            .I(N__31095));
    CascadeMux I__5670 (
            .O(N__31109),
            .I(N__31092));
    InMux I__5669 (
            .O(N__31108),
            .I(N__31085));
    InMux I__5668 (
            .O(N__31105),
            .I(N__31085));
    InMux I__5667 (
            .O(N__31102),
            .I(N__31085));
    InMux I__5666 (
            .O(N__31101),
            .I(N__31082));
    InMux I__5665 (
            .O(N__31100),
            .I(N__31079));
    InMux I__5664 (
            .O(N__31099),
            .I(N__31074));
    InMux I__5663 (
            .O(N__31098),
            .I(N__31074));
    InMux I__5662 (
            .O(N__31095),
            .I(N__31069));
    InMux I__5661 (
            .O(N__31092),
            .I(N__31069));
    LocalMux I__5660 (
            .O(N__31085),
            .I(N__31066));
    LocalMux I__5659 (
            .O(N__31082),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__5658 (
            .O(N__31079),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__5657 (
            .O(N__31074),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    LocalMux I__5656 (
            .O(N__31069),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    Odrv4 I__5655 (
            .O(N__31066),
            .I(\uart_pc.timer_CountZ0Z_4 ));
    IoInMux I__5654 (
            .O(N__31055),
            .I(N__31051));
    InMux I__5653 (
            .O(N__31054),
            .I(N__31043));
    LocalMux I__5652 (
            .O(N__31051),
            .I(N__31039));
    CascadeMux I__5651 (
            .O(N__31050),
            .I(N__31036));
    CascadeMux I__5650 (
            .O(N__31049),
            .I(N__31033));
    CascadeMux I__5649 (
            .O(N__31048),
            .I(N__31030));
    CascadeMux I__5648 (
            .O(N__31047),
            .I(N__31027));
    CascadeMux I__5647 (
            .O(N__31046),
            .I(N__31022));
    LocalMux I__5646 (
            .O(N__31043),
            .I(N__31018));
    InMux I__5645 (
            .O(N__31042),
            .I(N__31015));
    Span4Mux_s3_v I__5644 (
            .O(N__31039),
            .I(N__31012));
    InMux I__5643 (
            .O(N__31036),
            .I(N__30996));
    InMux I__5642 (
            .O(N__31033),
            .I(N__30996));
    InMux I__5641 (
            .O(N__31030),
            .I(N__30996));
    InMux I__5640 (
            .O(N__31027),
            .I(N__30996));
    InMux I__5639 (
            .O(N__31026),
            .I(N__30996));
    InMux I__5638 (
            .O(N__31025),
            .I(N__30996));
    InMux I__5637 (
            .O(N__31022),
            .I(N__30991));
    InMux I__5636 (
            .O(N__31021),
            .I(N__30991));
    Span4Mux_v I__5635 (
            .O(N__31018),
            .I(N__30986));
    LocalMux I__5634 (
            .O(N__31015),
            .I(N__30986));
    Span4Mux_v I__5633 (
            .O(N__31012),
            .I(N__30983));
    InMux I__5632 (
            .O(N__31011),
            .I(N__30980));
    InMux I__5631 (
            .O(N__31010),
            .I(N__30975));
    InMux I__5630 (
            .O(N__31009),
            .I(N__30975));
    LocalMux I__5629 (
            .O(N__30996),
            .I(N__30970));
    LocalMux I__5628 (
            .O(N__30991),
            .I(N__30970));
    Span4Mux_v I__5627 (
            .O(N__30986),
            .I(N__30967));
    Odrv4 I__5626 (
            .O(N__30983),
            .I(debug_CH0_16A_c));
    LocalMux I__5625 (
            .O(N__30980),
            .I(debug_CH0_16A_c));
    LocalMux I__5624 (
            .O(N__30975),
            .I(debug_CH0_16A_c));
    Odrv12 I__5623 (
            .O(N__30970),
            .I(debug_CH0_16A_c));
    Odrv4 I__5622 (
            .O(N__30967),
            .I(debug_CH0_16A_c));
    CascadeMux I__5621 (
            .O(N__30956),
            .I(\uart_drone.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__5620 (
            .O(N__30953),
            .I(N__30950));
    InMux I__5619 (
            .O(N__30950),
            .I(N__30947));
    LocalMux I__5618 (
            .O(N__30947),
            .I(N__30944));
    Span4Mux_h I__5617 (
            .O(N__30944),
            .I(N__30940));
    InMux I__5616 (
            .O(N__30943),
            .I(N__30937));
    Odrv4 I__5615 (
            .O(N__30940),
            .I(\uart_drone.stateZ0Z_0 ));
    LocalMux I__5614 (
            .O(N__30937),
            .I(\uart_drone.stateZ0Z_0 ));
    InMux I__5613 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__5612 (
            .O(N__30929),
            .I(N__30926));
    Odrv12 I__5611 (
            .O(N__30926),
            .I(\pid_side.un1_pid_prereg_cry_2_THRU_CO ));
    InMux I__5610 (
            .O(N__30923),
            .I(N__30919));
    InMux I__5609 (
            .O(N__30922),
            .I(N__30916));
    LocalMux I__5608 (
            .O(N__30919),
            .I(N__30913));
    LocalMux I__5607 (
            .O(N__30916),
            .I(N__30910));
    Span4Mux_v I__5606 (
            .O(N__30913),
            .I(N__30906));
    Span4Mux_v I__5605 (
            .O(N__30910),
            .I(N__30903));
    InMux I__5604 (
            .O(N__30909),
            .I(N__30900));
    Sp12to4 I__5603 (
            .O(N__30906),
            .I(N__30895));
    Sp12to4 I__5602 (
            .O(N__30903),
            .I(N__30895));
    LocalMux I__5601 (
            .O(N__30900),
            .I(\pid_side.error_p_regZ0Z_16 ));
    Odrv12 I__5600 (
            .O(N__30895),
            .I(\pid_side.error_p_regZ0Z_16 ));
    InMux I__5599 (
            .O(N__30890),
            .I(N__30887));
    LocalMux I__5598 (
            .O(N__30887),
            .I(N__30884));
    Span4Mux_h I__5597 (
            .O(N__30884),
            .I(N__30881));
    Odrv4 I__5596 (
            .O(N__30881),
            .I(\pid_side.un1_pid_prereg_cry_15_THRU_CO ));
    InMux I__5595 (
            .O(N__30878),
            .I(N__30875));
    LocalMux I__5594 (
            .O(N__30875),
            .I(N__30872));
    Odrv12 I__5593 (
            .O(N__30872),
            .I(\pid_side.un1_pid_prereg_cry_4_THRU_CO ));
    InMux I__5592 (
            .O(N__30869),
            .I(N__30866));
    LocalMux I__5591 (
            .O(N__30866),
            .I(N__30862));
    InMux I__5590 (
            .O(N__30865),
            .I(N__30859));
    Span4Mux_h I__5589 (
            .O(N__30862),
            .I(N__30854));
    LocalMux I__5588 (
            .O(N__30859),
            .I(N__30854));
    Span4Mux_h I__5587 (
            .O(N__30854),
            .I(N__30850));
    InMux I__5586 (
            .O(N__30853),
            .I(N__30847));
    Span4Mux_h I__5585 (
            .O(N__30850),
            .I(N__30844));
    LocalMux I__5584 (
            .O(N__30847),
            .I(\pid_side.error_p_regZ0Z_5 ));
    Odrv4 I__5583 (
            .O(N__30844),
            .I(\pid_side.error_p_regZ0Z_5 ));
    InMux I__5582 (
            .O(N__30839),
            .I(N__30836));
    LocalMux I__5581 (
            .O(N__30836),
            .I(N__30833));
    Span4Mux_v I__5580 (
            .O(N__30833),
            .I(N__30829));
    InMux I__5579 (
            .O(N__30832),
            .I(N__30826));
    Sp12to4 I__5578 (
            .O(N__30829),
            .I(N__30820));
    LocalMux I__5577 (
            .O(N__30826),
            .I(N__30820));
    InMux I__5576 (
            .O(N__30825),
            .I(N__30817));
    Span12Mux_h I__5575 (
            .O(N__30820),
            .I(N__30814));
    LocalMux I__5574 (
            .O(N__30817),
            .I(\pid_side.error_p_regZ0Z_13 ));
    Odrv12 I__5573 (
            .O(N__30814),
            .I(\pid_side.error_p_regZ0Z_13 ));
    InMux I__5572 (
            .O(N__30809),
            .I(N__30806));
    LocalMux I__5571 (
            .O(N__30806),
            .I(N__30803));
    Span4Mux_h I__5570 (
            .O(N__30803),
            .I(N__30800));
    Odrv4 I__5569 (
            .O(N__30800),
            .I(\pid_side.un1_pid_prereg_cry_12_THRU_CO ));
    InMux I__5568 (
            .O(N__30797),
            .I(N__30793));
    InMux I__5567 (
            .O(N__30796),
            .I(N__30790));
    LocalMux I__5566 (
            .O(N__30793),
            .I(N__30787));
    LocalMux I__5565 (
            .O(N__30790),
            .I(N__30784));
    Span4Mux_v I__5564 (
            .O(N__30787),
            .I(N__30781));
    Span4Mux_v I__5563 (
            .O(N__30784),
            .I(N__30778));
    Span4Mux_v I__5562 (
            .O(N__30781),
            .I(N__30775));
    Span4Mux_h I__5561 (
            .O(N__30778),
            .I(N__30772));
    Span4Mux_h I__5560 (
            .O(N__30775),
            .I(N__30769));
    Span4Mux_h I__5559 (
            .O(N__30772),
            .I(N__30766));
    Span4Mux_h I__5558 (
            .O(N__30769),
            .I(N__30761));
    Span4Mux_h I__5557 (
            .O(N__30766),
            .I(N__30761));
    Odrv4 I__5556 (
            .O(N__30761),
            .I(xy_kp_1));
    InMux I__5555 (
            .O(N__30758),
            .I(N__30754));
    InMux I__5554 (
            .O(N__30757),
            .I(N__30751));
    LocalMux I__5553 (
            .O(N__30754),
            .I(N__30748));
    LocalMux I__5552 (
            .O(N__30751),
            .I(N__30745));
    Span4Mux_h I__5551 (
            .O(N__30748),
            .I(N__30742));
    Span4Mux_s1_h I__5550 (
            .O(N__30745),
            .I(N__30739));
    Span4Mux_v I__5549 (
            .O(N__30742),
            .I(N__30736));
    Span4Mux_h I__5548 (
            .O(N__30739),
            .I(N__30733));
    Span4Mux_h I__5547 (
            .O(N__30736),
            .I(N__30730));
    Span4Mux_h I__5546 (
            .O(N__30733),
            .I(N__30727));
    Span4Mux_h I__5545 (
            .O(N__30730),
            .I(N__30722));
    Span4Mux_h I__5544 (
            .O(N__30727),
            .I(N__30722));
    Odrv4 I__5543 (
            .O(N__30722),
            .I(xy_kp_7));
    InMux I__5542 (
            .O(N__30719),
            .I(N__30716));
    LocalMux I__5541 (
            .O(N__30716),
            .I(\pid_alt.un1_reset_i_a5_1_10_8 ));
    InMux I__5540 (
            .O(N__30713),
            .I(N__30710));
    LocalMux I__5539 (
            .O(N__30710),
            .I(N__30707));
    Odrv12 I__5538 (
            .O(N__30707),
            .I(\pid_alt.un1_reset_i_a5_1_10_9 ));
    CascadeMux I__5537 (
            .O(N__30704),
            .I(\pid_alt.un1_reset_i_a5_0_6_cascade_ ));
    CascadeMux I__5536 (
            .O(N__30701),
            .I(\pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_ ));
    InMux I__5535 (
            .O(N__30698),
            .I(N__30695));
    LocalMux I__5534 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_h I__5533 (
            .O(N__30692),
            .I(N__30689));
    Odrv4 I__5532 (
            .O(N__30689),
            .I(\uart_drone.data_Auxce_0_5 ));
    InMux I__5531 (
            .O(N__30686),
            .I(N__30682));
    InMux I__5530 (
            .O(N__30685),
            .I(N__30679));
    LocalMux I__5529 (
            .O(N__30682),
            .I(\pid_alt.N_530 ));
    LocalMux I__5528 (
            .O(N__30679),
            .I(\pid_alt.N_530 ));
    CascadeMux I__5527 (
            .O(N__30674),
            .I(N__30671));
    InMux I__5526 (
            .O(N__30671),
            .I(N__30665));
    InMux I__5525 (
            .O(N__30670),
            .I(N__30665));
    LocalMux I__5524 (
            .O(N__30665),
            .I(N__30662));
    Odrv4 I__5523 (
            .O(N__30662),
            .I(\pid_alt.N_535 ));
    InMux I__5522 (
            .O(N__30659),
            .I(N__30652));
    InMux I__5521 (
            .O(N__30658),
            .I(N__30652));
    InMux I__5520 (
            .O(N__30657),
            .I(N__30649));
    LocalMux I__5519 (
            .O(N__30652),
            .I(N__30645));
    LocalMux I__5518 (
            .O(N__30649),
            .I(N__30642));
    CascadeMux I__5517 (
            .O(N__30648),
            .I(N__30639));
    Span4Mux_v I__5516 (
            .O(N__30645),
            .I(N__30633));
    Span4Mux_v I__5515 (
            .O(N__30642),
            .I(N__30633));
    InMux I__5514 (
            .O(N__30639),
            .I(N__30630));
    InMux I__5513 (
            .O(N__30638),
            .I(N__30627));
    Sp12to4 I__5512 (
            .O(N__30633),
            .I(N__30620));
    LocalMux I__5511 (
            .O(N__30630),
            .I(N__30620));
    LocalMux I__5510 (
            .O(N__30627),
            .I(N__30620));
    Odrv12 I__5509 (
            .O(N__30620),
            .I(\pid_alt.pid_preregZ0Z_5 ));
    CascadeMux I__5508 (
            .O(N__30617),
            .I(\pid_alt.N_535_cascade_ ));
    CascadeMux I__5507 (
            .O(N__30614),
            .I(N__30611));
    InMux I__5506 (
            .O(N__30611),
            .I(N__30606));
    InMux I__5505 (
            .O(N__30610),
            .I(N__30603));
    InMux I__5504 (
            .O(N__30609),
            .I(N__30600));
    LocalMux I__5503 (
            .O(N__30606),
            .I(N__30597));
    LocalMux I__5502 (
            .O(N__30603),
            .I(N__30594));
    LocalMux I__5501 (
            .O(N__30600),
            .I(N__30591));
    Span4Mux_h I__5500 (
            .O(N__30597),
            .I(N__30587));
    Span4Mux_v I__5499 (
            .O(N__30594),
            .I(N__30584));
    Span4Mux_v I__5498 (
            .O(N__30591),
            .I(N__30581));
    InMux I__5497 (
            .O(N__30590),
            .I(N__30578));
    Span4Mux_h I__5496 (
            .O(N__30587),
            .I(N__30575));
    Span4Mux_h I__5495 (
            .O(N__30584),
            .I(N__30572));
    Span4Mux_h I__5494 (
            .O(N__30581),
            .I(N__30567));
    LocalMux I__5493 (
            .O(N__30578),
            .I(N__30567));
    Odrv4 I__5492 (
            .O(N__30575),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    Odrv4 I__5491 (
            .O(N__30572),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    Odrv4 I__5490 (
            .O(N__30567),
            .I(\pid_alt.pid_preregZ0Z_4 ));
    InMux I__5489 (
            .O(N__30560),
            .I(N__30557));
    LocalMux I__5488 (
            .O(N__30557),
            .I(N__30554));
    Span4Mux_v I__5487 (
            .O(N__30554),
            .I(N__30551));
    Odrv4 I__5486 (
            .O(N__30551),
            .I(\uart_drone.data_Auxce_0_6 ));
    InMux I__5485 (
            .O(N__30548),
            .I(N__30544));
    InMux I__5484 (
            .O(N__30547),
            .I(N__30540));
    LocalMux I__5483 (
            .O(N__30544),
            .I(N__30537));
    CascadeMux I__5482 (
            .O(N__30543),
            .I(N__30533));
    LocalMux I__5481 (
            .O(N__30540),
            .I(N__30530));
    Span4Mux_v I__5480 (
            .O(N__30537),
            .I(N__30527));
    InMux I__5479 (
            .O(N__30536),
            .I(N__30524));
    InMux I__5478 (
            .O(N__30533),
            .I(N__30521));
    Span4Mux_h I__5477 (
            .O(N__30530),
            .I(N__30518));
    Sp12to4 I__5476 (
            .O(N__30527),
            .I(N__30511));
    LocalMux I__5475 (
            .O(N__30524),
            .I(N__30511));
    LocalMux I__5474 (
            .O(N__30521),
            .I(N__30511));
    Odrv4 I__5473 (
            .O(N__30518),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    Odrv12 I__5472 (
            .O(N__30511),
            .I(\pid_alt.pid_preregZ0Z_12 ));
    InMux I__5471 (
            .O(N__30506),
            .I(N__30500));
    InMux I__5470 (
            .O(N__30505),
            .I(N__30500));
    LocalMux I__5469 (
            .O(N__30500),
            .I(N__30496));
    InMux I__5468 (
            .O(N__30499),
            .I(N__30493));
    Span4Mux_v I__5467 (
            .O(N__30496),
            .I(N__30485));
    LocalMux I__5466 (
            .O(N__30493),
            .I(N__30485));
    InMux I__5465 (
            .O(N__30492),
            .I(N__30480));
    InMux I__5464 (
            .O(N__30491),
            .I(N__30480));
    InMux I__5463 (
            .O(N__30490),
            .I(N__30477));
    Span4Mux_h I__5462 (
            .O(N__30485),
            .I(N__30474));
    LocalMux I__5461 (
            .O(N__30480),
            .I(N__30469));
    LocalMux I__5460 (
            .O(N__30477),
            .I(N__30469));
    Span4Mux_h I__5459 (
            .O(N__30474),
            .I(N__30466));
    Odrv12 I__5458 (
            .O(N__30469),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    Odrv4 I__5457 (
            .O(N__30466),
            .I(\pid_alt.pid_preregZ0Z_13 ));
    CascadeMux I__5456 (
            .O(N__30461),
            .I(N__30455));
    CascadeMux I__5455 (
            .O(N__30460),
            .I(N__30452));
    InMux I__5454 (
            .O(N__30459),
            .I(N__30448));
    InMux I__5453 (
            .O(N__30458),
            .I(N__30443));
    InMux I__5452 (
            .O(N__30455),
            .I(N__30443));
    InMux I__5451 (
            .O(N__30452),
            .I(N__30438));
    InMux I__5450 (
            .O(N__30451),
            .I(N__30438));
    LocalMux I__5449 (
            .O(N__30448),
            .I(N__30435));
    LocalMux I__5448 (
            .O(N__30443),
            .I(N__30432));
    LocalMux I__5447 (
            .O(N__30438),
            .I(N__30429));
    Span4Mux_v I__5446 (
            .O(N__30435),
            .I(N__30426));
    Span4Mux_v I__5445 (
            .O(N__30432),
            .I(N__30423));
    Span12Mux_v I__5444 (
            .O(N__30429),
            .I(N__30420));
    Span4Mux_h I__5443 (
            .O(N__30426),
            .I(N__30415));
    Span4Mux_h I__5442 (
            .O(N__30423),
            .I(N__30415));
    Odrv12 I__5441 (
            .O(N__30420),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    Odrv4 I__5440 (
            .O(N__30415),
            .I(\pid_alt.pid_preregZ0Z_24 ));
    InMux I__5439 (
            .O(N__30410),
            .I(N__30403));
    InMux I__5438 (
            .O(N__30409),
            .I(N__30403));
    InMux I__5437 (
            .O(N__30408),
            .I(N__30400));
    LocalMux I__5436 (
            .O(N__30403),
            .I(N__30396));
    LocalMux I__5435 (
            .O(N__30400),
            .I(N__30393));
    InMux I__5434 (
            .O(N__30399),
            .I(N__30390));
    Span4Mux_v I__5433 (
            .O(N__30396),
            .I(N__30383));
    Span4Mux_v I__5432 (
            .O(N__30393),
            .I(N__30383));
    LocalMux I__5431 (
            .O(N__30390),
            .I(N__30383));
    Span4Mux_h I__5430 (
            .O(N__30383),
            .I(N__30380));
    Odrv4 I__5429 (
            .O(N__30380),
            .I(\pid_alt.N_551 ));
    InMux I__5428 (
            .O(N__30377),
            .I(N__30374));
    LocalMux I__5427 (
            .O(N__30374),
            .I(N__30371));
    Odrv12 I__5426 (
            .O(N__30371),
            .I(\pid_side.un1_pid_prereg_cry_6_THRU_CO ));
    InMux I__5425 (
            .O(N__30368),
            .I(N__30365));
    LocalMux I__5424 (
            .O(N__30365),
            .I(N__30362));
    Span4Mux_v I__5423 (
            .O(N__30362),
            .I(N__30358));
    InMux I__5422 (
            .O(N__30361),
            .I(N__30355));
    Span4Mux_h I__5421 (
            .O(N__30358),
            .I(N__30349));
    LocalMux I__5420 (
            .O(N__30355),
            .I(N__30349));
    InMux I__5419 (
            .O(N__30354),
            .I(N__30346));
    Span4Mux_v I__5418 (
            .O(N__30349),
            .I(N__30343));
    LocalMux I__5417 (
            .O(N__30346),
            .I(N__30338));
    Span4Mux_h I__5416 (
            .O(N__30343),
            .I(N__30338));
    Odrv4 I__5415 (
            .O(N__30338),
            .I(\pid_side.error_p_regZ0Z_7 ));
    InMux I__5414 (
            .O(N__30335),
            .I(N__30332));
    LocalMux I__5413 (
            .O(N__30332),
            .I(N__30329));
    Odrv4 I__5412 (
            .O(N__30329),
            .I(\uart_drone.data_Auxce_0_1 ));
    InMux I__5411 (
            .O(N__30326),
            .I(N__30323));
    LocalMux I__5410 (
            .O(N__30323),
            .I(\uart_drone.data_Auxce_0_3 ));
    InMux I__5409 (
            .O(N__30320),
            .I(N__30317));
    LocalMux I__5408 (
            .O(N__30317),
            .I(\uart_drone.data_Auxce_0_0_4 ));
    InMux I__5407 (
            .O(N__30314),
            .I(N__30311));
    LocalMux I__5406 (
            .O(N__30311),
            .I(\pid_alt.un1_reset_i_a5_0_6_3 ));
    InMux I__5405 (
            .O(N__30308),
            .I(N__30305));
    LocalMux I__5404 (
            .O(N__30305),
            .I(N__30302));
    Span4Mux_v I__5403 (
            .O(N__30302),
            .I(N__30299));
    Span4Mux_h I__5402 (
            .O(N__30299),
            .I(N__30295));
    InMux I__5401 (
            .O(N__30298),
            .I(N__30292));
    Span4Mux_v I__5400 (
            .O(N__30295),
            .I(N__30287));
    LocalMux I__5399 (
            .O(N__30292),
            .I(N__30287));
    Span4Mux_v I__5398 (
            .O(N__30287),
            .I(N__30284));
    Span4Mux_h I__5397 (
            .O(N__30284),
            .I(N__30281));
    Odrv4 I__5396 (
            .O(N__30281),
            .I(\pid_alt.N_306_5 ));
    CascadeMux I__5395 (
            .O(N__30278),
            .I(\pid_alt.un1_reset_i_a5_0_6_2_cascade_ ));
    InMux I__5394 (
            .O(N__30275),
            .I(N__30271));
    InMux I__5393 (
            .O(N__30274),
            .I(N__30268));
    LocalMux I__5392 (
            .O(N__30271),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    LocalMux I__5391 (
            .O(N__30268),
            .I(\uart_drone.data_AuxZ0Z_1 ));
    CascadeMux I__5390 (
            .O(N__30263),
            .I(N__30259));
    InMux I__5389 (
            .O(N__30262),
            .I(N__30256));
    InMux I__5388 (
            .O(N__30259),
            .I(N__30253));
    LocalMux I__5387 (
            .O(N__30256),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    LocalMux I__5386 (
            .O(N__30253),
            .I(\uart_drone.data_AuxZ0Z_2 ));
    InMux I__5385 (
            .O(N__30248),
            .I(N__30244));
    InMux I__5384 (
            .O(N__30247),
            .I(N__30241));
    LocalMux I__5383 (
            .O(N__30244),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    LocalMux I__5382 (
            .O(N__30241),
            .I(\uart_drone.data_AuxZ0Z_3 ));
    InMux I__5381 (
            .O(N__30236),
            .I(N__30232));
    InMux I__5380 (
            .O(N__30235),
            .I(N__30229));
    LocalMux I__5379 (
            .O(N__30232),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    LocalMux I__5378 (
            .O(N__30229),
            .I(\uart_drone.data_AuxZ0Z_4 ));
    InMux I__5377 (
            .O(N__30224),
            .I(N__30220));
    InMux I__5376 (
            .O(N__30223),
            .I(N__30217));
    LocalMux I__5375 (
            .O(N__30220),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    LocalMux I__5374 (
            .O(N__30217),
            .I(\uart_drone.data_AuxZ0Z_5 ));
    CascadeMux I__5373 (
            .O(N__30212),
            .I(N__30208));
    InMux I__5372 (
            .O(N__30211),
            .I(N__30205));
    InMux I__5371 (
            .O(N__30208),
            .I(N__30202));
    LocalMux I__5370 (
            .O(N__30205),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    LocalMux I__5369 (
            .O(N__30202),
            .I(\uart_drone.data_AuxZ0Z_6 ));
    InMux I__5368 (
            .O(N__30197),
            .I(N__30193));
    InMux I__5367 (
            .O(N__30196),
            .I(N__30190));
    LocalMux I__5366 (
            .O(N__30193),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    LocalMux I__5365 (
            .O(N__30190),
            .I(\uart_drone.data_AuxZ0Z_7 ));
    InMux I__5364 (
            .O(N__30185),
            .I(N__30182));
    LocalMux I__5363 (
            .O(N__30182),
            .I(N__30177));
    InMux I__5362 (
            .O(N__30181),
            .I(N__30172));
    InMux I__5361 (
            .O(N__30180),
            .I(N__30172));
    Span4Mux_v I__5360 (
            .O(N__30177),
            .I(N__30167));
    LocalMux I__5359 (
            .O(N__30172),
            .I(N__30167));
    Span4Mux_h I__5358 (
            .O(N__30167),
            .I(N__30164));
    Odrv4 I__5357 (
            .O(N__30164),
            .I(\pid_alt.pid_preregZ0Z_9 ));
    InMux I__5356 (
            .O(N__30161),
            .I(N__30158));
    LocalMux I__5355 (
            .O(N__30158),
            .I(\uart_drone.data_Auxce_0_0_0 ));
    CascadeMux I__5354 (
            .O(N__30155),
            .I(\uart_pc.N_152_cascade_ ));
    CascadeMux I__5353 (
            .O(N__30152),
            .I(N__30148));
    InMux I__5352 (
            .O(N__30151),
            .I(N__30145));
    InMux I__5351 (
            .O(N__30148),
            .I(N__30141));
    LocalMux I__5350 (
            .O(N__30145),
            .I(N__30133));
    InMux I__5349 (
            .O(N__30144),
            .I(N__30130));
    LocalMux I__5348 (
            .O(N__30141),
            .I(N__30127));
    InMux I__5347 (
            .O(N__30140),
            .I(N__30124));
    InMux I__5346 (
            .O(N__30139),
            .I(N__30121));
    InMux I__5345 (
            .O(N__30138),
            .I(N__30114));
    InMux I__5344 (
            .O(N__30137),
            .I(N__30114));
    InMux I__5343 (
            .O(N__30136),
            .I(N__30114));
    Odrv4 I__5342 (
            .O(N__30133),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__5341 (
            .O(N__30130),
            .I(\uart_pc.stateZ0Z_3 ));
    Odrv4 I__5340 (
            .O(N__30127),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__5339 (
            .O(N__30124),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__5338 (
            .O(N__30121),
            .I(\uart_pc.stateZ0Z_3 ));
    LocalMux I__5337 (
            .O(N__30114),
            .I(\uart_pc.stateZ0Z_3 ));
    CascadeMux I__5336 (
            .O(N__30101),
            .I(\uart_pc.CO0_cascade_ ));
    InMux I__5335 (
            .O(N__30098),
            .I(N__30089));
    InMux I__5334 (
            .O(N__30097),
            .I(N__30089));
    InMux I__5333 (
            .O(N__30096),
            .I(N__30089));
    LocalMux I__5332 (
            .O(N__30089),
            .I(N__30085));
    InMux I__5331 (
            .O(N__30088),
            .I(N__30082));
    Odrv4 I__5330 (
            .O(N__30085),
            .I(\uart_pc.un1_state_4_0 ));
    LocalMux I__5329 (
            .O(N__30082),
            .I(\uart_pc.un1_state_4_0 ));
    InMux I__5328 (
            .O(N__30077),
            .I(N__30071));
    InMux I__5327 (
            .O(N__30076),
            .I(N__30071));
    LocalMux I__5326 (
            .O(N__30071),
            .I(\uart_pc.un1_state_7_0 ));
    InMux I__5325 (
            .O(N__30068),
            .I(N__30065));
    LocalMux I__5324 (
            .O(N__30065),
            .I(N__30062));
    Span4Mux_h I__5323 (
            .O(N__30062),
            .I(N__30059));
    Odrv4 I__5322 (
            .O(N__30059),
            .I(\uart_pc.data_Auxce_0_0_0 ));
    CascadeMux I__5321 (
            .O(N__30056),
            .I(N__30053));
    InMux I__5320 (
            .O(N__30053),
            .I(N__30047));
    InMux I__5319 (
            .O(N__30052),
            .I(N__30047));
    LocalMux I__5318 (
            .O(N__30047),
            .I(N__30042));
    CascadeMux I__5317 (
            .O(N__30046),
            .I(N__30039));
    CascadeMux I__5316 (
            .O(N__30045),
            .I(N__30033));
    Span4Mux_h I__5315 (
            .O(N__30042),
            .I(N__30027));
    InMux I__5314 (
            .O(N__30039),
            .I(N__30020));
    InMux I__5313 (
            .O(N__30038),
            .I(N__30020));
    InMux I__5312 (
            .O(N__30037),
            .I(N__30020));
    InMux I__5311 (
            .O(N__30036),
            .I(N__30011));
    InMux I__5310 (
            .O(N__30033),
            .I(N__30011));
    InMux I__5309 (
            .O(N__30032),
            .I(N__30011));
    InMux I__5308 (
            .O(N__30031),
            .I(N__30011));
    InMux I__5307 (
            .O(N__30030),
            .I(N__30008));
    Odrv4 I__5306 (
            .O(N__30027),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5305 (
            .O(N__30020),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5304 (
            .O(N__30011),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    LocalMux I__5303 (
            .O(N__30008),
            .I(\uart_pc.bit_CountZ0Z_1 ));
    InMux I__5302 (
            .O(N__29999),
            .I(N__29992));
    InMux I__5301 (
            .O(N__29998),
            .I(N__29992));
    CascadeMux I__5300 (
            .O(N__29997),
            .I(N__29985));
    LocalMux I__5299 (
            .O(N__29992),
            .I(N__29980));
    InMux I__5298 (
            .O(N__29991),
            .I(N__29973));
    InMux I__5297 (
            .O(N__29990),
            .I(N__29973));
    InMux I__5296 (
            .O(N__29989),
            .I(N__29973));
    InMux I__5295 (
            .O(N__29988),
            .I(N__29966));
    InMux I__5294 (
            .O(N__29985),
            .I(N__29966));
    InMux I__5293 (
            .O(N__29984),
            .I(N__29966));
    InMux I__5292 (
            .O(N__29983),
            .I(N__29963));
    Odrv4 I__5291 (
            .O(N__29980),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5290 (
            .O(N__29973),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5289 (
            .O(N__29966),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    LocalMux I__5288 (
            .O(N__29963),
            .I(\uart_pc.bit_CountZ0Z_2 ));
    InMux I__5287 (
            .O(N__29954),
            .I(N__29948));
    InMux I__5286 (
            .O(N__29953),
            .I(N__29943));
    InMux I__5285 (
            .O(N__29952),
            .I(N__29943));
    CascadeMux I__5284 (
            .O(N__29951),
            .I(N__29937));
    LocalMux I__5283 (
            .O(N__29948),
            .I(N__29928));
    LocalMux I__5282 (
            .O(N__29943),
            .I(N__29928));
    InMux I__5281 (
            .O(N__29942),
            .I(N__29921));
    InMux I__5280 (
            .O(N__29941),
            .I(N__29921));
    InMux I__5279 (
            .O(N__29940),
            .I(N__29921));
    InMux I__5278 (
            .O(N__29937),
            .I(N__29912));
    InMux I__5277 (
            .O(N__29936),
            .I(N__29912));
    InMux I__5276 (
            .O(N__29935),
            .I(N__29912));
    InMux I__5275 (
            .O(N__29934),
            .I(N__29912));
    InMux I__5274 (
            .O(N__29933),
            .I(N__29909));
    Odrv4 I__5273 (
            .O(N__29928),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5272 (
            .O(N__29921),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5271 (
            .O(N__29912),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    LocalMux I__5270 (
            .O(N__29909),
            .I(\uart_pc.bit_CountZ0Z_0 ));
    InMux I__5269 (
            .O(N__29900),
            .I(N__29897));
    LocalMux I__5268 (
            .O(N__29897),
            .I(\uart_pc.data_Auxce_0_1 ));
    CascadeMux I__5267 (
            .O(N__29894),
            .I(N__29890));
    InMux I__5266 (
            .O(N__29893),
            .I(N__29887));
    InMux I__5265 (
            .O(N__29890),
            .I(N__29884));
    LocalMux I__5264 (
            .O(N__29887),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    LocalMux I__5263 (
            .O(N__29884),
            .I(\uart_drone.data_AuxZ0Z_0 ));
    InMux I__5262 (
            .O(N__29879),
            .I(N__29876));
    LocalMux I__5261 (
            .O(N__29876),
            .I(N__29871));
    InMux I__5260 (
            .O(N__29875),
            .I(N__29866));
    InMux I__5259 (
            .O(N__29874),
            .I(N__29866));
    Span4Mux_v I__5258 (
            .O(N__29871),
            .I(N__29863));
    LocalMux I__5257 (
            .O(N__29866),
            .I(N__29860));
    Span4Mux_h I__5256 (
            .O(N__29863),
            .I(N__29857));
    Span4Mux_v I__5255 (
            .O(N__29860),
            .I(N__29854));
    Odrv4 I__5254 (
            .O(N__29857),
            .I(\uart_drone.data_rdyc_1 ));
    Odrv4 I__5253 (
            .O(N__29854),
            .I(\uart_drone.data_rdyc_1 ));
    InMux I__5252 (
            .O(N__29849),
            .I(N__29846));
    LocalMux I__5251 (
            .O(N__29846),
            .I(N__29843));
    Odrv12 I__5250 (
            .O(N__29843),
            .I(\uart_drone_sync.aux_3__0__0_0 ));
    CascadeMux I__5249 (
            .O(N__29840),
            .I(\uart_drone.timer_Count_0_sqmuxa_cascade_ ));
    CascadeMux I__5248 (
            .O(N__29837),
            .I(\uart_pc.N_145_cascade_ ));
    InMux I__5247 (
            .O(N__29834),
            .I(N__29831));
    LocalMux I__5246 (
            .O(N__29831),
            .I(\uart_pc.N_144_1 ));
    CascadeMux I__5245 (
            .O(N__29828),
            .I(\uart_pc.N_144_1_cascade_ ));
    InMux I__5244 (
            .O(N__29825),
            .I(N__29822));
    LocalMux I__5243 (
            .O(N__29822),
            .I(N__29815));
    InMux I__5242 (
            .O(N__29821),
            .I(N__29812));
    InMux I__5241 (
            .O(N__29820),
            .I(N__29807));
    InMux I__5240 (
            .O(N__29819),
            .I(N__29807));
    InMux I__5239 (
            .O(N__29818),
            .I(N__29804));
    Odrv4 I__5238 (
            .O(N__29815),
            .I(\uart_pc.N_143 ));
    LocalMux I__5237 (
            .O(N__29812),
            .I(\uart_pc.N_143 ));
    LocalMux I__5236 (
            .O(N__29807),
            .I(\uart_pc.N_143 ));
    LocalMux I__5235 (
            .O(N__29804),
            .I(\uart_pc.N_143 ));
    InMux I__5234 (
            .O(N__29795),
            .I(N__29792));
    LocalMux I__5233 (
            .O(N__29792),
            .I(N__29784));
    InMux I__5232 (
            .O(N__29791),
            .I(N__29781));
    InMux I__5231 (
            .O(N__29790),
            .I(N__29778));
    InMux I__5230 (
            .O(N__29789),
            .I(N__29773));
    InMux I__5229 (
            .O(N__29788),
            .I(N__29773));
    InMux I__5228 (
            .O(N__29787),
            .I(N__29770));
    Odrv4 I__5227 (
            .O(N__29784),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5226 (
            .O(N__29781),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5225 (
            .O(N__29778),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5224 (
            .O(N__29773),
            .I(\uart_pc.stateZ0Z_4 ));
    LocalMux I__5223 (
            .O(N__29770),
            .I(\uart_pc.stateZ0Z_4 ));
    InMux I__5222 (
            .O(N__29759),
            .I(N__29756));
    LocalMux I__5221 (
            .O(N__29756),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_2 ));
    InMux I__5220 (
            .O(N__29753),
            .I(\uart_pc.un4_timer_Count_1_cry_1 ));
    InMux I__5219 (
            .O(N__29750),
            .I(N__29747));
    LocalMux I__5218 (
            .O(N__29747),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_3 ));
    InMux I__5217 (
            .O(N__29744),
            .I(\uart_pc.un4_timer_Count_1_cry_2 ));
    InMux I__5216 (
            .O(N__29741),
            .I(\uart_pc.un4_timer_Count_1_cry_3 ));
    InMux I__5215 (
            .O(N__29738),
            .I(N__29735));
    LocalMux I__5214 (
            .O(N__29735),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_4 ));
    CascadeMux I__5213 (
            .O(N__29732),
            .I(N__29729));
    InMux I__5212 (
            .O(N__29729),
            .I(N__29726));
    LocalMux I__5211 (
            .O(N__29726),
            .I(\uart_pc.un1_state_2_0_a3_0 ));
    InMux I__5210 (
            .O(N__29723),
            .I(N__29718));
    CascadeMux I__5209 (
            .O(N__29722),
            .I(N__29714));
    InMux I__5208 (
            .O(N__29721),
            .I(N__29711));
    LocalMux I__5207 (
            .O(N__29718),
            .I(N__29708));
    InMux I__5206 (
            .O(N__29717),
            .I(N__29703));
    InMux I__5205 (
            .O(N__29714),
            .I(N__29703));
    LocalMux I__5204 (
            .O(N__29711),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    Odrv4 I__5203 (
            .O(N__29708),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    LocalMux I__5202 (
            .O(N__29703),
            .I(\uart_pc.timer_CountZ0Z_0 ));
    InMux I__5201 (
            .O(N__29696),
            .I(N__29693));
    LocalMux I__5200 (
            .O(N__29693),
            .I(N__29686));
    CascadeMux I__5199 (
            .O(N__29692),
            .I(N__29683));
    InMux I__5198 (
            .O(N__29691),
            .I(N__29680));
    CascadeMux I__5197 (
            .O(N__29690),
            .I(N__29677));
    CascadeMux I__5196 (
            .O(N__29689),
            .I(N__29674));
    Span4Mux_v I__5195 (
            .O(N__29686),
            .I(N__29671));
    InMux I__5194 (
            .O(N__29683),
            .I(N__29668));
    LocalMux I__5193 (
            .O(N__29680),
            .I(N__29665));
    InMux I__5192 (
            .O(N__29677),
            .I(N__29660));
    InMux I__5191 (
            .O(N__29674),
            .I(N__29660));
    Odrv4 I__5190 (
            .O(N__29671),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__5189 (
            .O(N__29668),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    Odrv4 I__5188 (
            .O(N__29665),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    LocalMux I__5187 (
            .O(N__29660),
            .I(\uart_pc.timer_Count_0_sqmuxa ));
    CascadeMux I__5186 (
            .O(N__29651),
            .I(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ));
    InMux I__5185 (
            .O(N__29648),
            .I(N__29644));
    InMux I__5184 (
            .O(N__29647),
            .I(N__29641));
    LocalMux I__5183 (
            .O(N__29644),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    LocalMux I__5182 (
            .O(N__29641),
            .I(\uart_pc.timer_CountZ1Z_1 ));
    InMux I__5181 (
            .O(N__29636),
            .I(N__29633));
    LocalMux I__5180 (
            .O(N__29633),
            .I(N__29629));
    InMux I__5179 (
            .O(N__29632),
            .I(N__29626));
    Span4Mux_v I__5178 (
            .O(N__29629),
            .I(N__29623));
    LocalMux I__5177 (
            .O(N__29626),
            .I(N__29620));
    Span4Mux_h I__5176 (
            .O(N__29623),
            .I(N__29615));
    Span4Mux_h I__5175 (
            .O(N__29620),
            .I(N__29615));
    Odrv4 I__5174 (
            .O(N__29615),
            .I(drone_H_disp_side_13));
    CascadeMux I__5173 (
            .O(N__29612),
            .I(N__29608));
    InMux I__5172 (
            .O(N__29611),
            .I(N__29603));
    InMux I__5171 (
            .O(N__29608),
            .I(N__29603));
    LocalMux I__5170 (
            .O(N__29603),
            .I(N__29600));
    Span4Mux_h I__5169 (
            .O(N__29600),
            .I(N__29597));
    Span4Mux_h I__5168 (
            .O(N__29597),
            .I(N__29594));
    Odrv4 I__5167 (
            .O(N__29594),
            .I(drone_H_disp_side_14));
    CEMux I__5166 (
            .O(N__29591),
            .I(N__29588));
    LocalMux I__5165 (
            .O(N__29588),
            .I(N__29584));
    CEMux I__5164 (
            .O(N__29587),
            .I(N__29581));
    Span4Mux_v I__5163 (
            .O(N__29584),
            .I(N__29575));
    LocalMux I__5162 (
            .O(N__29581),
            .I(N__29575));
    CEMux I__5161 (
            .O(N__29580),
            .I(N__29572));
    Span4Mux_h I__5160 (
            .O(N__29575),
            .I(N__29569));
    LocalMux I__5159 (
            .O(N__29572),
            .I(N__29566));
    Span4Mux_h I__5158 (
            .O(N__29569),
            .I(N__29563));
    Span4Mux_v I__5157 (
            .O(N__29566),
            .I(N__29560));
    Span4Mux_v I__5156 (
            .O(N__29563),
            .I(N__29557));
    Span4Mux_v I__5155 (
            .O(N__29560),
            .I(N__29554));
    Odrv4 I__5154 (
            .O(N__29557),
            .I(\dron_frame_decoder_1.N_739_0 ));
    Odrv4 I__5153 (
            .O(N__29554),
            .I(\dron_frame_decoder_1.N_739_0 ));
    CascadeMux I__5152 (
            .O(N__29549),
            .I(N__29546));
    InMux I__5151 (
            .O(N__29546),
            .I(N__29543));
    LocalMux I__5150 (
            .O(N__29543),
            .I(N__29539));
    InMux I__5149 (
            .O(N__29542),
            .I(N__29535));
    Span12Mux_s10_h I__5148 (
            .O(N__29539),
            .I(N__29532));
    InMux I__5147 (
            .O(N__29538),
            .I(N__29529));
    LocalMux I__5146 (
            .O(N__29535),
            .I(drone_H_disp_side_12));
    Odrv12 I__5145 (
            .O(N__29532),
            .I(drone_H_disp_side_12));
    LocalMux I__5144 (
            .O(N__29529),
            .I(drone_H_disp_side_12));
    CascadeMux I__5143 (
            .O(N__29522),
            .I(N__29519));
    InMux I__5142 (
            .O(N__29519),
            .I(N__29516));
    LocalMux I__5141 (
            .O(N__29516),
            .I(N__29513));
    Odrv12 I__5140 (
            .O(N__29513),
            .I(drone_H_disp_side_i_12));
    InMux I__5139 (
            .O(N__29510),
            .I(N__29507));
    LocalMux I__5138 (
            .O(N__29507),
            .I(drone_H_disp_front_3));
    InMux I__5137 (
            .O(N__29504),
            .I(N__29500));
    InMux I__5136 (
            .O(N__29503),
            .I(N__29497));
    LocalMux I__5135 (
            .O(N__29500),
            .I(N__29494));
    LocalMux I__5134 (
            .O(N__29497),
            .I(N__29491));
    Span4Mux_v I__5133 (
            .O(N__29494),
            .I(N__29488));
    Span4Mux_v I__5132 (
            .O(N__29491),
            .I(N__29485));
    Sp12to4 I__5131 (
            .O(N__29488),
            .I(N__29482));
    Span4Mux_v I__5130 (
            .O(N__29485),
            .I(N__29479));
    Span12Mux_s3_h I__5129 (
            .O(N__29482),
            .I(N__29476));
    Sp12to4 I__5128 (
            .O(N__29479),
            .I(N__29473));
    Span12Mux_h I__5127 (
            .O(N__29476),
            .I(N__29470));
    Odrv12 I__5126 (
            .O(N__29473),
            .I(xy_kp_3));
    Odrv12 I__5125 (
            .O(N__29470),
            .I(xy_kp_3));
    InMux I__5124 (
            .O(N__29465),
            .I(N__29462));
    LocalMux I__5123 (
            .O(N__29462),
            .I(N__29459));
    Span4Mux_h I__5122 (
            .O(N__29459),
            .I(N__29456));
    Odrv4 I__5121 (
            .O(N__29456),
            .I(\uart_drone_sync.aux_2__0__0_0 ));
    CascadeMux I__5120 (
            .O(N__29453),
            .I(\pid_alt.un1_reset_i_a5_1_10_5_cascade_ ));
    InMux I__5119 (
            .O(N__29450),
            .I(N__29445));
    InMux I__5118 (
            .O(N__29449),
            .I(N__29440));
    InMux I__5117 (
            .O(N__29448),
            .I(N__29440));
    LocalMux I__5116 (
            .O(N__29445),
            .I(N__29437));
    LocalMux I__5115 (
            .O(N__29440),
            .I(N__29434));
    Span4Mux_h I__5114 (
            .O(N__29437),
            .I(N__29431));
    Span4Mux_h I__5113 (
            .O(N__29434),
            .I(N__29428));
    Span4Mux_h I__5112 (
            .O(N__29431),
            .I(N__29425));
    Span4Mux_h I__5111 (
            .O(N__29428),
            .I(N__29422));
    Odrv4 I__5110 (
            .O(N__29425),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    Odrv4 I__5109 (
            .O(N__29422),
            .I(\pid_alt.pid_preregZ0Z_6 ));
    InMux I__5108 (
            .O(N__29417),
            .I(N__29414));
    LocalMux I__5107 (
            .O(N__29414),
            .I(N__29411));
    Span4Mux_v I__5106 (
            .O(N__29411),
            .I(N__29408));
    Odrv4 I__5105 (
            .O(N__29408),
            .I(\pid_side.un1_pid_prereg_cry_9_THRU_CO ));
    InMux I__5104 (
            .O(N__29405),
            .I(N__29401));
    InMux I__5103 (
            .O(N__29404),
            .I(N__29398));
    LocalMux I__5102 (
            .O(N__29401),
            .I(N__29395));
    LocalMux I__5101 (
            .O(N__29398),
            .I(N__29392));
    Span4Mux_h I__5100 (
            .O(N__29395),
            .I(N__29388));
    Span12Mux_h I__5099 (
            .O(N__29392),
            .I(N__29385));
    InMux I__5098 (
            .O(N__29391),
            .I(N__29382));
    Span4Mux_h I__5097 (
            .O(N__29388),
            .I(N__29379));
    Odrv12 I__5096 (
            .O(N__29385),
            .I(\pid_side.error_p_regZ0Z_10 ));
    LocalMux I__5095 (
            .O(N__29382),
            .I(\pid_side.error_p_regZ0Z_10 ));
    Odrv4 I__5094 (
            .O(N__29379),
            .I(\pid_side.error_p_regZ0Z_10 ));
    CascadeMux I__5093 (
            .O(N__29372),
            .I(\pid_side.un1_reset_i_a2_3_cascade_ ));
    InMux I__5092 (
            .O(N__29369),
            .I(N__29365));
    InMux I__5091 (
            .O(N__29368),
            .I(N__29362));
    LocalMux I__5090 (
            .O(N__29365),
            .I(\pid_side.pid_preregZ0Z_18 ));
    LocalMux I__5089 (
            .O(N__29362),
            .I(\pid_side.pid_preregZ0Z_18 ));
    InMux I__5088 (
            .O(N__29357),
            .I(N__29353));
    InMux I__5087 (
            .O(N__29356),
            .I(N__29350));
    LocalMux I__5086 (
            .O(N__29353),
            .I(\pid_side.pid_preregZ0Z_17 ));
    LocalMux I__5085 (
            .O(N__29350),
            .I(\pid_side.pid_preregZ0Z_17 ));
    CascadeMux I__5084 (
            .O(N__29345),
            .I(N__29341));
    InMux I__5083 (
            .O(N__29344),
            .I(N__29338));
    InMux I__5082 (
            .O(N__29341),
            .I(N__29335));
    LocalMux I__5081 (
            .O(N__29338),
            .I(\pid_side.pid_preregZ0Z_19 ));
    LocalMux I__5080 (
            .O(N__29335),
            .I(\pid_side.pid_preregZ0Z_19 ));
    CascadeMux I__5079 (
            .O(N__29330),
            .I(N__29327));
    InMux I__5078 (
            .O(N__29327),
            .I(N__29323));
    InMux I__5077 (
            .O(N__29326),
            .I(N__29320));
    LocalMux I__5076 (
            .O(N__29323),
            .I(\pid_side.pid_preregZ0Z_20 ));
    LocalMux I__5075 (
            .O(N__29320),
            .I(\pid_side.pid_preregZ0Z_20 ));
    InMux I__5074 (
            .O(N__29315),
            .I(N__29311));
    InMux I__5073 (
            .O(N__29314),
            .I(N__29308));
    LocalMux I__5072 (
            .O(N__29311),
            .I(N__29305));
    LocalMux I__5071 (
            .O(N__29308),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    Odrv12 I__5070 (
            .O(N__29305),
            .I(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ));
    InMux I__5069 (
            .O(N__29300),
            .I(N__29294));
    InMux I__5068 (
            .O(N__29299),
            .I(N__29294));
    LocalMux I__5067 (
            .O(N__29294),
            .I(drone_H_disp_side_11));
    CEMux I__5066 (
            .O(N__29291),
            .I(N__29288));
    LocalMux I__5065 (
            .O(N__29288),
            .I(N__29285));
    Span4Mux_v I__5064 (
            .O(N__29285),
            .I(N__29281));
    CEMux I__5063 (
            .O(N__29284),
            .I(N__29278));
    Span4Mux_h I__5062 (
            .O(N__29281),
            .I(N__29275));
    LocalMux I__5061 (
            .O(N__29278),
            .I(N__29272));
    Odrv4 I__5060 (
            .O(N__29275),
            .I(\uart_drone.data_rdyc_1_0 ));
    Odrv12 I__5059 (
            .O(N__29272),
            .I(\uart_drone.data_rdyc_1_0 ));
    SRMux I__5058 (
            .O(N__29267),
            .I(N__29263));
    SRMux I__5057 (
            .O(N__29266),
            .I(N__29260));
    LocalMux I__5056 (
            .O(N__29263),
            .I(N__29257));
    LocalMux I__5055 (
            .O(N__29260),
            .I(N__29254));
    Span4Mux_h I__5054 (
            .O(N__29257),
            .I(N__29251));
    Span4Mux_h I__5053 (
            .O(N__29254),
            .I(N__29248));
    Odrv4 I__5052 (
            .O(N__29251),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    Odrv4 I__5051 (
            .O(N__29248),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ));
    CascadeMux I__5050 (
            .O(N__29243),
            .I(N__29240));
    InMux I__5049 (
            .O(N__29240),
            .I(N__29235));
    InMux I__5048 (
            .O(N__29239),
            .I(N__29232));
    InMux I__5047 (
            .O(N__29238),
            .I(N__29229));
    LocalMux I__5046 (
            .O(N__29235),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__5045 (
            .O(N__29232),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    LocalMux I__5044 (
            .O(N__29229),
            .I(\dron_frame_decoder_1.stateZ0Z_2 ));
    CascadeMux I__5043 (
            .O(N__29222),
            .I(N__29217));
    InMux I__5042 (
            .O(N__29221),
            .I(N__29214));
    InMux I__5041 (
            .O(N__29220),
            .I(N__29207));
    InMux I__5040 (
            .O(N__29217),
            .I(N__29200));
    LocalMux I__5039 (
            .O(N__29214),
            .I(N__29197));
    InMux I__5038 (
            .O(N__29213),
            .I(N__29192));
    InMux I__5037 (
            .O(N__29212),
            .I(N__29187));
    InMux I__5036 (
            .O(N__29211),
            .I(N__29187));
    InMux I__5035 (
            .O(N__29210),
            .I(N__29184));
    LocalMux I__5034 (
            .O(N__29207),
            .I(N__29181));
    InMux I__5033 (
            .O(N__29206),
            .I(N__29178));
    InMux I__5032 (
            .O(N__29205),
            .I(N__29171));
    InMux I__5031 (
            .O(N__29204),
            .I(N__29171));
    InMux I__5030 (
            .O(N__29203),
            .I(N__29171));
    LocalMux I__5029 (
            .O(N__29200),
            .I(N__29166));
    Span4Mux_v I__5028 (
            .O(N__29197),
            .I(N__29166));
    InMux I__5027 (
            .O(N__29196),
            .I(N__29161));
    InMux I__5026 (
            .O(N__29195),
            .I(N__29161));
    LocalMux I__5025 (
            .O(N__29192),
            .I(uart_drone_data_rdy));
    LocalMux I__5024 (
            .O(N__29187),
            .I(uart_drone_data_rdy));
    LocalMux I__5023 (
            .O(N__29184),
            .I(uart_drone_data_rdy));
    Odrv4 I__5022 (
            .O(N__29181),
            .I(uart_drone_data_rdy));
    LocalMux I__5021 (
            .O(N__29178),
            .I(uart_drone_data_rdy));
    LocalMux I__5020 (
            .O(N__29171),
            .I(uart_drone_data_rdy));
    Odrv4 I__5019 (
            .O(N__29166),
            .I(uart_drone_data_rdy));
    LocalMux I__5018 (
            .O(N__29161),
            .I(uart_drone_data_rdy));
    InMux I__5017 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__5016 (
            .O(N__29141),
            .I(N__29136));
    InMux I__5015 (
            .O(N__29140),
            .I(N__29133));
    InMux I__5014 (
            .O(N__29139),
            .I(N__29130));
    Span4Mux_v I__5013 (
            .O(N__29136),
            .I(N__29127));
    LocalMux I__5012 (
            .O(N__29133),
            .I(N__29124));
    LocalMux I__5011 (
            .O(N__29130),
            .I(N__29121));
    Span4Mux_h I__5010 (
            .O(N__29127),
            .I(N__29116));
    Span4Mux_v I__5009 (
            .O(N__29124),
            .I(N__29116));
    Span12Mux_h I__5008 (
            .O(N__29121),
            .I(N__29113));
    Odrv4 I__5007 (
            .O(N__29116),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    Odrv12 I__5006 (
            .O(N__29113),
            .I(\pid_alt.pid_preregZ0Z_10 ));
    CascadeMux I__5005 (
            .O(N__29108),
            .I(\pid_alt.un1_reset_i_a2_3_cascade_ ));
    InMux I__5004 (
            .O(N__29105),
            .I(N__29102));
    LocalMux I__5003 (
            .O(N__29102),
            .I(N__29099));
    Span4Mux_v I__5002 (
            .O(N__29099),
            .I(N__29094));
    InMux I__5001 (
            .O(N__29098),
            .I(N__29089));
    InMux I__5000 (
            .O(N__29097),
            .I(N__29089));
    Sp12to4 I__4999 (
            .O(N__29094),
            .I(N__29084));
    LocalMux I__4998 (
            .O(N__29089),
            .I(N__29084));
    Odrv12 I__4997 (
            .O(N__29084),
            .I(\pid_alt.pid_preregZ0Z_8 ));
    CascadeMux I__4996 (
            .O(N__29081),
            .I(N__29078));
    InMux I__4995 (
            .O(N__29078),
            .I(N__29075));
    LocalMux I__4994 (
            .O(N__29075),
            .I(N__29071));
    CascadeMux I__4993 (
            .O(N__29074),
            .I(N__29068));
    Span4Mux_h I__4992 (
            .O(N__29071),
            .I(N__29065));
    InMux I__4991 (
            .O(N__29068),
            .I(N__29062));
    Odrv4 I__4990 (
            .O(N__29065),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    LocalMux I__4989 (
            .O(N__29062),
            .I(\uart_pc.data_AuxZ0Z_5 ));
    InMux I__4988 (
            .O(N__29057),
            .I(N__29054));
    LocalMux I__4987 (
            .O(N__29054),
            .I(N__29051));
    Span4Mux_v I__4986 (
            .O(N__29051),
            .I(N__29048));
    Odrv4 I__4985 (
            .O(N__29048),
            .I(\uart_pc.data_Auxce_0_0_4 ));
    InMux I__4984 (
            .O(N__29045),
            .I(N__29042));
    LocalMux I__4983 (
            .O(N__29042),
            .I(\uart_pc.data_Auxce_0_5 ));
    InMux I__4982 (
            .O(N__29039),
            .I(N__29036));
    LocalMux I__4981 (
            .O(N__29036),
            .I(N__29033));
    Odrv4 I__4980 (
            .O(N__29033),
            .I(\uart_pc.data_Auxce_0_0_2 ));
    CascadeMux I__4979 (
            .O(N__29030),
            .I(N__29025));
    InMux I__4978 (
            .O(N__29029),
            .I(N__29022));
    InMux I__4977 (
            .O(N__29028),
            .I(N__29017));
    InMux I__4976 (
            .O(N__29025),
            .I(N__29017));
    LocalMux I__4975 (
            .O(N__29022),
            .I(\uart_drone.stateZ0Z_1 ));
    LocalMux I__4974 (
            .O(N__29017),
            .I(\uart_drone.stateZ0Z_1 ));
    CascadeMux I__4973 (
            .O(N__29012),
            .I(\uart_drone.state_srsts_i_0_2_cascade_ ));
    InMux I__4972 (
            .O(N__29009),
            .I(N__29004));
    CascadeMux I__4971 (
            .O(N__29008),
            .I(N__29001));
    InMux I__4970 (
            .O(N__29007),
            .I(N__28997));
    LocalMux I__4969 (
            .O(N__29004),
            .I(N__28994));
    InMux I__4968 (
            .O(N__29001),
            .I(N__28989));
    InMux I__4967 (
            .O(N__29000),
            .I(N__28989));
    LocalMux I__4966 (
            .O(N__28997),
            .I(\scaler_4.un2_source_data_0 ));
    Odrv4 I__4965 (
            .O(N__28994),
            .I(\scaler_4.un2_source_data_0 ));
    LocalMux I__4964 (
            .O(N__28989),
            .I(\scaler_4.un2_source_data_0 ));
    InMux I__4963 (
            .O(N__28982),
            .I(N__28978));
    InMux I__4962 (
            .O(N__28981),
            .I(N__28975));
    LocalMux I__4961 (
            .O(N__28978),
            .I(N__28969));
    LocalMux I__4960 (
            .O(N__28975),
            .I(N__28969));
    CascadeMux I__4959 (
            .O(N__28974),
            .I(N__28965));
    Span4Mux_v I__4958 (
            .O(N__28969),
            .I(N__28962));
    InMux I__4957 (
            .O(N__28968),
            .I(N__28959));
    InMux I__4956 (
            .O(N__28965),
            .I(N__28956));
    Odrv4 I__4955 (
            .O(N__28962),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__4954 (
            .O(N__28959),
            .I(frame_decoder_OFF4data_0));
    LocalMux I__4953 (
            .O(N__28956),
            .I(frame_decoder_OFF4data_0));
    InMux I__4952 (
            .O(N__28949),
            .I(N__28945));
    InMux I__4951 (
            .O(N__28948),
            .I(N__28942));
    LocalMux I__4950 (
            .O(N__28945),
            .I(N__28939));
    LocalMux I__4949 (
            .O(N__28942),
            .I(N__28934));
    Span4Mux_h I__4948 (
            .O(N__28939),
            .I(N__28931));
    InMux I__4947 (
            .O(N__28938),
            .I(N__28928));
    InMux I__4946 (
            .O(N__28937),
            .I(N__28925));
    Odrv4 I__4945 (
            .O(N__28934),
            .I(frame_decoder_CH4data_0));
    Odrv4 I__4944 (
            .O(N__28931),
            .I(frame_decoder_CH4data_0));
    LocalMux I__4943 (
            .O(N__28928),
            .I(frame_decoder_CH4data_0));
    LocalMux I__4942 (
            .O(N__28925),
            .I(frame_decoder_CH4data_0));
    CEMux I__4941 (
            .O(N__28916),
            .I(N__28913));
    LocalMux I__4940 (
            .O(N__28913),
            .I(N__28908));
    CEMux I__4939 (
            .O(N__28912),
            .I(N__28905));
    CEMux I__4938 (
            .O(N__28911),
            .I(N__28902));
    Span4Mux_h I__4937 (
            .O(N__28908),
            .I(N__28897));
    LocalMux I__4936 (
            .O(N__28905),
            .I(N__28897));
    LocalMux I__4935 (
            .O(N__28902),
            .I(N__28894));
    Span4Mux_v I__4934 (
            .O(N__28897),
            .I(N__28891));
    Span4Mux_h I__4933 (
            .O(N__28894),
            .I(N__28888));
    Span4Mux_h I__4932 (
            .O(N__28891),
            .I(N__28885));
    Span4Mux_v I__4931 (
            .O(N__28888),
            .I(N__28882));
    Span4Mux_h I__4930 (
            .O(N__28885),
            .I(N__28879));
    Odrv4 I__4929 (
            .O(N__28882),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    Odrv4 I__4928 (
            .O(N__28879),
            .I(\scaler_4.debug_CH3_20A_c_0 ));
    InMux I__4927 (
            .O(N__28874),
            .I(N__28870));
    CascadeMux I__4926 (
            .O(N__28873),
            .I(N__28867));
    LocalMux I__4925 (
            .O(N__28870),
            .I(N__28864));
    InMux I__4924 (
            .O(N__28867),
            .I(N__28861));
    Odrv12 I__4923 (
            .O(N__28864),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    LocalMux I__4922 (
            .O(N__28861),
            .I(\uart_pc.data_AuxZ1Z_2 ));
    CascadeMux I__4921 (
            .O(N__28856),
            .I(N__28853));
    InMux I__4920 (
            .O(N__28853),
            .I(N__28849));
    CascadeMux I__4919 (
            .O(N__28852),
            .I(N__28846));
    LocalMux I__4918 (
            .O(N__28849),
            .I(N__28843));
    InMux I__4917 (
            .O(N__28846),
            .I(N__28840));
    Odrv4 I__4916 (
            .O(N__28843),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    LocalMux I__4915 (
            .O(N__28840),
            .I(\uart_pc.data_AuxZ1Z_1 ));
    InMux I__4914 (
            .O(N__28835),
            .I(N__28832));
    LocalMux I__4913 (
            .O(N__28832),
            .I(\uart_pc.data_Auxce_0_3 ));
    InMux I__4912 (
            .O(N__28829),
            .I(N__28825));
    CascadeMux I__4911 (
            .O(N__28828),
            .I(N__28822));
    LocalMux I__4910 (
            .O(N__28825),
            .I(N__28819));
    InMux I__4909 (
            .O(N__28822),
            .I(N__28816));
    Odrv4 I__4908 (
            .O(N__28819),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    LocalMux I__4907 (
            .O(N__28816),
            .I(\uart_pc.data_AuxZ0Z_3 ));
    CEMux I__4906 (
            .O(N__28811),
            .I(N__28808));
    LocalMux I__4905 (
            .O(N__28808),
            .I(\pid_alt.state_1_0_0 ));
    CascadeMux I__4904 (
            .O(N__28805),
            .I(\uart_pc.state_srsts_0_0_0_cascade_ ));
    CascadeMux I__4903 (
            .O(N__28802),
            .I(\uart_pc.N_143_cascade_ ));
    InMux I__4902 (
            .O(N__28799),
            .I(N__28796));
    LocalMux I__4901 (
            .O(N__28796),
            .I(N__28793));
    Span4Mux_h I__4900 (
            .O(N__28793),
            .I(N__28788));
    InMux I__4899 (
            .O(N__28792),
            .I(N__28783));
    InMux I__4898 (
            .O(N__28791),
            .I(N__28783));
    Odrv4 I__4897 (
            .O(N__28788),
            .I(\uart_pc.data_rdyc_1 ));
    LocalMux I__4896 (
            .O(N__28783),
            .I(\uart_pc.data_rdyc_1 ));
    CascadeMux I__4895 (
            .O(N__28778),
            .I(\uart_pc.data_rdyc_1_cascade_ ));
    InMux I__4894 (
            .O(N__28775),
            .I(N__28770));
    InMux I__4893 (
            .O(N__28774),
            .I(N__28766));
    InMux I__4892 (
            .O(N__28773),
            .I(N__28763));
    LocalMux I__4891 (
            .O(N__28770),
            .I(N__28760));
    InMux I__4890 (
            .O(N__28769),
            .I(N__28757));
    LocalMux I__4889 (
            .O(N__28766),
            .I(N__28753));
    LocalMux I__4888 (
            .O(N__28763),
            .I(N__28750));
    Span4Mux_v I__4887 (
            .O(N__28760),
            .I(N__28745));
    LocalMux I__4886 (
            .O(N__28757),
            .I(N__28745));
    InMux I__4885 (
            .O(N__28756),
            .I(N__28742));
    Span4Mux_v I__4884 (
            .O(N__28753),
            .I(N__28736));
    Span4Mux_v I__4883 (
            .O(N__28750),
            .I(N__28736));
    Span4Mux_h I__4882 (
            .O(N__28745),
            .I(N__28731));
    LocalMux I__4881 (
            .O(N__28742),
            .I(N__28731));
    CascadeMux I__4880 (
            .O(N__28741),
            .I(N__28727));
    Span4Mux_v I__4879 (
            .O(N__28736),
            .I(N__28724));
    Span4Mux_h I__4878 (
            .O(N__28731),
            .I(N__28721));
    InMux I__4877 (
            .O(N__28730),
            .I(N__28716));
    InMux I__4876 (
            .O(N__28727),
            .I(N__28716));
    Odrv4 I__4875 (
            .O(N__28724),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    Odrv4 I__4874 (
            .O(N__28721),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    LocalMux I__4873 (
            .O(N__28716),
            .I(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ));
    InMux I__4872 (
            .O(N__28709),
            .I(N__28705));
    InMux I__4871 (
            .O(N__28708),
            .I(N__28702));
    LocalMux I__4870 (
            .O(N__28705),
            .I(N__28699));
    LocalMux I__4869 (
            .O(N__28702),
            .I(N__28696));
    Span4Mux_v I__4868 (
            .O(N__28699),
            .I(N__28692));
    Span12Mux_h I__4867 (
            .O(N__28696),
            .I(N__28689));
    InMux I__4866 (
            .O(N__28695),
            .I(N__28686));
    Span4Mux_h I__4865 (
            .O(N__28692),
            .I(N__28683));
    Odrv12 I__4864 (
            .O(N__28689),
            .I(\pid_side.error_p_regZ0Z_12 ));
    LocalMux I__4863 (
            .O(N__28686),
            .I(\pid_side.error_p_regZ0Z_12 ));
    Odrv4 I__4862 (
            .O(N__28683),
            .I(\pid_side.error_p_regZ0Z_12 ));
    InMux I__4861 (
            .O(N__28676),
            .I(N__28673));
    LocalMux I__4860 (
            .O(N__28673),
            .I(\pid_side.un1_pid_prereg_cry_11_THRU_CO ));
    InMux I__4859 (
            .O(N__28670),
            .I(N__28667));
    LocalMux I__4858 (
            .O(N__28667),
            .I(\pid_side.un1_pid_prereg_cry_17_THRU_CO ));
    CascadeMux I__4857 (
            .O(N__28664),
            .I(N__28661));
    InMux I__4856 (
            .O(N__28661),
            .I(N__28658));
    LocalMux I__4855 (
            .O(N__28658),
            .I(N__28654));
    InMux I__4854 (
            .O(N__28657),
            .I(N__28651));
    Span4Mux_h I__4853 (
            .O(N__28654),
            .I(N__28646));
    LocalMux I__4852 (
            .O(N__28651),
            .I(N__28646));
    Span4Mux_h I__4851 (
            .O(N__28646),
            .I(N__28642));
    InMux I__4850 (
            .O(N__28645),
            .I(N__28639));
    Span4Mux_h I__4849 (
            .O(N__28642),
            .I(N__28636));
    LocalMux I__4848 (
            .O(N__28639),
            .I(\pid_side.error_p_regZ0Z_18 ));
    Odrv4 I__4847 (
            .O(N__28636),
            .I(\pid_side.error_p_regZ0Z_18 ));
    InMux I__4846 (
            .O(N__28631),
            .I(N__28628));
    LocalMux I__4845 (
            .O(N__28628),
            .I(N__28625));
    Span12Mux_v I__4844 (
            .O(N__28625),
            .I(N__28621));
    InMux I__4843 (
            .O(N__28624),
            .I(N__28618));
    Odrv12 I__4842 (
            .O(N__28621),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    LocalMux I__4841 (
            .O(N__28618),
            .I(\pid_alt.error_d_reg_prevZ0Z_15 ));
    InMux I__4840 (
            .O(N__28613),
            .I(N__28609));
    CascadeMux I__4839 (
            .O(N__28612),
            .I(N__28606));
    LocalMux I__4838 (
            .O(N__28609),
            .I(N__28603));
    InMux I__4837 (
            .O(N__28606),
            .I(N__28600));
    Span4Mux_v I__4836 (
            .O(N__28603),
            .I(N__28597));
    LocalMux I__4835 (
            .O(N__28600),
            .I(N__28594));
    Span4Mux_h I__4834 (
            .O(N__28597),
            .I(N__28591));
    Span12Mux_v I__4833 (
            .O(N__28594),
            .I(N__28588));
    Odrv4 I__4832 (
            .O(N__28591),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    Odrv12 I__4831 (
            .O(N__28588),
            .I(\pid_alt.error_p_regZ0Z_15 ));
    InMux I__4830 (
            .O(N__28583),
            .I(N__28580));
    LocalMux I__4829 (
            .O(N__28580),
            .I(N__28577));
    Span4Mux_v I__4828 (
            .O(N__28577),
            .I(N__28573));
    InMux I__4827 (
            .O(N__28576),
            .I(N__28569));
    Span4Mux_h I__4826 (
            .O(N__28573),
            .I(N__28566));
    InMux I__4825 (
            .O(N__28572),
            .I(N__28563));
    LocalMux I__4824 (
            .O(N__28569),
            .I(N__28558));
    Span4Mux_v I__4823 (
            .O(N__28566),
            .I(N__28558));
    LocalMux I__4822 (
            .O(N__28563),
            .I(N__28555));
    Span4Mux_v I__4821 (
            .O(N__28558),
            .I(N__28552));
    Span4Mux_v I__4820 (
            .O(N__28555),
            .I(N__28549));
    Span4Mux_h I__4819 (
            .O(N__28552),
            .I(N__28546));
    Span4Mux_v I__4818 (
            .O(N__28549),
            .I(N__28543));
    Odrv4 I__4817 (
            .O(N__28546),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    Odrv4 I__4816 (
            .O(N__28543),
            .I(\pid_alt.error_d_regZ0Z_15 ));
    InMux I__4815 (
            .O(N__28538),
            .I(N__28532));
    InMux I__4814 (
            .O(N__28537),
            .I(N__28532));
    LocalMux I__4813 (
            .O(N__28532),
            .I(N__28529));
    Span4Mux_h I__4812 (
            .O(N__28529),
            .I(N__28526));
    Span4Mux_h I__4811 (
            .O(N__28526),
            .I(N__28523));
    Odrv4 I__4810 (
            .O(N__28523),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ));
    InMux I__4809 (
            .O(N__28520),
            .I(N__28517));
    LocalMux I__4808 (
            .O(N__28517),
            .I(N__28514));
    Span4Mux_h I__4807 (
            .O(N__28514),
            .I(N__28511));
    Span4Mux_h I__4806 (
            .O(N__28511),
            .I(N__28508));
    Odrv4 I__4805 (
            .O(N__28508),
            .I(\pid_side.error_axb_8_l_ofxZ0 ));
    CascadeMux I__4804 (
            .O(N__28505),
            .I(N__28502));
    InMux I__4803 (
            .O(N__28502),
            .I(N__28496));
    InMux I__4802 (
            .O(N__28501),
            .I(N__28496));
    LocalMux I__4801 (
            .O(N__28496),
            .I(side_command_7));
    InMux I__4800 (
            .O(N__28493),
            .I(N__28490));
    LocalMux I__4799 (
            .O(N__28490),
            .I(N__28487));
    Span4Mux_h I__4798 (
            .O(N__28487),
            .I(N__28484));
    Span4Mux_h I__4797 (
            .O(N__28484),
            .I(N__28481));
    Odrv4 I__4796 (
            .O(N__28481),
            .I(\pid_side.error_axbZ0Z_7 ));
    InMux I__4795 (
            .O(N__28478),
            .I(N__28475));
    LocalMux I__4794 (
            .O(N__28475),
            .I(drone_H_disp_front_2));
    InMux I__4793 (
            .O(N__28472),
            .I(N__28469));
    LocalMux I__4792 (
            .O(N__28469),
            .I(drone_H_disp_side_1));
    InMux I__4791 (
            .O(N__28466),
            .I(N__28463));
    LocalMux I__4790 (
            .O(N__28463),
            .I(N__28460));
    Odrv12 I__4789 (
            .O(N__28460),
            .I(\pid_side.error_axbZ0Z_1 ));
    InMux I__4788 (
            .O(N__28457),
            .I(N__28454));
    LocalMux I__4787 (
            .O(N__28454),
            .I(\pid_side.un1_pid_prereg_cry_7_THRU_CO ));
    InMux I__4786 (
            .O(N__28451),
            .I(N__28447));
    InMux I__4785 (
            .O(N__28450),
            .I(N__28444));
    LocalMux I__4784 (
            .O(N__28447),
            .I(N__28439));
    LocalMux I__4783 (
            .O(N__28444),
            .I(N__28439));
    Span4Mux_v I__4782 (
            .O(N__28439),
            .I(N__28435));
    InMux I__4781 (
            .O(N__28438),
            .I(N__28432));
    Span4Mux_h I__4780 (
            .O(N__28435),
            .I(N__28429));
    LocalMux I__4779 (
            .O(N__28432),
            .I(\pid_side.error_p_regZ0Z_8 ));
    Odrv4 I__4778 (
            .O(N__28429),
            .I(\pid_side.error_p_regZ0Z_8 ));
    InMux I__4777 (
            .O(N__28424),
            .I(N__28421));
    LocalMux I__4776 (
            .O(N__28421),
            .I(N__28417));
    InMux I__4775 (
            .O(N__28420),
            .I(N__28414));
    Span4Mux_v I__4774 (
            .O(N__28417),
            .I(N__28409));
    LocalMux I__4773 (
            .O(N__28414),
            .I(N__28409));
    Span4Mux_h I__4772 (
            .O(N__28409),
            .I(N__28405));
    InMux I__4771 (
            .O(N__28408),
            .I(N__28402));
    Span4Mux_h I__4770 (
            .O(N__28405),
            .I(N__28399));
    LocalMux I__4769 (
            .O(N__28402),
            .I(\pid_side.error_p_regZ0Z_11 ));
    Odrv4 I__4768 (
            .O(N__28399),
            .I(\pid_side.error_p_regZ0Z_11 ));
    InMux I__4767 (
            .O(N__28394),
            .I(N__28391));
    LocalMux I__4766 (
            .O(N__28391),
            .I(\pid_side.un1_pid_prereg_cry_10_THRU_CO ));
    InMux I__4765 (
            .O(N__28388),
            .I(N__28385));
    LocalMux I__4764 (
            .O(N__28385),
            .I(\pid_side.un1_pid_prereg_cry_3_THRU_CO ));
    InMux I__4763 (
            .O(N__28382),
            .I(N__28378));
    InMux I__4762 (
            .O(N__28381),
            .I(N__28375));
    LocalMux I__4761 (
            .O(N__28378),
            .I(N__28372));
    LocalMux I__4760 (
            .O(N__28375),
            .I(N__28369));
    Span4Mux_v I__4759 (
            .O(N__28372),
            .I(N__28363));
    Span4Mux_v I__4758 (
            .O(N__28369),
            .I(N__28363));
    InMux I__4757 (
            .O(N__28368),
            .I(N__28360));
    Span4Mux_h I__4756 (
            .O(N__28363),
            .I(N__28357));
    LocalMux I__4755 (
            .O(N__28360),
            .I(\pid_side.error_p_regZ0Z_4 ));
    Odrv4 I__4754 (
            .O(N__28357),
            .I(\pid_side.error_p_regZ0Z_4 ));
    InMux I__4753 (
            .O(N__28352),
            .I(N__28349));
    LocalMux I__4752 (
            .O(N__28349),
            .I(N__28345));
    InMux I__4751 (
            .O(N__28348),
            .I(N__28342));
    Span4Mux_h I__4750 (
            .O(N__28345),
            .I(N__28337));
    LocalMux I__4749 (
            .O(N__28342),
            .I(N__28337));
    Span4Mux_h I__4748 (
            .O(N__28337),
            .I(N__28333));
    InMux I__4747 (
            .O(N__28336),
            .I(N__28330));
    Span4Mux_h I__4746 (
            .O(N__28333),
            .I(N__28327));
    LocalMux I__4745 (
            .O(N__28330),
            .I(\pid_side.error_p_regZ0Z_6 ));
    Odrv4 I__4744 (
            .O(N__28327),
            .I(\pid_side.error_p_regZ0Z_6 ));
    InMux I__4743 (
            .O(N__28322),
            .I(N__28319));
    LocalMux I__4742 (
            .O(N__28319),
            .I(\pid_side.un1_pid_prereg_cry_5_THRU_CO ));
    InMux I__4741 (
            .O(N__28316),
            .I(N__28313));
    LocalMux I__4740 (
            .O(N__28313),
            .I(\pid_side.un1_pid_prereg_cry_18_THRU_CO ));
    CascadeMux I__4739 (
            .O(N__28310),
            .I(N__28307));
    InMux I__4738 (
            .O(N__28307),
            .I(N__28303));
    InMux I__4737 (
            .O(N__28306),
            .I(N__28300));
    LocalMux I__4736 (
            .O(N__28303),
            .I(N__28297));
    LocalMux I__4735 (
            .O(N__28300),
            .I(N__28294));
    Span4Mux_v I__4734 (
            .O(N__28297),
            .I(N__28290));
    Span4Mux_v I__4733 (
            .O(N__28294),
            .I(N__28287));
    InMux I__4732 (
            .O(N__28293),
            .I(N__28284));
    Sp12to4 I__4731 (
            .O(N__28290),
            .I(N__28279));
    Sp12to4 I__4730 (
            .O(N__28287),
            .I(N__28279));
    LocalMux I__4729 (
            .O(N__28284),
            .I(\pid_side.error_p_regZ0Z_19 ));
    Odrv12 I__4728 (
            .O(N__28279),
            .I(\pid_side.error_p_regZ0Z_19 ));
    InMux I__4727 (
            .O(N__28274),
            .I(N__28271));
    LocalMux I__4726 (
            .O(N__28271),
            .I(N__28268));
    Span4Mux_h I__4725 (
            .O(N__28268),
            .I(N__28264));
    InMux I__4724 (
            .O(N__28267),
            .I(N__28261));
    Sp12to4 I__4723 (
            .O(N__28264),
            .I(N__28255));
    LocalMux I__4722 (
            .O(N__28261),
            .I(N__28255));
    InMux I__4721 (
            .O(N__28260),
            .I(N__28252));
    Span12Mux_v I__4720 (
            .O(N__28255),
            .I(N__28249));
    LocalMux I__4719 (
            .O(N__28252),
            .I(\pid_side.error_p_regZ0Z_15 ));
    Odrv12 I__4718 (
            .O(N__28249),
            .I(\pid_side.error_p_regZ0Z_15 ));
    InMux I__4717 (
            .O(N__28244),
            .I(N__28241));
    LocalMux I__4716 (
            .O(N__28241),
            .I(\pid_side.un1_pid_prereg_cry_14_THRU_CO ));
    InMux I__4715 (
            .O(N__28238),
            .I(N__28235));
    LocalMux I__4714 (
            .O(N__28235),
            .I(N__28231));
    InMux I__4713 (
            .O(N__28234),
            .I(N__28228));
    Span4Mux_h I__4712 (
            .O(N__28231),
            .I(N__28223));
    LocalMux I__4711 (
            .O(N__28228),
            .I(N__28223));
    Span4Mux_h I__4710 (
            .O(N__28223),
            .I(N__28220));
    Span4Mux_h I__4709 (
            .O(N__28220),
            .I(N__28216));
    InMux I__4708 (
            .O(N__28219),
            .I(N__28213));
    Span4Mux_s1_h I__4707 (
            .O(N__28216),
            .I(N__28210));
    LocalMux I__4706 (
            .O(N__28213),
            .I(\pid_side.error_p_regZ0Z_14 ));
    Odrv4 I__4705 (
            .O(N__28210),
            .I(\pid_side.error_p_regZ0Z_14 ));
    InMux I__4704 (
            .O(N__28205),
            .I(N__28202));
    LocalMux I__4703 (
            .O(N__28202),
            .I(\pid_side.un1_pid_prereg_cry_13_THRU_CO ));
    InMux I__4702 (
            .O(N__28199),
            .I(N__28196));
    LocalMux I__4701 (
            .O(N__28196),
            .I(\pid_side.un1_pid_prereg_cry_16_THRU_CO ));
    InMux I__4700 (
            .O(N__28193),
            .I(N__28190));
    LocalMux I__4699 (
            .O(N__28190),
            .I(N__28186));
    InMux I__4698 (
            .O(N__28189),
            .I(N__28183));
    Span4Mux_v I__4697 (
            .O(N__28186),
            .I(N__28180));
    LocalMux I__4696 (
            .O(N__28183),
            .I(N__28177));
    Span4Mux_h I__4695 (
            .O(N__28180),
            .I(N__28173));
    Span4Mux_v I__4694 (
            .O(N__28177),
            .I(N__28170));
    InMux I__4693 (
            .O(N__28176),
            .I(N__28167));
    Span4Mux_h I__4692 (
            .O(N__28173),
            .I(N__28164));
    Span4Mux_h I__4691 (
            .O(N__28170),
            .I(N__28161));
    LocalMux I__4690 (
            .O(N__28167),
            .I(\pid_side.error_p_regZ0Z_17 ));
    Odrv4 I__4689 (
            .O(N__28164),
            .I(\pid_side.error_p_regZ0Z_17 ));
    Odrv4 I__4688 (
            .O(N__28161),
            .I(\pid_side.error_p_regZ0Z_17 ));
    InMux I__4687 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__4686 (
            .O(N__28151),
            .I(\pid_side.un1_pid_prereg_cry_19_THRU_CO ));
    InMux I__4685 (
            .O(N__28148),
            .I(N__28143));
    InMux I__4684 (
            .O(N__28147),
            .I(N__28138));
    InMux I__4683 (
            .O(N__28146),
            .I(N__28138));
    LocalMux I__4682 (
            .O(N__28143),
            .I(N__28132));
    LocalMux I__4681 (
            .O(N__28138),
            .I(N__28132));
    InMux I__4680 (
            .O(N__28137),
            .I(N__28129));
    Span4Mux_h I__4679 (
            .O(N__28132),
            .I(N__28126));
    LocalMux I__4678 (
            .O(N__28129),
            .I(\pid_side.error_p_regZ0Z_20 ));
    Odrv4 I__4677 (
            .O(N__28126),
            .I(\pid_side.error_p_regZ0Z_20 ));
    CascadeMux I__4676 (
            .O(N__28121),
            .I(N__28115));
    InMux I__4675 (
            .O(N__28120),
            .I(N__28109));
    InMux I__4674 (
            .O(N__28119),
            .I(N__28109));
    InMux I__4673 (
            .O(N__28118),
            .I(N__28102));
    InMux I__4672 (
            .O(N__28115),
            .I(N__28102));
    InMux I__4671 (
            .O(N__28114),
            .I(N__28102));
    LocalMux I__4670 (
            .O(N__28109),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    LocalMux I__4669 (
            .O(N__28102),
            .I(\dron_frame_decoder_1.stateZ0Z_4 ));
    InMux I__4668 (
            .O(N__28097),
            .I(N__28094));
    LocalMux I__4667 (
            .O(N__28094),
            .I(N__28091));
    Span4Mux_h I__4666 (
            .O(N__28091),
            .I(N__28088));
    Span4Mux_v I__4665 (
            .O(N__28088),
            .I(N__28085));
    Odrv4 I__4664 (
            .O(N__28085),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ));
    CascadeMux I__4663 (
            .O(N__28082),
            .I(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ));
    CascadeMux I__4662 (
            .O(N__28079),
            .I(N__28074));
    CascadeMux I__4661 (
            .O(N__28078),
            .I(N__28071));
    InMux I__4660 (
            .O(N__28077),
            .I(N__28066));
    InMux I__4659 (
            .O(N__28074),
            .I(N__28066));
    InMux I__4658 (
            .O(N__28071),
            .I(N__28063));
    LocalMux I__4657 (
            .O(N__28066),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    LocalMux I__4656 (
            .O(N__28063),
            .I(\dron_frame_decoder_1.stateZ0Z_7 ));
    InMux I__4655 (
            .O(N__28058),
            .I(N__28055));
    LocalMux I__4654 (
            .O(N__28055),
            .I(N__28047));
    InMux I__4653 (
            .O(N__28054),
            .I(N__28042));
    InMux I__4652 (
            .O(N__28053),
            .I(N__28042));
    InMux I__4651 (
            .O(N__28052),
            .I(N__28037));
    InMux I__4650 (
            .O(N__28051),
            .I(N__28037));
    InMux I__4649 (
            .O(N__28050),
            .I(N__28034));
    Odrv4 I__4648 (
            .O(N__28047),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__4647 (
            .O(N__28042),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__4646 (
            .O(N__28037),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    LocalMux I__4645 (
            .O(N__28034),
            .I(\dron_frame_decoder_1.stateZ0Z_6 ));
    InMux I__4644 (
            .O(N__28025),
            .I(N__28022));
    LocalMux I__4643 (
            .O(N__28022),
            .I(N__28019));
    Odrv4 I__4642 (
            .O(N__28019),
            .I(\dron_frame_decoder_1.N_412_4 ));
    CascadeMux I__4641 (
            .O(N__28016),
            .I(N__28013));
    InMux I__4640 (
            .O(N__28013),
            .I(N__28010));
    LocalMux I__4639 (
            .O(N__28010),
            .I(\dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0 ));
    InMux I__4638 (
            .O(N__28007),
            .I(N__28004));
    LocalMux I__4637 (
            .O(N__28004),
            .I(\dron_frame_decoder_1.N_175 ));
    InMux I__4636 (
            .O(N__28001),
            .I(N__27995));
    InMux I__4635 (
            .O(N__28000),
            .I(N__27990));
    InMux I__4634 (
            .O(N__27999),
            .I(N__27990));
    InMux I__4633 (
            .O(N__27998),
            .I(N__27987));
    LocalMux I__4632 (
            .O(N__27995),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    LocalMux I__4631 (
            .O(N__27990),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    LocalMux I__4630 (
            .O(N__27987),
            .I(\dron_frame_decoder_1.stateZ0Z_5 ));
    InMux I__4629 (
            .O(N__27980),
            .I(N__27977));
    LocalMux I__4628 (
            .O(N__27977),
            .I(N__27973));
    InMux I__4627 (
            .O(N__27976),
            .I(N__27970));
    Odrv4 I__4626 (
            .O(N__27973),
            .I(\dron_frame_decoder_1.N_431 ));
    LocalMux I__4625 (
            .O(N__27970),
            .I(\dron_frame_decoder_1.N_431 ));
    InMux I__4624 (
            .O(N__27965),
            .I(N__27960));
    InMux I__4623 (
            .O(N__27964),
            .I(N__27957));
    InMux I__4622 (
            .O(N__27963),
            .I(N__27954));
    LocalMux I__4621 (
            .O(N__27960),
            .I(\dron_frame_decoder_1.N_435 ));
    LocalMux I__4620 (
            .O(N__27957),
            .I(\dron_frame_decoder_1.N_435 ));
    LocalMux I__4619 (
            .O(N__27954),
            .I(\dron_frame_decoder_1.N_435 ));
    CascadeMux I__4618 (
            .O(N__27947),
            .I(N__27943));
    CascadeMux I__4617 (
            .O(N__27946),
            .I(N__27939));
    InMux I__4616 (
            .O(N__27943),
            .I(N__27936));
    InMux I__4615 (
            .O(N__27942),
            .I(N__27933));
    InMux I__4614 (
            .O(N__27939),
            .I(N__27930));
    LocalMux I__4613 (
            .O(N__27936),
            .I(N__27925));
    LocalMux I__4612 (
            .O(N__27933),
            .I(N__27925));
    LocalMux I__4611 (
            .O(N__27930),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    Odrv4 I__4610 (
            .O(N__27925),
            .I(\dron_frame_decoder_1.stateZ0Z_1 ));
    InMux I__4609 (
            .O(N__27920),
            .I(N__27917));
    LocalMux I__4608 (
            .O(N__27917),
            .I(N__27914));
    Span4Mux_h I__4607 (
            .O(N__27914),
            .I(N__27911));
    Odrv4 I__4606 (
            .O(N__27911),
            .I(\pid_side.un1_pid_prereg_cry_8_THRU_CO ));
    InMux I__4605 (
            .O(N__27908),
            .I(N__27904));
    CascadeMux I__4604 (
            .O(N__27907),
            .I(N__27901));
    LocalMux I__4603 (
            .O(N__27904),
            .I(N__27898));
    InMux I__4602 (
            .O(N__27901),
            .I(N__27895));
    Span4Mux_h I__4601 (
            .O(N__27898),
            .I(N__27889));
    LocalMux I__4600 (
            .O(N__27895),
            .I(N__27889));
    InMux I__4599 (
            .O(N__27894),
            .I(N__27886));
    Span4Mux_v I__4598 (
            .O(N__27889),
            .I(N__27883));
    LocalMux I__4597 (
            .O(N__27886),
            .I(N__27878));
    Span4Mux_h I__4596 (
            .O(N__27883),
            .I(N__27878));
    Odrv4 I__4595 (
            .O(N__27878),
            .I(\pid_side.error_p_regZ0Z_9 ));
    InMux I__4594 (
            .O(N__27875),
            .I(N__27863));
    InMux I__4593 (
            .O(N__27874),
            .I(N__27863));
    InMux I__4592 (
            .O(N__27873),
            .I(N__27863));
    InMux I__4591 (
            .O(N__27872),
            .I(N__27856));
    InMux I__4590 (
            .O(N__27871),
            .I(N__27856));
    InMux I__4589 (
            .O(N__27870),
            .I(N__27856));
    LocalMux I__4588 (
            .O(N__27863),
            .I(N__27849));
    LocalMux I__4587 (
            .O(N__27856),
            .I(N__27849));
    InMux I__4586 (
            .O(N__27855),
            .I(N__27844));
    InMux I__4585 (
            .O(N__27854),
            .I(N__27844));
    Odrv4 I__4584 (
            .O(N__27849),
            .I(\dron_frame_decoder_1.N_428 ));
    LocalMux I__4583 (
            .O(N__27844),
            .I(\dron_frame_decoder_1.N_428 ));
    CascadeMux I__4582 (
            .O(N__27839),
            .I(N__27836));
    InMux I__4581 (
            .O(N__27836),
            .I(N__27831));
    InMux I__4580 (
            .O(N__27835),
            .I(N__27828));
    CascadeMux I__4579 (
            .O(N__27834),
            .I(N__27825));
    LocalMux I__4578 (
            .O(N__27831),
            .I(N__27822));
    LocalMux I__4577 (
            .O(N__27828),
            .I(N__27819));
    InMux I__4576 (
            .O(N__27825),
            .I(N__27816));
    Span4Mux_v I__4575 (
            .O(N__27822),
            .I(N__27813));
    Odrv12 I__4574 (
            .O(N__27819),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    LocalMux I__4573 (
            .O(N__27816),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    Odrv4 I__4572 (
            .O(N__27813),
            .I(\dron_frame_decoder_1.stateZ0Z_3 ));
    CascadeMux I__4571 (
            .O(N__27806),
            .I(\dron_frame_decoder_1.N_412_4_cascade_ ));
    InMux I__4570 (
            .O(N__27803),
            .I(N__27798));
    InMux I__4569 (
            .O(N__27802),
            .I(N__27795));
    InMux I__4568 (
            .O(N__27801),
            .I(N__27792));
    LocalMux I__4567 (
            .O(N__27798),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__4566 (
            .O(N__27795),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    LocalMux I__4565 (
            .O(N__27792),
            .I(\dron_frame_decoder_1.WDTZ0Z_15 ));
    CascadeMux I__4564 (
            .O(N__27785),
            .I(N__27781));
    InMux I__4563 (
            .O(N__27784),
            .I(N__27777));
    InMux I__4562 (
            .O(N__27781),
            .I(N__27774));
    InMux I__4561 (
            .O(N__27780),
            .I(N__27771));
    LocalMux I__4560 (
            .O(N__27777),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__4559 (
            .O(N__27774),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    LocalMux I__4558 (
            .O(N__27771),
            .I(\dron_frame_decoder_1.WDTZ0Z_14 ));
    InMux I__4557 (
            .O(N__27764),
            .I(N__27761));
    LocalMux I__4556 (
            .O(N__27761),
            .I(N__27758));
    Odrv4 I__4555 (
            .O(N__27758),
            .I(\dron_frame_decoder_1.WDT10lt14_0 ));
    CascadeMux I__4554 (
            .O(N__27755),
            .I(\dron_frame_decoder_1.N_177_cascade_ ));
    InMux I__4553 (
            .O(N__27752),
            .I(N__27746));
    InMux I__4552 (
            .O(N__27751),
            .I(N__27743));
    InMux I__4551 (
            .O(N__27750),
            .I(N__27740));
    InMux I__4550 (
            .O(N__27749),
            .I(N__27737));
    LocalMux I__4549 (
            .O(N__27746),
            .I(N__27734));
    LocalMux I__4548 (
            .O(N__27743),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__4547 (
            .O(N__27740),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    LocalMux I__4546 (
            .O(N__27737),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    Odrv4 I__4545 (
            .O(N__27734),
            .I(\dron_frame_decoder_1.stateZ0Z_0 ));
    InMux I__4544 (
            .O(N__27725),
            .I(N__27722));
    LocalMux I__4543 (
            .O(N__27722),
            .I(\dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3 ));
    CascadeMux I__4542 (
            .O(N__27719),
            .I(N__27716));
    InMux I__4541 (
            .O(N__27716),
            .I(N__27710));
    InMux I__4540 (
            .O(N__27715),
            .I(N__27710));
    LocalMux I__4539 (
            .O(N__27710),
            .I(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ));
    InMux I__4538 (
            .O(N__27707),
            .I(\scaler_4.un2_source_data_0_cry_3 ));
    CascadeMux I__4537 (
            .O(N__27704),
            .I(N__27701));
    InMux I__4536 (
            .O(N__27701),
            .I(N__27695));
    InMux I__4535 (
            .O(N__27700),
            .I(N__27695));
    LocalMux I__4534 (
            .O(N__27695),
            .I(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ));
    InMux I__4533 (
            .O(N__27692),
            .I(\scaler_4.un2_source_data_0_cry_4 ));
    CascadeMux I__4532 (
            .O(N__27689),
            .I(N__27686));
    InMux I__4531 (
            .O(N__27686),
            .I(N__27680));
    InMux I__4530 (
            .O(N__27685),
            .I(N__27680));
    LocalMux I__4529 (
            .O(N__27680),
            .I(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ));
    InMux I__4528 (
            .O(N__27677),
            .I(\scaler_4.un2_source_data_0_cry_5 ));
    CascadeMux I__4527 (
            .O(N__27674),
            .I(N__27671));
    InMux I__4526 (
            .O(N__27671),
            .I(N__27665));
    InMux I__4525 (
            .O(N__27670),
            .I(N__27665));
    LocalMux I__4524 (
            .O(N__27665),
            .I(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ));
    InMux I__4523 (
            .O(N__27662),
            .I(\scaler_4.un2_source_data_0_cry_6 ));
    CascadeMux I__4522 (
            .O(N__27659),
            .I(N__27656));
    InMux I__4521 (
            .O(N__27656),
            .I(N__27650));
    InMux I__4520 (
            .O(N__27655),
            .I(N__27650));
    LocalMux I__4519 (
            .O(N__27650),
            .I(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ));
    InMux I__4518 (
            .O(N__27647),
            .I(\scaler_4.un2_source_data_0_cry_7 ));
    InMux I__4517 (
            .O(N__27644),
            .I(N__27640));
    InMux I__4516 (
            .O(N__27643),
            .I(N__27637));
    LocalMux I__4515 (
            .O(N__27640),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    LocalMux I__4514 (
            .O(N__27637),
            .I(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ));
    CascadeMux I__4513 (
            .O(N__27632),
            .I(N__27629));
    InMux I__4512 (
            .O(N__27629),
            .I(N__27626));
    LocalMux I__4511 (
            .O(N__27626),
            .I(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ));
    InMux I__4510 (
            .O(N__27623),
            .I(bfn_9_11_0_));
    InMux I__4509 (
            .O(N__27620),
            .I(\scaler_4.un2_source_data_0_cry_9 ));
    CascadeMux I__4508 (
            .O(N__27617),
            .I(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ));
    InMux I__4507 (
            .O(N__27614),
            .I(N__27594));
    InMux I__4506 (
            .O(N__27613),
            .I(N__27591));
    InMux I__4505 (
            .O(N__27612),
            .I(N__27588));
    InMux I__4504 (
            .O(N__27611),
            .I(N__27585));
    InMux I__4503 (
            .O(N__27610),
            .I(N__27582));
    InMux I__4502 (
            .O(N__27609),
            .I(N__27579));
    CascadeMux I__4501 (
            .O(N__27608),
            .I(N__27574));
    InMux I__4500 (
            .O(N__27607),
            .I(N__27569));
    InMux I__4499 (
            .O(N__27606),
            .I(N__27569));
    InMux I__4498 (
            .O(N__27605),
            .I(N__27564));
    InMux I__4497 (
            .O(N__27604),
            .I(N__27551));
    InMux I__4496 (
            .O(N__27603),
            .I(N__27551));
    InMux I__4495 (
            .O(N__27602),
            .I(N__27551));
    InMux I__4494 (
            .O(N__27601),
            .I(N__27551));
    InMux I__4493 (
            .O(N__27600),
            .I(N__27551));
    InMux I__4492 (
            .O(N__27599),
            .I(N__27551));
    InMux I__4491 (
            .O(N__27598),
            .I(N__27546));
    InMux I__4490 (
            .O(N__27597),
            .I(N__27546));
    LocalMux I__4489 (
            .O(N__27594),
            .I(N__27541));
    LocalMux I__4488 (
            .O(N__27591),
            .I(N__27541));
    LocalMux I__4487 (
            .O(N__27588),
            .I(N__27538));
    LocalMux I__4486 (
            .O(N__27585),
            .I(N__27530));
    LocalMux I__4485 (
            .O(N__27582),
            .I(N__27530));
    LocalMux I__4484 (
            .O(N__27579),
            .I(N__27527));
    InMux I__4483 (
            .O(N__27578),
            .I(N__27524));
    InMux I__4482 (
            .O(N__27577),
            .I(N__27519));
    InMux I__4481 (
            .O(N__27574),
            .I(N__27519));
    LocalMux I__4480 (
            .O(N__27569),
            .I(N__27516));
    InMux I__4479 (
            .O(N__27568),
            .I(N__27511));
    InMux I__4478 (
            .O(N__27567),
            .I(N__27511));
    LocalMux I__4477 (
            .O(N__27564),
            .I(N__27508));
    LocalMux I__4476 (
            .O(N__27551),
            .I(N__27505));
    LocalMux I__4475 (
            .O(N__27546),
            .I(N__27498));
    Span4Mux_h I__4474 (
            .O(N__27541),
            .I(N__27498));
    Span4Mux_h I__4473 (
            .O(N__27538),
            .I(N__27498));
    InMux I__4472 (
            .O(N__27537),
            .I(N__27495));
    InMux I__4471 (
            .O(N__27536),
            .I(N__27492));
    InMux I__4470 (
            .O(N__27535),
            .I(N__27488));
    Span12Mux_v I__4469 (
            .O(N__27530),
            .I(N__27485));
    Span4Mux_h I__4468 (
            .O(N__27527),
            .I(N__27478));
    LocalMux I__4467 (
            .O(N__27524),
            .I(N__27478));
    LocalMux I__4466 (
            .O(N__27519),
            .I(N__27478));
    Span4Mux_v I__4465 (
            .O(N__27516),
            .I(N__27471));
    LocalMux I__4464 (
            .O(N__27511),
            .I(N__27471));
    Span4Mux_v I__4463 (
            .O(N__27508),
            .I(N__27471));
    Span4Mux_v I__4462 (
            .O(N__27505),
            .I(N__27468));
    Span4Mux_v I__4461 (
            .O(N__27498),
            .I(N__27461));
    LocalMux I__4460 (
            .O(N__27495),
            .I(N__27461));
    LocalMux I__4459 (
            .O(N__27492),
            .I(N__27461));
    InMux I__4458 (
            .O(N__27491),
            .I(N__27458));
    LocalMux I__4457 (
            .O(N__27488),
            .I(uart_pc_data_rdy));
    Odrv12 I__4456 (
            .O(N__27485),
            .I(uart_pc_data_rdy));
    Odrv4 I__4455 (
            .O(N__27478),
            .I(uart_pc_data_rdy));
    Odrv4 I__4454 (
            .O(N__27471),
            .I(uart_pc_data_rdy));
    Odrv4 I__4453 (
            .O(N__27468),
            .I(uart_pc_data_rdy));
    Odrv4 I__4452 (
            .O(N__27461),
            .I(uart_pc_data_rdy));
    LocalMux I__4451 (
            .O(N__27458),
            .I(uart_pc_data_rdy));
    CascadeMux I__4450 (
            .O(N__27443),
            .I(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ));
    InMux I__4449 (
            .O(N__27440),
            .I(N__27435));
    InMux I__4448 (
            .O(N__27439),
            .I(N__27430));
    InMux I__4447 (
            .O(N__27438),
            .I(N__27430));
    LocalMux I__4446 (
            .O(N__27435),
            .I(N__27425));
    LocalMux I__4445 (
            .O(N__27430),
            .I(N__27425));
    Odrv12 I__4444 (
            .O(N__27425),
            .I(\Commands_frame_decoder.N_422 ));
    InMux I__4443 (
            .O(N__27422),
            .I(N__27416));
    InMux I__4442 (
            .O(N__27421),
            .I(N__27413));
    InMux I__4441 (
            .O(N__27420),
            .I(N__27410));
    InMux I__4440 (
            .O(N__27419),
            .I(N__27407));
    LocalMux I__4439 (
            .O(N__27416),
            .I(N__27403));
    LocalMux I__4438 (
            .O(N__27413),
            .I(N__27400));
    LocalMux I__4437 (
            .O(N__27410),
            .I(N__27397));
    LocalMux I__4436 (
            .O(N__27407),
            .I(N__27394));
    InMux I__4435 (
            .O(N__27406),
            .I(N__27391));
    Span12Mux_v I__4434 (
            .O(N__27403),
            .I(N__27386));
    Span4Mux_h I__4433 (
            .O(N__27400),
            .I(N__27383));
    Span4Mux_h I__4432 (
            .O(N__27397),
            .I(N__27376));
    Span4Mux_v I__4431 (
            .O(N__27394),
            .I(N__27376));
    LocalMux I__4430 (
            .O(N__27391),
            .I(N__27376));
    InMux I__4429 (
            .O(N__27390),
            .I(N__27371));
    InMux I__4428 (
            .O(N__27389),
            .I(N__27371));
    Odrv12 I__4427 (
            .O(N__27386),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__4426 (
            .O(N__27383),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    Odrv4 I__4425 (
            .O(N__27376),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    LocalMux I__4424 (
            .O(N__27371),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ));
    CascadeMux I__4423 (
            .O(N__27362),
            .I(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ));
    CascadeMux I__4422 (
            .O(N__27359),
            .I(N__27355));
    InMux I__4421 (
            .O(N__27358),
            .I(N__27352));
    InMux I__4420 (
            .O(N__27355),
            .I(N__27349));
    LocalMux I__4419 (
            .O(N__27352),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    LocalMux I__4418 (
            .O(N__27349),
            .I(\uart_pc.data_AuxZ0Z_4 ));
    CascadeMux I__4417 (
            .O(N__27344),
            .I(N__27341));
    InMux I__4416 (
            .O(N__27341),
            .I(N__27338));
    LocalMux I__4415 (
            .O(N__27338),
            .I(N__27335));
    Span4Mux_v I__4414 (
            .O(N__27335),
            .I(N__27331));
    InMux I__4413 (
            .O(N__27334),
            .I(N__27328));
    Odrv4 I__4412 (
            .O(N__27331),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    LocalMux I__4411 (
            .O(N__27328),
            .I(\uart_pc.data_AuxZ1Z_0 ));
    CascadeMux I__4410 (
            .O(N__27323),
            .I(N__27320));
    InMux I__4409 (
            .O(N__27320),
            .I(N__27317));
    LocalMux I__4408 (
            .O(N__27317),
            .I(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ));
    InMux I__4407 (
            .O(N__27314),
            .I(\scaler_4.un2_source_data_0_cry_1 ));
    CascadeMux I__4406 (
            .O(N__27311),
            .I(N__27308));
    InMux I__4405 (
            .O(N__27308),
            .I(N__27302));
    InMux I__4404 (
            .O(N__27307),
            .I(N__27302));
    LocalMux I__4403 (
            .O(N__27302),
            .I(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ));
    InMux I__4402 (
            .O(N__27299),
            .I(\scaler_4.un2_source_data_0_cry_2 ));
    InMux I__4401 (
            .O(N__27296),
            .I(N__27293));
    LocalMux I__4400 (
            .O(N__27293),
            .I(uart_input_pc_c));
    InMux I__4399 (
            .O(N__27290),
            .I(N__27287));
    LocalMux I__4398 (
            .O(N__27287),
            .I(\uart_pc_sync.aux_0__0_Z0Z_0 ));
    InMux I__4397 (
            .O(N__27284),
            .I(N__27281));
    LocalMux I__4396 (
            .O(N__27281),
            .I(\uart_pc_sync.aux_1__0_Z0Z_0 ));
    InMux I__4395 (
            .O(N__27278),
            .I(N__27275));
    LocalMux I__4394 (
            .O(N__27275),
            .I(\uart_pc_sync.aux_2__0_Z0Z_0 ));
    InMux I__4393 (
            .O(N__27272),
            .I(N__27269));
    LocalMux I__4392 (
            .O(N__27269),
            .I(\uart_pc_sync.aux_3__0_Z0Z_0 ));
    InMux I__4391 (
            .O(N__27266),
            .I(N__27262));
    InMux I__4390 (
            .O(N__27265),
            .I(N__27259));
    LocalMux I__4389 (
            .O(N__27262),
            .I(N__27256));
    LocalMux I__4388 (
            .O(N__27259),
            .I(N__27251));
    Span4Mux_h I__4387 (
            .O(N__27256),
            .I(N__27248));
    InMux I__4386 (
            .O(N__27255),
            .I(N__27245));
    InMux I__4385 (
            .O(N__27254),
            .I(N__27242));
    Span4Mux_h I__4384 (
            .O(N__27251),
            .I(N__27239));
    Odrv4 I__4383 (
            .O(N__27248),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__4382 (
            .O(N__27245),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    LocalMux I__4381 (
            .O(N__27242),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    Odrv4 I__4380 (
            .O(N__27239),
            .I(\Commands_frame_decoder.stateZ0Z_14 ));
    InMux I__4379 (
            .O(N__27230),
            .I(N__27226));
    CascadeMux I__4378 (
            .O(N__27229),
            .I(N__27223));
    LocalMux I__4377 (
            .O(N__27226),
            .I(N__27220));
    InMux I__4376 (
            .O(N__27223),
            .I(N__27216));
    Span4Mux_v I__4375 (
            .O(N__27220),
            .I(N__27213));
    InMux I__4374 (
            .O(N__27219),
            .I(N__27210));
    LocalMux I__4373 (
            .O(N__27216),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    Odrv4 I__4372 (
            .O(N__27213),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    LocalMux I__4371 (
            .O(N__27210),
            .I(\Commands_frame_decoder.countZ0Z_0 ));
    IoInMux I__4370 (
            .O(N__27203),
            .I(N__27200));
    LocalMux I__4369 (
            .O(N__27200),
            .I(N__27197));
    Span4Mux_s1_v I__4368 (
            .O(N__27197),
            .I(N__27194));
    Span4Mux_v I__4367 (
            .O(N__27194),
            .I(N__27190));
    InMux I__4366 (
            .O(N__27193),
            .I(N__27187));
    Span4Mux_h I__4365 (
            .O(N__27190),
            .I(N__27183));
    LocalMux I__4364 (
            .O(N__27187),
            .I(N__27180));
    CascadeMux I__4363 (
            .O(N__27186),
            .I(N__27177));
    Span4Mux_h I__4362 (
            .O(N__27183),
            .I(N__27171));
    Span4Mux_v I__4361 (
            .O(N__27180),
            .I(N__27171));
    InMux I__4360 (
            .O(N__27177),
            .I(N__27168));
    InMux I__4359 (
            .O(N__27176),
            .I(N__27165));
    Odrv4 I__4358 (
            .O(N__27171),
            .I(debug_CH3_20A_c));
    LocalMux I__4357 (
            .O(N__27168),
            .I(debug_CH3_20A_c));
    LocalMux I__4356 (
            .O(N__27165),
            .I(debug_CH3_20A_c));
    InMux I__4355 (
            .O(N__27158),
            .I(N__27155));
    LocalMux I__4354 (
            .O(N__27155),
            .I(N__27151));
    InMux I__4353 (
            .O(N__27154),
            .I(N__27148));
    Span12Mux_s8_h I__4352 (
            .O(N__27151),
            .I(N__27145));
    LocalMux I__4351 (
            .O(N__27148),
            .I(N__27142));
    Odrv12 I__4350 (
            .O(N__27145),
            .I(drone_H_disp_side_0));
    Odrv12 I__4349 (
            .O(N__27142),
            .I(drone_H_disp_side_0));
    InMux I__4348 (
            .O(N__27137),
            .I(N__27134));
    LocalMux I__4347 (
            .O(N__27134),
            .I(drone_H_disp_side_2));
    InMux I__4346 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__4345 (
            .O(N__27128),
            .I(drone_H_disp_side_3));
    InMux I__4344 (
            .O(N__27125),
            .I(N__27122));
    LocalMux I__4343 (
            .O(N__27122),
            .I(\dron_frame_decoder_1.drone_H_disp_side_4 ));
    InMux I__4342 (
            .O(N__27119),
            .I(N__27116));
    LocalMux I__4341 (
            .O(N__27116),
            .I(\dron_frame_decoder_1.drone_H_disp_side_5 ));
    InMux I__4340 (
            .O(N__27113),
            .I(N__27110));
    LocalMux I__4339 (
            .O(N__27110),
            .I(N__27107));
    Odrv4 I__4338 (
            .O(N__27107),
            .I(\dron_frame_decoder_1.drone_H_disp_side_6 ));
    InMux I__4337 (
            .O(N__27104),
            .I(N__27101));
    LocalMux I__4336 (
            .O(N__27101),
            .I(\dron_frame_decoder_1.drone_H_disp_side_7 ));
    CEMux I__4335 (
            .O(N__27098),
            .I(N__27095));
    LocalMux I__4334 (
            .O(N__27095),
            .I(N__27092));
    Odrv12 I__4333 (
            .O(N__27092),
            .I(\dron_frame_decoder_1.N_747_0 ));
    InMux I__4332 (
            .O(N__27089),
            .I(N__27086));
    LocalMux I__4331 (
            .O(N__27086),
            .I(N__27083));
    Span4Mux_s1_h I__4330 (
            .O(N__27083),
            .I(N__27080));
    Sp12to4 I__4329 (
            .O(N__27080),
            .I(N__27077));
    Span12Mux_v I__4328 (
            .O(N__27077),
            .I(N__27074));
    Odrv12 I__4327 (
            .O(N__27074),
            .I(alt_ki_7));
    InMux I__4326 (
            .O(N__27071),
            .I(\pid_side.un1_pid_prereg_cry_13 ));
    InMux I__4325 (
            .O(N__27068),
            .I(\pid_side.un1_pid_prereg_cry_14 ));
    InMux I__4324 (
            .O(N__27065),
            .I(\pid_side.un1_pid_prereg_cry_15 ));
    InMux I__4323 (
            .O(N__27062),
            .I(bfn_8_19_0_));
    InMux I__4322 (
            .O(N__27059),
            .I(\pid_side.un1_pid_prereg_cry_17 ));
    InMux I__4321 (
            .O(N__27056),
            .I(\pid_side.un1_pid_prereg_cry_18 ));
    InMux I__4320 (
            .O(N__27053),
            .I(\pid_side.un1_pid_prereg_cry_19 ));
    InMux I__4319 (
            .O(N__27050),
            .I(\pid_side.un1_pid_prereg_cry_20 ));
    CEMux I__4318 (
            .O(N__27047),
            .I(N__27044));
    LocalMux I__4317 (
            .O(N__27044),
            .I(N__27041));
    Span4Mux_v I__4316 (
            .O(N__27041),
            .I(N__27038));
    Span4Mux_h I__4315 (
            .O(N__27038),
            .I(N__27034));
    CEMux I__4314 (
            .O(N__27037),
            .I(N__27031));
    Odrv4 I__4313 (
            .O(N__27034),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    LocalMux I__4312 (
            .O(N__27031),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ));
    InMux I__4311 (
            .O(N__27026),
            .I(\pid_side.un1_pid_prereg_cry_4 ));
    InMux I__4310 (
            .O(N__27023),
            .I(\pid_side.un1_pid_prereg_cry_5 ));
    InMux I__4309 (
            .O(N__27020),
            .I(\pid_side.un1_pid_prereg_cry_6 ));
    InMux I__4308 (
            .O(N__27017),
            .I(\pid_side.un1_pid_prereg_cry_7 ));
    InMux I__4307 (
            .O(N__27014),
            .I(bfn_8_18_0_));
    InMux I__4306 (
            .O(N__27011),
            .I(\pid_side.un1_pid_prereg_cry_9 ));
    InMux I__4305 (
            .O(N__27008),
            .I(\pid_side.un1_pid_prereg_cry_10 ));
    InMux I__4304 (
            .O(N__27005),
            .I(\pid_side.un1_pid_prereg_cry_11 ));
    InMux I__4303 (
            .O(N__27002),
            .I(\pid_side.un1_pid_prereg_cry_12 ));
    CascadeMux I__4302 (
            .O(N__26999),
            .I(N__26995));
    CascadeMux I__4301 (
            .O(N__26998),
            .I(N__26992));
    InMux I__4300 (
            .O(N__26995),
            .I(N__26987));
    InMux I__4299 (
            .O(N__26992),
            .I(N__26980));
    InMux I__4298 (
            .O(N__26991),
            .I(N__26980));
    InMux I__4297 (
            .O(N__26990),
            .I(N__26980));
    LocalMux I__4296 (
            .O(N__26987),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    LocalMux I__4295 (
            .O(N__26980),
            .I(\Commands_frame_decoder.stateZ0Z_7 ));
    CascadeMux I__4294 (
            .O(N__26975),
            .I(N__26971));
    InMux I__4293 (
            .O(N__26974),
            .I(N__26966));
    InMux I__4292 (
            .O(N__26971),
            .I(N__26966));
    LocalMux I__4291 (
            .O(N__26966),
            .I(\Commands_frame_decoder.stateZ0Z_8 ));
    CEMux I__4290 (
            .O(N__26963),
            .I(N__26960));
    LocalMux I__4289 (
            .O(N__26960),
            .I(N__26957));
    Span4Mux_v I__4288 (
            .O(N__26957),
            .I(N__26953));
    CEMux I__4287 (
            .O(N__26956),
            .I(N__26950));
    Span4Mux_h I__4286 (
            .O(N__26953),
            .I(N__26947));
    LocalMux I__4285 (
            .O(N__26950),
            .I(N__26944));
    Span4Mux_h I__4284 (
            .O(N__26947),
            .I(N__26939));
    Span4Mux_v I__4283 (
            .O(N__26944),
            .I(N__26939));
    Odrv4 I__4282 (
            .O(N__26939),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ));
    InMux I__4281 (
            .O(N__26936),
            .I(N__26930));
    InMux I__4280 (
            .O(N__26935),
            .I(N__26930));
    LocalMux I__4279 (
            .O(N__26930),
            .I(\Commands_frame_decoder.stateZ0Z_9 ));
    InMux I__4278 (
            .O(N__26927),
            .I(N__26924));
    LocalMux I__4277 (
            .O(N__26924),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa ));
    CascadeMux I__4276 (
            .O(N__26921),
            .I(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ));
    InMux I__4275 (
            .O(N__26918),
            .I(N__26904));
    InMux I__4274 (
            .O(N__26917),
            .I(N__26904));
    InMux I__4273 (
            .O(N__26916),
            .I(N__26904));
    InMux I__4272 (
            .O(N__26915),
            .I(N__26904));
    InMux I__4271 (
            .O(N__26914),
            .I(N__26898));
    InMux I__4270 (
            .O(N__26913),
            .I(N__26895));
    LocalMux I__4269 (
            .O(N__26904),
            .I(N__26890));
    InMux I__4268 (
            .O(N__26903),
            .I(N__26887));
    InMux I__4267 (
            .O(N__26902),
            .I(N__26884));
    InMux I__4266 (
            .O(N__26901),
            .I(N__26881));
    LocalMux I__4265 (
            .O(N__26898),
            .I(N__26876));
    LocalMux I__4264 (
            .O(N__26895),
            .I(N__26873));
    InMux I__4263 (
            .O(N__26894),
            .I(N__26868));
    InMux I__4262 (
            .O(N__26893),
            .I(N__26868));
    Span4Mux_v I__4261 (
            .O(N__26890),
            .I(N__26865));
    LocalMux I__4260 (
            .O(N__26887),
            .I(N__26860));
    LocalMux I__4259 (
            .O(N__26884),
            .I(N__26860));
    LocalMux I__4258 (
            .O(N__26881),
            .I(N__26857));
    InMux I__4257 (
            .O(N__26880),
            .I(N__26852));
    InMux I__4256 (
            .O(N__26879),
            .I(N__26852));
    Span4Mux_v I__4255 (
            .O(N__26876),
            .I(N__26844));
    Span4Mux_h I__4254 (
            .O(N__26873),
            .I(N__26844));
    LocalMux I__4253 (
            .O(N__26868),
            .I(N__26844));
    Span4Mux_v I__4252 (
            .O(N__26865),
            .I(N__26835));
    Span4Mux_v I__4251 (
            .O(N__26860),
            .I(N__26835));
    Span4Mux_h I__4250 (
            .O(N__26857),
            .I(N__26835));
    LocalMux I__4249 (
            .O(N__26852),
            .I(N__26835));
    InMux I__4248 (
            .O(N__26851),
            .I(N__26832));
    Odrv4 I__4247 (
            .O(N__26844),
            .I(\Commands_frame_decoder.N_415 ));
    Odrv4 I__4246 (
            .O(N__26835),
            .I(\Commands_frame_decoder.N_415 ));
    LocalMux I__4245 (
            .O(N__26832),
            .I(\Commands_frame_decoder.N_415 ));
    CascadeMux I__4244 (
            .O(N__26825),
            .I(N__26822));
    InMux I__4243 (
            .O(N__26822),
            .I(N__26819));
    LocalMux I__4242 (
            .O(N__26819),
            .I(N__26815));
    InMux I__4241 (
            .O(N__26818),
            .I(N__26812));
    Span4Mux_h I__4240 (
            .O(N__26815),
            .I(N__26808));
    LocalMux I__4239 (
            .O(N__26812),
            .I(N__26805));
    InMux I__4238 (
            .O(N__26811),
            .I(N__26802));
    Span4Mux_v I__4237 (
            .O(N__26808),
            .I(N__26799));
    Span12Mux_s8_h I__4236 (
            .O(N__26805),
            .I(N__26796));
    LocalMux I__4235 (
            .O(N__26802),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv4 I__4234 (
            .O(N__26799),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    Odrv12 I__4233 (
            .O(N__26796),
            .I(\Commands_frame_decoder.stateZ0Z_10 ));
    InMux I__4232 (
            .O(N__26789),
            .I(\pid_side.un1_pid_prereg_cry_1 ));
    InMux I__4231 (
            .O(N__26786),
            .I(\pid_side.un1_pid_prereg_cry_2 ));
    InMux I__4230 (
            .O(N__26783),
            .I(\pid_side.un1_pid_prereg_cry_3 ));
    InMux I__4229 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__4228 (
            .O(N__26777),
            .I(N__26774));
    Span4Mux_v I__4227 (
            .O(N__26774),
            .I(N__26771));
    Odrv4 I__4226 (
            .O(N__26771),
            .I(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ));
    CascadeMux I__4225 (
            .O(N__26768),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_ ));
    InMux I__4224 (
            .O(N__26765),
            .I(N__26759));
    InMux I__4223 (
            .O(N__26764),
            .I(N__26759));
    LocalMux I__4222 (
            .O(N__26759),
            .I(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0 ));
    InMux I__4221 (
            .O(N__26756),
            .I(N__26752));
    InMux I__4220 (
            .O(N__26755),
            .I(N__26749));
    LocalMux I__4219 (
            .O(N__26752),
            .I(N__26746));
    LocalMux I__4218 (
            .O(N__26749),
            .I(N__26742));
    Span12Mux_s5_h I__4217 (
            .O(N__26746),
            .I(N__26739));
    InMux I__4216 (
            .O(N__26745),
            .I(N__26736));
    Span4Mux_s3_h I__4215 (
            .O(N__26742),
            .I(N__26733));
    Span12Mux_h I__4214 (
            .O(N__26739),
            .I(N__26730));
    LocalMux I__4213 (
            .O(N__26736),
            .I(N__26725));
    Span4Mux_h I__4212 (
            .O(N__26733),
            .I(N__26725));
    Odrv12 I__4211 (
            .O(N__26730),
            .I(xy_kp_4));
    Odrv4 I__4210 (
            .O(N__26725),
            .I(xy_kp_4));
    CascadeMux I__4209 (
            .O(N__26720),
            .I(N__26716));
    CascadeMux I__4208 (
            .O(N__26719),
            .I(N__26713));
    InMux I__4207 (
            .O(N__26716),
            .I(N__26709));
    InMux I__4206 (
            .O(N__26713),
            .I(N__26706));
    InMux I__4205 (
            .O(N__26712),
            .I(N__26703));
    LocalMux I__4204 (
            .O(N__26709),
            .I(N__26699));
    LocalMux I__4203 (
            .O(N__26706),
            .I(N__26694));
    LocalMux I__4202 (
            .O(N__26703),
            .I(N__26694));
    InMux I__4201 (
            .O(N__26702),
            .I(N__26691));
    Span4Mux_v I__4200 (
            .O(N__26699),
            .I(N__26688));
    Span12Mux_s10_v I__4199 (
            .O(N__26694),
            .I(N__26685));
    LocalMux I__4198 (
            .O(N__26691),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv4 I__4197 (
            .O(N__26688),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    Odrv12 I__4196 (
            .O(N__26685),
            .I(\Commands_frame_decoder.stateZ0Z_6 ));
    InMux I__4195 (
            .O(N__26678),
            .I(N__26673));
    InMux I__4194 (
            .O(N__26677),
            .I(N__26668));
    InMux I__4193 (
            .O(N__26676),
            .I(N__26668));
    LocalMux I__4192 (
            .O(N__26673),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    LocalMux I__4191 (
            .O(N__26668),
            .I(\dron_frame_decoder_1.WDTZ0Z_12 ));
    InMux I__4190 (
            .O(N__26663),
            .I(\dron_frame_decoder_1.un1_WDT_cry_11 ));
    CascadeMux I__4189 (
            .O(N__26660),
            .I(N__26656));
    InMux I__4188 (
            .O(N__26659),
            .I(N__26653));
    InMux I__4187 (
            .O(N__26656),
            .I(N__26650));
    LocalMux I__4186 (
            .O(N__26653),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    LocalMux I__4185 (
            .O(N__26650),
            .I(\dron_frame_decoder_1.WDTZ0Z_13 ));
    InMux I__4184 (
            .O(N__26645),
            .I(\dron_frame_decoder_1.un1_WDT_cry_12 ));
    InMux I__4183 (
            .O(N__26642),
            .I(\dron_frame_decoder_1.un1_WDT_cry_13 ));
    InMux I__4182 (
            .O(N__26639),
            .I(\dron_frame_decoder_1.un1_WDT_cry_14 ));
    CascadeMux I__4181 (
            .O(N__26636),
            .I(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ));
    SRMux I__4180 (
            .O(N__26633),
            .I(N__26630));
    LocalMux I__4179 (
            .O(N__26630),
            .I(N__26627));
    Span4Mux_h I__4178 (
            .O(N__26627),
            .I(N__26624));
    Span4Mux_h I__4177 (
            .O(N__26624),
            .I(N__26620));
    SRMux I__4176 (
            .O(N__26623),
            .I(N__26617));
    Odrv4 I__4175 (
            .O(N__26620),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    LocalMux I__4174 (
            .O(N__26617),
            .I(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ));
    InMux I__4173 (
            .O(N__26612),
            .I(N__26609));
    LocalMux I__4172 (
            .O(N__26609),
            .I(\dron_frame_decoder_1.WDTZ0Z_3 ));
    InMux I__4171 (
            .O(N__26606),
            .I(\dron_frame_decoder_1.un1_WDT_cry_2 ));
    CascadeMux I__4170 (
            .O(N__26603),
            .I(N__26599));
    InMux I__4169 (
            .O(N__26602),
            .I(N__26596));
    InMux I__4168 (
            .O(N__26599),
            .I(N__26593));
    LocalMux I__4167 (
            .O(N__26596),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    LocalMux I__4166 (
            .O(N__26593),
            .I(\dron_frame_decoder_1.WDTZ0Z_4 ));
    InMux I__4165 (
            .O(N__26588),
            .I(\dron_frame_decoder_1.un1_WDT_cry_3 ));
    InMux I__4164 (
            .O(N__26585),
            .I(N__26581));
    InMux I__4163 (
            .O(N__26584),
            .I(N__26578));
    LocalMux I__4162 (
            .O(N__26581),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    LocalMux I__4161 (
            .O(N__26578),
            .I(\dron_frame_decoder_1.WDTZ0Z_5 ));
    InMux I__4160 (
            .O(N__26573),
            .I(\dron_frame_decoder_1.un1_WDT_cry_4 ));
    InMux I__4159 (
            .O(N__26570),
            .I(N__26566));
    InMux I__4158 (
            .O(N__26569),
            .I(N__26563));
    LocalMux I__4157 (
            .O(N__26566),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    LocalMux I__4156 (
            .O(N__26563),
            .I(\dron_frame_decoder_1.WDTZ0Z_6 ));
    InMux I__4155 (
            .O(N__26558),
            .I(\dron_frame_decoder_1.un1_WDT_cry_5 ));
    InMux I__4154 (
            .O(N__26555),
            .I(N__26551));
    InMux I__4153 (
            .O(N__26554),
            .I(N__26548));
    LocalMux I__4152 (
            .O(N__26551),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    LocalMux I__4151 (
            .O(N__26548),
            .I(\dron_frame_decoder_1.WDTZ0Z_7 ));
    InMux I__4150 (
            .O(N__26543),
            .I(\dron_frame_decoder_1.un1_WDT_cry_6 ));
    InMux I__4149 (
            .O(N__26540),
            .I(N__26536));
    InMux I__4148 (
            .O(N__26539),
            .I(N__26533));
    LocalMux I__4147 (
            .O(N__26536),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    LocalMux I__4146 (
            .O(N__26533),
            .I(\dron_frame_decoder_1.WDTZ0Z_8 ));
    InMux I__4145 (
            .O(N__26528),
            .I(bfn_8_12_0_));
    InMux I__4144 (
            .O(N__26525),
            .I(N__26521));
    InMux I__4143 (
            .O(N__26524),
            .I(N__26518));
    LocalMux I__4142 (
            .O(N__26521),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    LocalMux I__4141 (
            .O(N__26518),
            .I(\dron_frame_decoder_1.WDTZ0Z_9 ));
    InMux I__4140 (
            .O(N__26513),
            .I(\dron_frame_decoder_1.un1_WDT_cry_8 ));
    InMux I__4139 (
            .O(N__26510),
            .I(N__26506));
    InMux I__4138 (
            .O(N__26509),
            .I(N__26503));
    LocalMux I__4137 (
            .O(N__26506),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    LocalMux I__4136 (
            .O(N__26503),
            .I(\dron_frame_decoder_1.WDTZ0Z_10 ));
    InMux I__4135 (
            .O(N__26498),
            .I(\dron_frame_decoder_1.un1_WDT_cry_9 ));
    InMux I__4134 (
            .O(N__26495),
            .I(N__26490));
    InMux I__4133 (
            .O(N__26494),
            .I(N__26485));
    InMux I__4132 (
            .O(N__26493),
            .I(N__26485));
    LocalMux I__4131 (
            .O(N__26490),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    LocalMux I__4130 (
            .O(N__26485),
            .I(\dron_frame_decoder_1.WDTZ0Z_11 ));
    InMux I__4129 (
            .O(N__26480),
            .I(\dron_frame_decoder_1.un1_WDT_cry_10 ));
    InMux I__4128 (
            .O(N__26477),
            .I(N__26474));
    LocalMux I__4127 (
            .O(N__26474),
            .I(N__26471));
    Odrv4 I__4126 (
            .O(N__26471),
            .I(\scaler_4.N_1684_i_l_ofxZ0 ));
    InMux I__4125 (
            .O(N__26468),
            .I(bfn_8_10_0_));
    InMux I__4124 (
            .O(N__26465),
            .I(\scaler_4.un3_source_data_0_cry_8 ));
    SRMux I__4123 (
            .O(N__26462),
            .I(N__26459));
    LocalMux I__4122 (
            .O(N__26459),
            .I(N__26455));
    SRMux I__4121 (
            .O(N__26458),
            .I(N__26452));
    Span4Mux_v I__4120 (
            .O(N__26455),
            .I(N__26449));
    LocalMux I__4119 (
            .O(N__26452),
            .I(N__26446));
    Span4Mux_h I__4118 (
            .O(N__26449),
            .I(N__26441));
    Span4Mux_h I__4117 (
            .O(N__26446),
            .I(N__26441));
    Odrv4 I__4116 (
            .O(N__26441),
            .I(\Commands_frame_decoder.un1_state57_iZ0 ));
    CascadeMux I__4115 (
            .O(N__26438),
            .I(N__26434));
    InMux I__4114 (
            .O(N__26437),
            .I(N__26431));
    InMux I__4113 (
            .O(N__26434),
            .I(N__26428));
    LocalMux I__4112 (
            .O(N__26431),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    LocalMux I__4111 (
            .O(N__26428),
            .I(\dron_frame_decoder_1.WDT10_0_i ));
    InMux I__4110 (
            .O(N__26423),
            .I(N__26420));
    LocalMux I__4109 (
            .O(N__26420),
            .I(\dron_frame_decoder_1.WDTZ0Z_0 ));
    InMux I__4108 (
            .O(N__26417),
            .I(N__26414));
    LocalMux I__4107 (
            .O(N__26414),
            .I(\dron_frame_decoder_1.WDTZ0Z_1 ));
    InMux I__4106 (
            .O(N__26411),
            .I(\dron_frame_decoder_1.un1_WDT_cry_0 ));
    InMux I__4105 (
            .O(N__26408),
            .I(N__26405));
    LocalMux I__4104 (
            .O(N__26405),
            .I(\dron_frame_decoder_1.WDTZ0Z_2 ));
    InMux I__4103 (
            .O(N__26402),
            .I(\dron_frame_decoder_1.un1_WDT_cry_1 ));
    InMux I__4102 (
            .O(N__26399),
            .I(N__26396));
    LocalMux I__4101 (
            .O(N__26396),
            .I(frame_decoder_CH4data_1));
    CascadeMux I__4100 (
            .O(N__26393),
            .I(N__26390));
    InMux I__4099 (
            .O(N__26390),
            .I(N__26387));
    LocalMux I__4098 (
            .O(N__26387),
            .I(frame_decoder_OFF4data_1));
    InMux I__4097 (
            .O(N__26384),
            .I(\scaler_4.un3_source_data_0_cry_0 ));
    InMux I__4096 (
            .O(N__26381),
            .I(N__26378));
    LocalMux I__4095 (
            .O(N__26378),
            .I(frame_decoder_CH4data_2));
    CascadeMux I__4094 (
            .O(N__26375),
            .I(N__26372));
    InMux I__4093 (
            .O(N__26372),
            .I(N__26369));
    LocalMux I__4092 (
            .O(N__26369),
            .I(frame_decoder_OFF4data_2));
    InMux I__4091 (
            .O(N__26366),
            .I(\scaler_4.un3_source_data_0_cry_1 ));
    InMux I__4090 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__4089 (
            .O(N__26360),
            .I(frame_decoder_CH4data_3));
    CascadeMux I__4088 (
            .O(N__26357),
            .I(N__26354));
    InMux I__4087 (
            .O(N__26354),
            .I(N__26351));
    LocalMux I__4086 (
            .O(N__26351),
            .I(frame_decoder_OFF4data_3));
    InMux I__4085 (
            .O(N__26348),
            .I(\scaler_4.un3_source_data_0_cry_2 ));
    InMux I__4084 (
            .O(N__26345),
            .I(N__26342));
    LocalMux I__4083 (
            .O(N__26342),
            .I(frame_decoder_CH4data_4));
    CascadeMux I__4082 (
            .O(N__26339),
            .I(N__26336));
    InMux I__4081 (
            .O(N__26336),
            .I(N__26333));
    LocalMux I__4080 (
            .O(N__26333),
            .I(frame_decoder_OFF4data_4));
    InMux I__4079 (
            .O(N__26330),
            .I(\scaler_4.un3_source_data_0_cry_3 ));
    InMux I__4078 (
            .O(N__26327),
            .I(N__26324));
    LocalMux I__4077 (
            .O(N__26324),
            .I(N__26321));
    Span4Mux_h I__4076 (
            .O(N__26321),
            .I(N__26318));
    Odrv4 I__4075 (
            .O(N__26318),
            .I(frame_decoder_CH4data_5));
    CascadeMux I__4074 (
            .O(N__26315),
            .I(N__26312));
    InMux I__4073 (
            .O(N__26312),
            .I(N__26309));
    LocalMux I__4072 (
            .O(N__26309),
            .I(frame_decoder_OFF4data_5));
    InMux I__4071 (
            .O(N__26306),
            .I(\scaler_4.un3_source_data_0_cry_4 ));
    InMux I__4070 (
            .O(N__26303),
            .I(N__26300));
    LocalMux I__4069 (
            .O(N__26300),
            .I(frame_decoder_CH4data_6));
    CascadeMux I__4068 (
            .O(N__26297),
            .I(N__26294));
    InMux I__4067 (
            .O(N__26294),
            .I(N__26291));
    LocalMux I__4066 (
            .O(N__26291),
            .I(N__26288));
    Span4Mux_h I__4065 (
            .O(N__26288),
            .I(N__26285));
    Span4Mux_h I__4064 (
            .O(N__26285),
            .I(N__26282));
    Odrv4 I__4063 (
            .O(N__26282),
            .I(frame_decoder_OFF4data_6));
    InMux I__4062 (
            .O(N__26279),
            .I(\scaler_4.un3_source_data_0_cry_5 ));
    InMux I__4061 (
            .O(N__26276),
            .I(N__26273));
    LocalMux I__4060 (
            .O(N__26273),
            .I(N__26270));
    Span12Mux_s9_v I__4059 (
            .O(N__26270),
            .I(N__26267));
    Odrv12 I__4058 (
            .O(N__26267),
            .I(\scaler_4.un3_source_data_0_axb_7 ));
    InMux I__4057 (
            .O(N__26264),
            .I(\scaler_4.un3_source_data_0_cry_6 ));
    InMux I__4056 (
            .O(N__26261),
            .I(N__26257));
    InMux I__4055 (
            .O(N__26260),
            .I(N__26254));
    LocalMux I__4054 (
            .O(N__26257),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    LocalMux I__4053 (
            .O(N__26254),
            .I(\Commands_frame_decoder.WDTZ0Z_7 ));
    InMux I__4052 (
            .O(N__26249),
            .I(\Commands_frame_decoder.un1_WDT_cry_6 ));
    InMux I__4051 (
            .O(N__26246),
            .I(N__26242));
    InMux I__4050 (
            .O(N__26245),
            .I(N__26239));
    LocalMux I__4049 (
            .O(N__26242),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    LocalMux I__4048 (
            .O(N__26239),
            .I(\Commands_frame_decoder.WDTZ0Z_8 ));
    InMux I__4047 (
            .O(N__26234),
            .I(bfn_8_8_0_));
    CascadeMux I__4046 (
            .O(N__26231),
            .I(N__26227));
    InMux I__4045 (
            .O(N__26230),
            .I(N__26224));
    InMux I__4044 (
            .O(N__26227),
            .I(N__26221));
    LocalMux I__4043 (
            .O(N__26224),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    LocalMux I__4042 (
            .O(N__26221),
            .I(\Commands_frame_decoder.WDTZ0Z_9 ));
    InMux I__4041 (
            .O(N__26216),
            .I(\Commands_frame_decoder.un1_WDT_cry_8 ));
    InMux I__4040 (
            .O(N__26213),
            .I(N__26209));
    InMux I__4039 (
            .O(N__26212),
            .I(N__26206));
    LocalMux I__4038 (
            .O(N__26209),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    LocalMux I__4037 (
            .O(N__26206),
            .I(\Commands_frame_decoder.WDTZ0Z_10 ));
    InMux I__4036 (
            .O(N__26201),
            .I(\Commands_frame_decoder.un1_WDT_cry_9 ));
    InMux I__4035 (
            .O(N__26198),
            .I(N__26193));
    InMux I__4034 (
            .O(N__26197),
            .I(N__26188));
    InMux I__4033 (
            .O(N__26196),
            .I(N__26188));
    LocalMux I__4032 (
            .O(N__26193),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    LocalMux I__4031 (
            .O(N__26188),
            .I(\Commands_frame_decoder.WDTZ0Z_11 ));
    InMux I__4030 (
            .O(N__26183),
            .I(\Commands_frame_decoder.un1_WDT_cry_10 ));
    InMux I__4029 (
            .O(N__26180),
            .I(N__26175));
    InMux I__4028 (
            .O(N__26179),
            .I(N__26170));
    InMux I__4027 (
            .O(N__26178),
            .I(N__26170));
    LocalMux I__4026 (
            .O(N__26175),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    LocalMux I__4025 (
            .O(N__26170),
            .I(\Commands_frame_decoder.WDTZ0Z_12 ));
    InMux I__4024 (
            .O(N__26165),
            .I(\Commands_frame_decoder.un1_WDT_cry_11 ));
    CascadeMux I__4023 (
            .O(N__26162),
            .I(N__26158));
    InMux I__4022 (
            .O(N__26161),
            .I(N__26155));
    InMux I__4021 (
            .O(N__26158),
            .I(N__26152));
    LocalMux I__4020 (
            .O(N__26155),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    LocalMux I__4019 (
            .O(N__26152),
            .I(\Commands_frame_decoder.WDTZ0Z_13 ));
    InMux I__4018 (
            .O(N__26147),
            .I(\Commands_frame_decoder.un1_WDT_cry_12 ));
    InMux I__4017 (
            .O(N__26144),
            .I(N__26138));
    InMux I__4016 (
            .O(N__26143),
            .I(N__26131));
    InMux I__4015 (
            .O(N__26142),
            .I(N__26131));
    InMux I__4014 (
            .O(N__26141),
            .I(N__26131));
    LocalMux I__4013 (
            .O(N__26138),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    LocalMux I__4012 (
            .O(N__26131),
            .I(\Commands_frame_decoder.WDTZ0Z_14 ));
    InMux I__4011 (
            .O(N__26126),
            .I(\Commands_frame_decoder.un1_WDT_cry_13 ));
    InMux I__4010 (
            .O(N__26123),
            .I(\Commands_frame_decoder.un1_WDT_cry_14 ));
    CascadeMux I__4009 (
            .O(N__26120),
            .I(N__26117));
    InMux I__4008 (
            .O(N__26117),
            .I(N__26109));
    InMux I__4007 (
            .O(N__26116),
            .I(N__26109));
    InMux I__4006 (
            .O(N__26115),
            .I(N__26106));
    InMux I__4005 (
            .O(N__26114),
            .I(N__26103));
    LocalMux I__4004 (
            .O(N__26109),
            .I(N__26100));
    LocalMux I__4003 (
            .O(N__26106),
            .I(N__26097));
    LocalMux I__4002 (
            .O(N__26103),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__4001 (
            .O(N__26100),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    Odrv4 I__4000 (
            .O(N__26097),
            .I(\Commands_frame_decoder.WDTZ0Z_15 ));
    InMux I__3999 (
            .O(N__26090),
            .I(N__26087));
    LocalMux I__3998 (
            .O(N__26087),
            .I(\Commands_frame_decoder.count_1_sqmuxa ));
    CascadeMux I__3997 (
            .O(N__26084),
            .I(N__26080));
    InMux I__3996 (
            .O(N__26083),
            .I(N__26077));
    InMux I__3995 (
            .O(N__26080),
            .I(N__26074));
    LocalMux I__3994 (
            .O(N__26077),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    LocalMux I__3993 (
            .O(N__26074),
            .I(\Commands_frame_decoder.state_0_sqmuxa ));
    InMux I__3992 (
            .O(N__26069),
            .I(N__26066));
    LocalMux I__3991 (
            .O(N__26066),
            .I(\Commands_frame_decoder.WDTZ0Z_0 ));
    InMux I__3990 (
            .O(N__26063),
            .I(N__26060));
    LocalMux I__3989 (
            .O(N__26060),
            .I(\Commands_frame_decoder.WDTZ0Z_1 ));
    InMux I__3988 (
            .O(N__26057),
            .I(\Commands_frame_decoder.un1_WDT_cry_0 ));
    InMux I__3987 (
            .O(N__26054),
            .I(N__26051));
    LocalMux I__3986 (
            .O(N__26051),
            .I(\Commands_frame_decoder.WDTZ0Z_2 ));
    InMux I__3985 (
            .O(N__26048),
            .I(\Commands_frame_decoder.un1_WDT_cry_1 ));
    InMux I__3984 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__3983 (
            .O(N__26042),
            .I(\Commands_frame_decoder.WDTZ0Z_3 ));
    InMux I__3982 (
            .O(N__26039),
            .I(\Commands_frame_decoder.un1_WDT_cry_2 ));
    InMux I__3981 (
            .O(N__26036),
            .I(N__26032));
    InMux I__3980 (
            .O(N__26035),
            .I(N__26029));
    LocalMux I__3979 (
            .O(N__26032),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    LocalMux I__3978 (
            .O(N__26029),
            .I(\Commands_frame_decoder.WDTZ0Z_4 ));
    InMux I__3977 (
            .O(N__26024),
            .I(\Commands_frame_decoder.un1_WDT_cry_3 ));
    InMux I__3976 (
            .O(N__26021),
            .I(N__26017));
    InMux I__3975 (
            .O(N__26020),
            .I(N__26014));
    LocalMux I__3974 (
            .O(N__26017),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    LocalMux I__3973 (
            .O(N__26014),
            .I(\Commands_frame_decoder.WDTZ0Z_5 ));
    InMux I__3972 (
            .O(N__26009),
            .I(\Commands_frame_decoder.un1_WDT_cry_4 ));
    InMux I__3971 (
            .O(N__26006),
            .I(N__26002));
    InMux I__3970 (
            .O(N__26005),
            .I(N__25999));
    LocalMux I__3969 (
            .O(N__26002),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    LocalMux I__3968 (
            .O(N__25999),
            .I(\Commands_frame_decoder.WDTZ0Z_6 ));
    InMux I__3967 (
            .O(N__25994),
            .I(\Commands_frame_decoder.un1_WDT_cry_5 ));
    InMux I__3966 (
            .O(N__25991),
            .I(N__25988));
    LocalMux I__3965 (
            .O(N__25988),
            .I(N__25985));
    Odrv4 I__3964 (
            .O(N__25985),
            .I(\pid_side.error_axbZ0Z_2 ));
    InMux I__3963 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__3962 (
            .O(N__25979),
            .I(N__25976));
    Odrv4 I__3961 (
            .O(N__25976),
            .I(\pid_side.error_axbZ0Z_3 ));
    InMux I__3960 (
            .O(N__25973),
            .I(N__25970));
    LocalMux I__3959 (
            .O(N__25970),
            .I(N__25967));
    Span4Mux_s3_h I__3958 (
            .O(N__25967),
            .I(N__25963));
    InMux I__3957 (
            .O(N__25966),
            .I(N__25960));
    Span4Mux_h I__3956 (
            .O(N__25963),
            .I(N__25957));
    LocalMux I__3955 (
            .O(N__25960),
            .I(alt_kp_4));
    Odrv4 I__3954 (
            .O(N__25957),
            .I(alt_kp_4));
    CEMux I__3953 (
            .O(N__25952),
            .I(N__25949));
    LocalMux I__3952 (
            .O(N__25949),
            .I(N__25944));
    CEMux I__3951 (
            .O(N__25948),
            .I(N__25941));
    CEMux I__3950 (
            .O(N__25947),
            .I(N__25938));
    Span4Mux_s3_h I__3949 (
            .O(N__25944),
            .I(N__25933));
    LocalMux I__3948 (
            .O(N__25941),
            .I(N__25933));
    LocalMux I__3947 (
            .O(N__25938),
            .I(N__25930));
    Span4Mux_h I__3946 (
            .O(N__25933),
            .I(N__25925));
    Span4Mux_h I__3945 (
            .O(N__25930),
            .I(N__25925));
    Odrv4 I__3944 (
            .O(N__25925),
            .I(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ));
    InMux I__3943 (
            .O(N__25922),
            .I(N__25919));
    LocalMux I__3942 (
            .O(N__25919),
            .I(N__25916));
    Span12Mux_s8_v I__3941 (
            .O(N__25916),
            .I(N__25913));
    Odrv12 I__3940 (
            .O(N__25913),
            .I(\pid_alt.state_RNIFCSD1Z0Z_0 ));
    IoInMux I__3939 (
            .O(N__25910),
            .I(N__25907));
    LocalMux I__3938 (
            .O(N__25907),
            .I(N__25904));
    Span4Mux_s1_v I__3937 (
            .O(N__25904),
            .I(N__25901));
    Odrv4 I__3936 (
            .O(N__25901),
            .I(\pid_alt.N_850_0 ));
    InMux I__3935 (
            .O(N__25898),
            .I(N__25895));
    LocalMux I__3934 (
            .O(N__25895),
            .I(uart_input_drone_c));
    InMux I__3933 (
            .O(N__25892),
            .I(N__25889));
    LocalMux I__3932 (
            .O(N__25889),
            .I(\uart_drone_sync.aux_0__0__0_0 ));
    InMux I__3931 (
            .O(N__25886),
            .I(N__25883));
    LocalMux I__3930 (
            .O(N__25883),
            .I(\uart_drone_sync.aux_1__0__0_0 ));
    CEMux I__3929 (
            .O(N__25880),
            .I(N__25877));
    LocalMux I__3928 (
            .O(N__25877),
            .I(N__25874));
    Span4Mux_v I__3927 (
            .O(N__25874),
            .I(N__25871));
    Span4Mux_h I__3926 (
            .O(N__25871),
            .I(N__25868));
    Odrv4 I__3925 (
            .O(N__25868),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ));
    InMux I__3924 (
            .O(N__25865),
            .I(N__25862));
    LocalMux I__3923 (
            .O(N__25862),
            .I(N__25859));
    Span4Mux_h I__3922 (
            .O(N__25859),
            .I(N__25856));
    Odrv4 I__3921 (
            .O(N__25856),
            .I(\pid_alt.pid_preregZ0Z_14 ));
    InMux I__3920 (
            .O(N__25853),
            .I(N__25850));
    LocalMux I__3919 (
            .O(N__25850),
            .I(N__25847));
    Odrv4 I__3918 (
            .O(N__25847),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ));
    CascadeMux I__3917 (
            .O(N__25844),
            .I(N__25841));
    InMux I__3916 (
            .O(N__25841),
            .I(N__25838));
    LocalMux I__3915 (
            .O(N__25838),
            .I(N__25835));
    Odrv4 I__3914 (
            .O(N__25835),
            .I(\pid_alt.pid_preregZ0Z_16 ));
    InMux I__3913 (
            .O(N__25832),
            .I(N__25829));
    LocalMux I__3912 (
            .O(N__25829),
            .I(N__25826));
    Odrv4 I__3911 (
            .O(N__25826),
            .I(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5 ));
    CEMux I__3910 (
            .O(N__25823),
            .I(N__25820));
    LocalMux I__3909 (
            .O(N__25820),
            .I(N__25816));
    CEMux I__3908 (
            .O(N__25819),
            .I(N__25813));
    Span4Mux_s3_h I__3907 (
            .O(N__25816),
            .I(N__25810));
    LocalMux I__3906 (
            .O(N__25813),
            .I(N__25807));
    Span4Mux_h I__3905 (
            .O(N__25810),
            .I(N__25804));
    Span4Mux_v I__3904 (
            .O(N__25807),
            .I(N__25801));
    Odrv4 I__3903 (
            .O(N__25804),
            .I(\dron_frame_decoder_1.N_755_0 ));
    Odrv4 I__3902 (
            .O(N__25801),
            .I(\dron_frame_decoder_1.N_755_0 ));
    InMux I__3901 (
            .O(N__25796),
            .I(N__25793));
    LocalMux I__3900 (
            .O(N__25793),
            .I(N__25790));
    Odrv12 I__3899 (
            .O(N__25790),
            .I(\dron_frame_decoder_1.drone_altitude_7 ));
    InMux I__3898 (
            .O(N__25787),
            .I(N__25783));
    InMux I__3897 (
            .O(N__25786),
            .I(N__25780));
    LocalMux I__3896 (
            .O(N__25783),
            .I(N__25777));
    LocalMux I__3895 (
            .O(N__25780),
            .I(N__25774));
    Span4Mux_v I__3894 (
            .O(N__25777),
            .I(N__25771));
    Odrv4 I__3893 (
            .O(N__25774),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    Odrv4 I__3892 (
            .O(N__25771),
            .I(\Commands_frame_decoder.source_CH2data_1_sqmuxa ));
    CascadeMux I__3891 (
            .O(N__25766),
            .I(N__25763));
    InMux I__3890 (
            .O(N__25763),
            .I(N__25760));
    LocalMux I__3889 (
            .O(N__25760),
            .I(N__25757));
    Odrv4 I__3888 (
            .O(N__25757),
            .I(drone_H_disp_side_i_4));
    CascadeMux I__3887 (
            .O(N__25754),
            .I(N__25751));
    InMux I__3886 (
            .O(N__25751),
            .I(N__25748));
    LocalMux I__3885 (
            .O(N__25748),
            .I(N__25745));
    Odrv4 I__3884 (
            .O(N__25745),
            .I(drone_H_disp_side_i_7));
    CascadeMux I__3883 (
            .O(N__25742),
            .I(N__25739));
    InMux I__3882 (
            .O(N__25739),
            .I(N__25736));
    LocalMux I__3881 (
            .O(N__25736),
            .I(N__25733));
    Odrv4 I__3880 (
            .O(N__25733),
            .I(drone_H_disp_side_i_5));
    InMux I__3879 (
            .O(N__25730),
            .I(N__25727));
    LocalMux I__3878 (
            .O(N__25727),
            .I(N__25724));
    Odrv4 I__3877 (
            .O(N__25724),
            .I(\pid_alt.m7_e_4 ));
    InMux I__3876 (
            .O(N__25721),
            .I(N__25718));
    LocalMux I__3875 (
            .O(N__25718),
            .I(N__25715));
    Span4Mux_h I__3874 (
            .O(N__25715),
            .I(N__25710));
    InMux I__3873 (
            .O(N__25714),
            .I(N__25705));
    InMux I__3872 (
            .O(N__25713),
            .I(N__25705));
    Odrv4 I__3871 (
            .O(N__25710),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    LocalMux I__3870 (
            .O(N__25705),
            .I(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ));
    CascadeMux I__3869 (
            .O(N__25700),
            .I(N__25697));
    InMux I__3868 (
            .O(N__25697),
            .I(N__25694));
    LocalMux I__3867 (
            .O(N__25694),
            .I(\pid_alt.error_i_acumm_preregZ0Z_19 ));
    CascadeMux I__3866 (
            .O(N__25691),
            .I(\pid_alt.un1_reset_i_a5_1_10_7_cascade_ ));
    InMux I__3865 (
            .O(N__25688),
            .I(N__25685));
    LocalMux I__3864 (
            .O(N__25685),
            .I(N__25680));
    InMux I__3863 (
            .O(N__25684),
            .I(N__25675));
    InMux I__3862 (
            .O(N__25683),
            .I(N__25675));
    Odrv12 I__3861 (
            .O(N__25680),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    LocalMux I__3860 (
            .O(N__25675),
            .I(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ));
    InMux I__3859 (
            .O(N__25670),
            .I(N__25667));
    LocalMux I__3858 (
            .O(N__25667),
            .I(\pid_alt.error_i_acumm_preregZ0Z_18 ));
    InMux I__3857 (
            .O(N__25664),
            .I(N__25661));
    LocalMux I__3856 (
            .O(N__25661),
            .I(N__25656));
    InMux I__3855 (
            .O(N__25660),
            .I(N__25651));
    InMux I__3854 (
            .O(N__25659),
            .I(N__25651));
    Odrv12 I__3853 (
            .O(N__25656),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    LocalMux I__3852 (
            .O(N__25651),
            .I(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ));
    InMux I__3851 (
            .O(N__25646),
            .I(N__25643));
    LocalMux I__3850 (
            .O(N__25643),
            .I(\pid_alt.error_i_acumm_preregZ0Z_17 ));
    InMux I__3849 (
            .O(N__25640),
            .I(N__25637));
    LocalMux I__3848 (
            .O(N__25637),
            .I(N__25632));
    InMux I__3847 (
            .O(N__25636),
            .I(N__25627));
    InMux I__3846 (
            .O(N__25635),
            .I(N__25627));
    Span4Mux_v I__3845 (
            .O(N__25632),
            .I(N__25622));
    LocalMux I__3844 (
            .O(N__25627),
            .I(N__25622));
    Span4Mux_h I__3843 (
            .O(N__25622),
            .I(N__25619));
    Odrv4 I__3842 (
            .O(N__25619),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ));
    CascadeMux I__3841 (
            .O(N__25616),
            .I(N__25613));
    InMux I__3840 (
            .O(N__25613),
            .I(N__25610));
    LocalMux I__3839 (
            .O(N__25610),
            .I(N__25607));
    Span4Mux_h I__3838 (
            .O(N__25607),
            .I(N__25604));
    Odrv4 I__3837 (
            .O(N__25604),
            .I(\pid_alt.error_i_acumm_preregZ0Z_20 ));
    InMux I__3836 (
            .O(N__25601),
            .I(N__25598));
    LocalMux I__3835 (
            .O(N__25598),
            .I(N__25593));
    InMux I__3834 (
            .O(N__25597),
            .I(N__25588));
    InMux I__3833 (
            .O(N__25596),
            .I(N__25588));
    Odrv12 I__3832 (
            .O(N__25593),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    LocalMux I__3831 (
            .O(N__25588),
            .I(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ));
    InMux I__3830 (
            .O(N__25583),
            .I(N__25580));
    LocalMux I__3829 (
            .O(N__25580),
            .I(\pid_alt.error_i_acumm_preregZ0Z_16 ));
    CEMux I__3828 (
            .O(N__25577),
            .I(N__25505));
    CEMux I__3827 (
            .O(N__25576),
            .I(N__25505));
    CEMux I__3826 (
            .O(N__25575),
            .I(N__25505));
    CEMux I__3825 (
            .O(N__25574),
            .I(N__25505));
    CEMux I__3824 (
            .O(N__25573),
            .I(N__25505));
    CEMux I__3823 (
            .O(N__25572),
            .I(N__25505));
    CEMux I__3822 (
            .O(N__25571),
            .I(N__25505));
    CEMux I__3821 (
            .O(N__25570),
            .I(N__25505));
    CEMux I__3820 (
            .O(N__25569),
            .I(N__25505));
    CEMux I__3819 (
            .O(N__25568),
            .I(N__25505));
    CEMux I__3818 (
            .O(N__25567),
            .I(N__25505));
    CEMux I__3817 (
            .O(N__25566),
            .I(N__25505));
    CEMux I__3816 (
            .O(N__25565),
            .I(N__25505));
    CEMux I__3815 (
            .O(N__25564),
            .I(N__25505));
    CEMux I__3814 (
            .O(N__25563),
            .I(N__25505));
    CEMux I__3813 (
            .O(N__25562),
            .I(N__25505));
    CEMux I__3812 (
            .O(N__25561),
            .I(N__25505));
    CEMux I__3811 (
            .O(N__25560),
            .I(N__25505));
    CEMux I__3810 (
            .O(N__25559),
            .I(N__25505));
    CEMux I__3809 (
            .O(N__25558),
            .I(N__25505));
    CEMux I__3808 (
            .O(N__25557),
            .I(N__25505));
    CEMux I__3807 (
            .O(N__25556),
            .I(N__25505));
    CEMux I__3806 (
            .O(N__25555),
            .I(N__25505));
    CEMux I__3805 (
            .O(N__25554),
            .I(N__25505));
    GlobalMux I__3804 (
            .O(N__25505),
            .I(N__25502));
    gio2CtrlBuf I__3803 (
            .O(N__25502),
            .I(\pid_alt.state_0_g_0 ));
    InMux I__3802 (
            .O(N__25499),
            .I(N__25487));
    InMux I__3801 (
            .O(N__25498),
            .I(N__25487));
    InMux I__3800 (
            .O(N__25497),
            .I(N__25487));
    InMux I__3799 (
            .O(N__25496),
            .I(N__25487));
    LocalMux I__3798 (
            .O(N__25487),
            .I(N__25483));
    InMux I__3797 (
            .O(N__25486),
            .I(N__25480));
    Span4Mux_v I__3796 (
            .O(N__25483),
            .I(N__25477));
    LocalMux I__3795 (
            .O(N__25480),
            .I(N__25474));
    Odrv4 I__3794 (
            .O(N__25477),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    Odrv4 I__3793 (
            .O(N__25474),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0 ));
    CascadeMux I__3792 (
            .O(N__25469),
            .I(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ));
    InMux I__3791 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__3790 (
            .O(N__25463),
            .I(\dron_frame_decoder_1.WDT10lto13_1 ));
    CascadeMux I__3789 (
            .O(N__25460),
            .I(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ));
    InMux I__3788 (
            .O(N__25457),
            .I(N__25454));
    LocalMux I__3787 (
            .O(N__25454),
            .I(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ));
    InMux I__3786 (
            .O(N__25451),
            .I(N__25447));
    InMux I__3785 (
            .O(N__25450),
            .I(N__25444));
    LocalMux I__3784 (
            .O(N__25447),
            .I(N__25441));
    LocalMux I__3783 (
            .O(N__25444),
            .I(N__25438));
    Odrv12 I__3782 (
            .O(N__25441),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    Odrv4 I__3781 (
            .O(N__25438),
            .I(\Commands_frame_decoder.source_CH3data_1_sqmuxa ));
    InMux I__3780 (
            .O(N__25433),
            .I(N__25430));
    LocalMux I__3779 (
            .O(N__25430),
            .I(N__25426));
    CascadeMux I__3778 (
            .O(N__25429),
            .I(N__25423));
    Span4Mux_h I__3777 (
            .O(N__25426),
            .I(N__25420));
    InMux I__3776 (
            .O(N__25423),
            .I(N__25417));
    Span4Mux_v I__3775 (
            .O(N__25420),
            .I(N__25414));
    LocalMux I__3774 (
            .O(N__25417),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    Odrv4 I__3773 (
            .O(N__25414),
            .I(\Commands_frame_decoder.stateZ0Z_2 ));
    CascadeMux I__3772 (
            .O(N__25409),
            .I(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ));
    InMux I__3771 (
            .O(N__25406),
            .I(N__25402));
    InMux I__3770 (
            .O(N__25405),
            .I(N__25399));
    LocalMux I__3769 (
            .O(N__25402),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    LocalMux I__3768 (
            .O(N__25399),
            .I(\Commands_frame_decoder.stateZ0Z_3 ));
    InMux I__3767 (
            .O(N__25394),
            .I(N__25390));
    InMux I__3766 (
            .O(N__25393),
            .I(N__25387));
    LocalMux I__3765 (
            .O(N__25390),
            .I(N__25382));
    LocalMux I__3764 (
            .O(N__25387),
            .I(N__25382));
    Odrv12 I__3763 (
            .O(N__25382),
            .I(frame_decoder_OFF4data_7));
    InMux I__3762 (
            .O(N__25379),
            .I(N__25376));
    LocalMux I__3761 (
            .O(N__25376),
            .I(N__25373));
    Odrv4 I__3760 (
            .O(N__25373),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa ));
    InMux I__3759 (
            .O(N__25370),
            .I(N__25364));
    InMux I__3758 (
            .O(N__25369),
            .I(N__25364));
    LocalMux I__3757 (
            .O(N__25364),
            .I(\Commands_frame_decoder.stateZ0Z_4 ));
    InMux I__3756 (
            .O(N__25361),
            .I(N__25355));
    InMux I__3755 (
            .O(N__25360),
            .I(N__25355));
    LocalMux I__3754 (
            .O(N__25355),
            .I(\Commands_frame_decoder.WDT8lt14_0 ));
    InMux I__3753 (
            .O(N__25352),
            .I(N__25349));
    LocalMux I__3752 (
            .O(N__25349),
            .I(N__25346));
    Odrv4 I__3751 (
            .O(N__25346),
            .I(\Commands_frame_decoder.N_377_0 ));
    CascadeMux I__3750 (
            .O(N__25343),
            .I(\Commands_frame_decoder.N_377_0_cascade_ ));
    InMux I__3749 (
            .O(N__25340),
            .I(N__25337));
    LocalMux I__3748 (
            .O(N__25337),
            .I(N__25333));
    InMux I__3747 (
            .O(N__25336),
            .I(N__25330));
    Odrv4 I__3746 (
            .O(N__25333),
            .I(\Commands_frame_decoder.N_384 ));
    LocalMux I__3745 (
            .O(N__25330),
            .I(\Commands_frame_decoder.N_384 ));
    CEMux I__3744 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__3743 (
            .O(N__25322),
            .I(N__25319));
    Span4Mux_v I__3742 (
            .O(N__25319),
            .I(N__25315));
    CEMux I__3741 (
            .O(N__25318),
            .I(N__25312));
    Odrv4 I__3740 (
            .O(N__25315),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    LocalMux I__3739 (
            .O(N__25312),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ));
    CascadeMux I__3738 (
            .O(N__25307),
            .I(N__25303));
    CascadeMux I__3737 (
            .O(N__25306),
            .I(N__25300));
    InMux I__3736 (
            .O(N__25303),
            .I(N__25297));
    InMux I__3735 (
            .O(N__25300),
            .I(N__25294));
    LocalMux I__3734 (
            .O(N__25297),
            .I(N__25291));
    LocalMux I__3733 (
            .O(N__25294),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    Odrv4 I__3732 (
            .O(N__25291),
            .I(\Commands_frame_decoder.stateZ0Z_12 ));
    InMux I__3731 (
            .O(N__25286),
            .I(N__25280));
    InMux I__3730 (
            .O(N__25285),
            .I(N__25280));
    LocalMux I__3729 (
            .O(N__25280),
            .I(\Commands_frame_decoder.stateZ0Z_13 ));
    InMux I__3728 (
            .O(N__25277),
            .I(N__25274));
    LocalMux I__3727 (
            .O(N__25274),
            .I(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ));
    CascadeMux I__3726 (
            .O(N__25271),
            .I(\Commands_frame_decoder.WDT8lto13_1_cascade_ ));
    InMux I__3725 (
            .O(N__25268),
            .I(N__25265));
    LocalMux I__3724 (
            .O(N__25265),
            .I(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ));
    InMux I__3723 (
            .O(N__25262),
            .I(N__25258));
    InMux I__3722 (
            .O(N__25261),
            .I(N__25255));
    LocalMux I__3721 (
            .O(N__25258),
            .I(N__25252));
    LocalMux I__3720 (
            .O(N__25255),
            .I(N__25248));
    Span4Mux_h I__3719 (
            .O(N__25252),
            .I(N__25245));
    InMux I__3718 (
            .O(N__25251),
            .I(N__25242));
    Span4Mux_h I__3717 (
            .O(N__25248),
            .I(N__25239));
    Odrv4 I__3716 (
            .O(N__25245),
            .I(\Commands_frame_decoder.preinitZ0 ));
    LocalMux I__3715 (
            .O(N__25242),
            .I(\Commands_frame_decoder.preinitZ0 ));
    Odrv4 I__3714 (
            .O(N__25239),
            .I(\Commands_frame_decoder.preinitZ0 ));
    CascadeMux I__3713 (
            .O(N__25232),
            .I(\Commands_frame_decoder.WDT8lt14_0_cascade_ ));
    InMux I__3712 (
            .O(N__25229),
            .I(N__25226));
    LocalMux I__3711 (
            .O(N__25226),
            .I(drone_H_disp_side_i_6));
    InMux I__3710 (
            .O(N__25223),
            .I(N__25220));
    LocalMux I__3709 (
            .O(N__25220),
            .I(N__25217));
    Odrv4 I__3708 (
            .O(N__25217),
            .I(side_command_0));
    InMux I__3707 (
            .O(N__25214),
            .I(N__25211));
    LocalMux I__3706 (
            .O(N__25211),
            .I(side_command_1));
    CascadeMux I__3705 (
            .O(N__25208),
            .I(N__25205));
    InMux I__3704 (
            .O(N__25205),
            .I(N__25202));
    LocalMux I__3703 (
            .O(N__25202),
            .I(side_command_2));
    InMux I__3702 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3701 (
            .O(N__25196),
            .I(side_command_3));
    CascadeMux I__3700 (
            .O(N__25193),
            .I(N__25190));
    InMux I__3699 (
            .O(N__25190),
            .I(N__25187));
    LocalMux I__3698 (
            .O(N__25187),
            .I(side_command_4));
    CascadeMux I__3697 (
            .O(N__25184),
            .I(N__25181));
    InMux I__3696 (
            .O(N__25181),
            .I(N__25178));
    LocalMux I__3695 (
            .O(N__25178),
            .I(side_command_5));
    InMux I__3694 (
            .O(N__25175),
            .I(N__25172));
    LocalMux I__3693 (
            .O(N__25172),
            .I(side_command_6));
    InMux I__3692 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__3691 (
            .O(N__25166),
            .I(N__25163));
    Odrv4 I__3690 (
            .O(N__25163),
            .I(drone_H_disp_side_15));
    InMux I__3689 (
            .O(N__25160),
            .I(N__25157));
    LocalMux I__3688 (
            .O(N__25157),
            .I(N__25154));
    Odrv4 I__3687 (
            .O(N__25154),
            .I(\dron_frame_decoder_1.drone_altitude_5 ));
    InMux I__3686 (
            .O(N__25151),
            .I(N__25148));
    LocalMux I__3685 (
            .O(N__25148),
            .I(N__25145));
    Odrv4 I__3684 (
            .O(N__25145),
            .I(\dron_frame_decoder_1.drone_altitude_6 ));
    InMux I__3683 (
            .O(N__25142),
            .I(N__25138));
    InMux I__3682 (
            .O(N__25141),
            .I(N__25135));
    LocalMux I__3681 (
            .O(N__25138),
            .I(N__25132));
    LocalMux I__3680 (
            .O(N__25135),
            .I(N__25129));
    Span12Mux_s10_v I__3679 (
            .O(N__25132),
            .I(N__25126));
    Span4Mux_s3_h I__3678 (
            .O(N__25129),
            .I(N__25123));
    Span12Mux_h I__3677 (
            .O(N__25126),
            .I(N__25120));
    Span4Mux_v I__3676 (
            .O(N__25123),
            .I(N__25117));
    Odrv12 I__3675 (
            .O(N__25120),
            .I(xy_kp_0));
    Odrv4 I__3674 (
            .O(N__25117),
            .I(xy_kp_0));
    InMux I__3673 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__3672 (
            .O(N__25109),
            .I(N__25106));
    Span4Mux_s1_h I__3671 (
            .O(N__25106),
            .I(N__25102));
    InMux I__3670 (
            .O(N__25105),
            .I(N__25099));
    Span4Mux_v I__3669 (
            .O(N__25102),
            .I(N__25096));
    LocalMux I__3668 (
            .O(N__25099),
            .I(N__25093));
    Sp12to4 I__3667 (
            .O(N__25096),
            .I(N__25090));
    Span4Mux_s2_h I__3666 (
            .O(N__25093),
            .I(N__25087));
    Span12Mux_h I__3665 (
            .O(N__25090),
            .I(N__25084));
    Span4Mux_h I__3664 (
            .O(N__25087),
            .I(N__25081));
    Odrv12 I__3663 (
            .O(N__25084),
            .I(xy_kp_2));
    Odrv4 I__3662 (
            .O(N__25081),
            .I(xy_kp_2));
    InMux I__3661 (
            .O(N__25076),
            .I(N__25073));
    LocalMux I__3660 (
            .O(N__25073),
            .I(N__25070));
    Span4Mux_s3_h I__3659 (
            .O(N__25070),
            .I(N__25066));
    InMux I__3658 (
            .O(N__25069),
            .I(N__25063));
    Span4Mux_h I__3657 (
            .O(N__25066),
            .I(N__25060));
    LocalMux I__3656 (
            .O(N__25063),
            .I(N__25057));
    Span4Mux_v I__3655 (
            .O(N__25060),
            .I(N__25054));
    Span4Mux_s2_h I__3654 (
            .O(N__25057),
            .I(N__25051));
    Sp12to4 I__3653 (
            .O(N__25054),
            .I(N__25048));
    Span4Mux_v I__3652 (
            .O(N__25051),
            .I(N__25045));
    Odrv12 I__3651 (
            .O(N__25048),
            .I(xy_kp_6));
    Odrv4 I__3650 (
            .O(N__25045),
            .I(xy_kp_6));
    InMux I__3649 (
            .O(N__25040),
            .I(N__25037));
    LocalMux I__3648 (
            .O(N__25037),
            .I(\dron_frame_decoder_1.drone_altitude_4 ));
    InMux I__3647 (
            .O(N__25034),
            .I(N__25031));
    LocalMux I__3646 (
            .O(N__25031),
            .I(N__25028));
    Span4Mux_h I__3645 (
            .O(N__25028),
            .I(N__25025));
    Odrv4 I__3644 (
            .O(N__25025),
            .I(drone_altitude_i_4));
    InMux I__3643 (
            .O(N__25022),
            .I(N__25019));
    LocalMux I__3642 (
            .O(N__25019),
            .I(N__25016));
    Span4Mux_v I__3641 (
            .O(N__25016),
            .I(N__25012));
    CascadeMux I__3640 (
            .O(N__25015),
            .I(N__25009));
    Span4Mux_v I__3639 (
            .O(N__25012),
            .I(N__25006));
    InMux I__3638 (
            .O(N__25009),
            .I(N__25003));
    Odrv4 I__3637 (
            .O(N__25006),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    LocalMux I__3636 (
            .O(N__25003),
            .I(\pid_alt.error_i_regZ0Z_0 ));
    InMux I__3635 (
            .O(N__24998),
            .I(N__24995));
    LocalMux I__3634 (
            .O(N__24995),
            .I(N__24992));
    Span4Mux_v I__3633 (
            .O(N__24992),
            .I(N__24989));
    Span4Mux_v I__3632 (
            .O(N__24989),
            .I(N__24985));
    InMux I__3631 (
            .O(N__24988),
            .I(N__24982));
    Odrv4 I__3630 (
            .O(N__24985),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    LocalMux I__3629 (
            .O(N__24982),
            .I(\pid_alt.error_i_acummZ0Z_0 ));
    InMux I__3628 (
            .O(N__24977),
            .I(N__24974));
    LocalMux I__3627 (
            .O(N__24974),
            .I(N__24970));
    InMux I__3626 (
            .O(N__24973),
            .I(N__24967));
    Span4Mux_v I__3625 (
            .O(N__24970),
            .I(N__24964));
    LocalMux I__3624 (
            .O(N__24967),
            .I(N__24961));
    Odrv4 I__3623 (
            .O(N__24964),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    Odrv12 I__3622 (
            .O(N__24961),
            .I(\pid_alt.error_i_acumm_preregZ0Z_0 ));
    InMux I__3621 (
            .O(N__24956),
            .I(N__24953));
    LocalMux I__3620 (
            .O(N__24953),
            .I(drone_H_disp_side_i_13));
    InMux I__3619 (
            .O(N__24950),
            .I(N__24946));
    CascadeMux I__3618 (
            .O(N__24949),
            .I(N__24943));
    LocalMux I__3617 (
            .O(N__24946),
            .I(N__24940));
    InMux I__3616 (
            .O(N__24943),
            .I(N__24937));
    Span4Mux_v I__3615 (
            .O(N__24940),
            .I(N__24932));
    LocalMux I__3614 (
            .O(N__24937),
            .I(N__24932));
    Odrv4 I__3613 (
            .O(N__24932),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ));
    CascadeMux I__3612 (
            .O(N__24929),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ));
    InMux I__3611 (
            .O(N__24926),
            .I(N__24923));
    LocalMux I__3610 (
            .O(N__24923),
            .I(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ));
    InMux I__3609 (
            .O(N__24920),
            .I(N__24914));
    InMux I__3608 (
            .O(N__24919),
            .I(N__24914));
    LocalMux I__3607 (
            .O(N__24914),
            .I(N__24911));
    Span4Mux_v I__3606 (
            .O(N__24911),
            .I(N__24907));
    InMux I__3605 (
            .O(N__24910),
            .I(N__24904));
    Span4Mux_h I__3604 (
            .O(N__24907),
            .I(N__24899));
    LocalMux I__3603 (
            .O(N__24904),
            .I(N__24899));
    Span4Mux_v I__3602 (
            .O(N__24899),
            .I(N__24896));
    Span4Mux_v I__3601 (
            .O(N__24896),
            .I(N__24893));
    Odrv4 I__3600 (
            .O(N__24893),
            .I(\pid_alt.error_d_regZ0Z_19 ));
    InMux I__3599 (
            .O(N__24890),
            .I(N__24887));
    LocalMux I__3598 (
            .O(N__24887),
            .I(N__24883));
    InMux I__3597 (
            .O(N__24886),
            .I(N__24880));
    Span4Mux_h I__3596 (
            .O(N__24883),
            .I(N__24877));
    LocalMux I__3595 (
            .O(N__24880),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    Odrv4 I__3594 (
            .O(N__24877),
            .I(\pid_alt.error_d_reg_prevZ0Z_19 ));
    InMux I__3593 (
            .O(N__24872),
            .I(N__24866));
    InMux I__3592 (
            .O(N__24871),
            .I(N__24866));
    LocalMux I__3591 (
            .O(N__24866),
            .I(\pid_alt.error_d_reg_prevZ0Z_20 ));
    InMux I__3590 (
            .O(N__24863),
            .I(N__24857));
    InMux I__3589 (
            .O(N__24862),
            .I(N__24857));
    LocalMux I__3588 (
            .O(N__24857),
            .I(N__24854));
    Span4Mux_h I__3587 (
            .O(N__24854),
            .I(N__24851));
    Span4Mux_v I__3586 (
            .O(N__24851),
            .I(N__24848));
    Odrv4 I__3585 (
            .O(N__24848),
            .I(\pid_alt.error_p_regZ0Z_20 ));
    InMux I__3584 (
            .O(N__24845),
            .I(N__24840));
    InMux I__3583 (
            .O(N__24844),
            .I(N__24835));
    InMux I__3582 (
            .O(N__24843),
            .I(N__24835));
    LocalMux I__3581 (
            .O(N__24840),
            .I(N__24830));
    LocalMux I__3580 (
            .O(N__24835),
            .I(N__24830));
    Span12Mux_v I__3579 (
            .O(N__24830),
            .I(N__24827));
    Odrv12 I__3578 (
            .O(N__24827),
            .I(\pid_alt.error_d_regZ0Z_20 ));
    InMux I__3577 (
            .O(N__24824),
            .I(N__24821));
    LocalMux I__3576 (
            .O(N__24821),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ));
    CascadeMux I__3575 (
            .O(N__24818),
            .I(\pid_alt.un1_pid_prereg_236_1_cascade_ ));
    CascadeMux I__3574 (
            .O(N__24815),
            .I(N__24812));
    InMux I__3573 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__3572 (
            .O(N__24809),
            .I(N__24806));
    Odrv4 I__3571 (
            .O(N__24806),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ));
    InMux I__3570 (
            .O(N__24803),
            .I(N__24793));
    InMux I__3569 (
            .O(N__24802),
            .I(N__24793));
    InMux I__3568 (
            .O(N__24801),
            .I(N__24793));
    CascadeMux I__3567 (
            .O(N__24800),
            .I(N__24790));
    LocalMux I__3566 (
            .O(N__24793),
            .I(N__24787));
    InMux I__3565 (
            .O(N__24790),
            .I(N__24782));
    Span4Mux_h I__3564 (
            .O(N__24787),
            .I(N__24779));
    InMux I__3563 (
            .O(N__24786),
            .I(N__24774));
    InMux I__3562 (
            .O(N__24785),
            .I(N__24774));
    LocalMux I__3561 (
            .O(N__24782),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    Odrv4 I__3560 (
            .O(N__24779),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    LocalMux I__3559 (
            .O(N__24774),
            .I(\pid_alt.un1_pid_prereg_236_1 ));
    CascadeMux I__3558 (
            .O(N__24767),
            .I(N__24764));
    InMux I__3557 (
            .O(N__24764),
            .I(N__24755));
    InMux I__3556 (
            .O(N__24763),
            .I(N__24755));
    InMux I__3555 (
            .O(N__24762),
            .I(N__24755));
    LocalMux I__3554 (
            .O(N__24755),
            .I(N__24751));
    InMux I__3553 (
            .O(N__24754),
            .I(N__24747));
    Span4Mux_h I__3552 (
            .O(N__24751),
            .I(N__24744));
    InMux I__3551 (
            .O(N__24750),
            .I(N__24741));
    LocalMux I__3550 (
            .O(N__24747),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    Odrv4 I__3549 (
            .O(N__24744),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    LocalMux I__3548 (
            .O(N__24741),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ));
    CascadeMux I__3547 (
            .O(N__24734),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_ ));
    InMux I__3546 (
            .O(N__24731),
            .I(N__24717));
    InMux I__3545 (
            .O(N__24730),
            .I(N__24717));
    InMux I__3544 (
            .O(N__24729),
            .I(N__24717));
    InMux I__3543 (
            .O(N__24728),
            .I(N__24717));
    InMux I__3542 (
            .O(N__24727),
            .I(N__24714));
    InMux I__3541 (
            .O(N__24726),
            .I(N__24711));
    LocalMux I__3540 (
            .O(N__24717),
            .I(N__24708));
    LocalMux I__3539 (
            .O(N__24714),
            .I(N__24703));
    LocalMux I__3538 (
            .O(N__24711),
            .I(N__24703));
    Span4Mux_s3_h I__3537 (
            .O(N__24708),
            .I(N__24698));
    Span4Mux_h I__3536 (
            .O(N__24703),
            .I(N__24698));
    Odrv4 I__3535 (
            .O(N__24698),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ));
    InMux I__3534 (
            .O(N__24695),
            .I(N__24692));
    LocalMux I__3533 (
            .O(N__24692),
            .I(\pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ));
    InMux I__3532 (
            .O(N__24689),
            .I(N__24686));
    LocalMux I__3531 (
            .O(N__24686),
            .I(drone_altitude_1));
    InMux I__3530 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3529 (
            .O(N__24680),
            .I(drone_altitude_2));
    InMux I__3528 (
            .O(N__24677),
            .I(N__24674));
    LocalMux I__3527 (
            .O(N__24674),
            .I(drone_altitude_3));
    CascadeMux I__3526 (
            .O(N__24671),
            .I(N__24667));
    CascadeMux I__3525 (
            .O(N__24670),
            .I(N__24664));
    InMux I__3524 (
            .O(N__24667),
            .I(N__24661));
    InMux I__3523 (
            .O(N__24664),
            .I(N__24658));
    LocalMux I__3522 (
            .O(N__24661),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    LocalMux I__3521 (
            .O(N__24658),
            .I(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ));
    InMux I__3520 (
            .O(N__24653),
            .I(N__24644));
    InMux I__3519 (
            .O(N__24652),
            .I(N__24644));
    InMux I__3518 (
            .O(N__24651),
            .I(N__24644));
    LocalMux I__3517 (
            .O(N__24644),
            .I(N__24641));
    Span4Mux_h I__3516 (
            .O(N__24641),
            .I(N__24638));
    Span4Mux_v I__3515 (
            .O(N__24638),
            .I(N__24635));
    Span4Mux_v I__3514 (
            .O(N__24635),
            .I(N__24632));
    Odrv4 I__3513 (
            .O(N__24632),
            .I(\pid_alt.error_d_regZ0Z_7 ));
    CascadeMux I__3512 (
            .O(N__24629),
            .I(N__24626));
    InMux I__3511 (
            .O(N__24626),
            .I(N__24620));
    InMux I__3510 (
            .O(N__24625),
            .I(N__24620));
    LocalMux I__3509 (
            .O(N__24620),
            .I(\pid_alt.error_d_reg_prevZ0Z_7 ));
    InMux I__3508 (
            .O(N__24617),
            .I(N__24611));
    InMux I__3507 (
            .O(N__24616),
            .I(N__24611));
    LocalMux I__3506 (
            .O(N__24611),
            .I(N__24608));
    Span4Mux_h I__3505 (
            .O(N__24608),
            .I(N__24605));
    Span4Mux_v I__3504 (
            .O(N__24605),
            .I(N__24602));
    Odrv4 I__3503 (
            .O(N__24602),
            .I(\pid_alt.error_p_regZ0Z_7 ));
    CascadeMux I__3502 (
            .O(N__24599),
            .I(N__24596));
    InMux I__3501 (
            .O(N__24596),
            .I(N__24593));
    LocalMux I__3500 (
            .O(N__24593),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ));
    InMux I__3499 (
            .O(N__24590),
            .I(N__24584));
    InMux I__3498 (
            .O(N__24589),
            .I(N__24584));
    LocalMux I__3497 (
            .O(N__24584),
            .I(N__24581));
    Span4Mux_h I__3496 (
            .O(N__24581),
            .I(N__24578));
    Odrv4 I__3495 (
            .O(N__24578),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ));
    CascadeMux I__3494 (
            .O(N__24575),
            .I(N__24571));
    InMux I__3493 (
            .O(N__24574),
            .I(N__24568));
    InMux I__3492 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__3491 (
            .O(N__24568),
            .I(N__24560));
    LocalMux I__3490 (
            .O(N__24565),
            .I(N__24560));
    Span4Mux_v I__3489 (
            .O(N__24560),
            .I(N__24557));
    Odrv4 I__3488 (
            .O(N__24557),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ));
    CascadeMux I__3487 (
            .O(N__24554),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ));
    InMux I__3486 (
            .O(N__24551),
            .I(N__24545));
    InMux I__3485 (
            .O(N__24550),
            .I(N__24545));
    LocalMux I__3484 (
            .O(N__24545),
            .I(N__24541));
    InMux I__3483 (
            .O(N__24544),
            .I(N__24538));
    Span4Mux_h I__3482 (
            .O(N__24541),
            .I(N__24535));
    LocalMux I__3481 (
            .O(N__24538),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    Odrv4 I__3480 (
            .O(N__24535),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ));
    InMux I__3479 (
            .O(N__24530),
            .I(N__24527));
    LocalMux I__3478 (
            .O(N__24527),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ));
    InMux I__3477 (
            .O(N__24524),
            .I(N__24521));
    LocalMux I__3476 (
            .O(N__24521),
            .I(\pid_alt.pid_preregZ0Z_20 ));
    InMux I__3475 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__3474 (
            .O(N__24515),
            .I(\pid_alt.pid_preregZ0Z_19 ));
    CascadeMux I__3473 (
            .O(N__24512),
            .I(N__24509));
    InMux I__3472 (
            .O(N__24509),
            .I(N__24506));
    LocalMux I__3471 (
            .O(N__24506),
            .I(\pid_alt.pid_preregZ0Z_22 ));
    InMux I__3470 (
            .O(N__24503),
            .I(N__24500));
    LocalMux I__3469 (
            .O(N__24500),
            .I(\pid_alt.pid_preregZ0Z_17 ));
    InMux I__3468 (
            .O(N__24497),
            .I(N__24494));
    LocalMux I__3467 (
            .O(N__24494),
            .I(\pid_alt.pid_preregZ0Z_21 ));
    InMux I__3466 (
            .O(N__24491),
            .I(N__24488));
    LocalMux I__3465 (
            .O(N__24488),
            .I(\pid_alt.pid_preregZ0Z_15 ));
    CascadeMux I__3464 (
            .O(N__24485),
            .I(N__24482));
    InMux I__3463 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__3462 (
            .O(N__24479),
            .I(\pid_alt.pid_preregZ0Z_23 ));
    InMux I__3461 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__3460 (
            .O(N__24473),
            .I(\pid_alt.pid_preregZ0Z_18 ));
    InMux I__3459 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__3458 (
            .O(N__24467),
            .I(N__24463));
    InMux I__3457 (
            .O(N__24466),
            .I(N__24460));
    Span4Mux_v I__3456 (
            .O(N__24463),
            .I(N__24457));
    LocalMux I__3455 (
            .O(N__24460),
            .I(N__24454));
    Span4Mux_h I__3454 (
            .O(N__24457),
            .I(N__24449));
    Span4Mux_v I__3453 (
            .O(N__24454),
            .I(N__24449));
    Odrv4 I__3452 (
            .O(N__24449),
            .I(\pid_alt.error_p_regZ0Z_19 ));
    InMux I__3451 (
            .O(N__24446),
            .I(N__24443));
    LocalMux I__3450 (
            .O(N__24443),
            .I(\pid_alt.error_i_acumm_preregZ0Z_15 ));
    InMux I__3449 (
            .O(N__24440),
            .I(N__24437));
    LocalMux I__3448 (
            .O(N__24437),
            .I(\pid_alt.error_i_acumm_preregZ0Z_14 ));
    InMux I__3447 (
            .O(N__24434),
            .I(N__24431));
    LocalMux I__3446 (
            .O(N__24431),
            .I(N__24428));
    Span4Mux_v I__3445 (
            .O(N__24428),
            .I(N__24425));
    Odrv4 I__3444 (
            .O(N__24425),
            .I(\pid_alt.un1_reset_1_i_a5_0_9 ));
    InMux I__3443 (
            .O(N__24422),
            .I(N__24419));
    LocalMux I__3442 (
            .O(N__24419),
            .I(N__24416));
    Span4Mux_h I__3441 (
            .O(N__24416),
            .I(N__24413));
    Odrv4 I__3440 (
            .O(N__24413),
            .I(\pid_alt.un1_reset_1_i_a5_0_8 ));
    CascadeMux I__3439 (
            .O(N__24410),
            .I(\pid_alt.N_557_cascade_ ));
    InMux I__3438 (
            .O(N__24407),
            .I(N__24404));
    LocalMux I__3437 (
            .O(N__24404),
            .I(\pid_alt.un1_reset_1_i_a5_0_10 ));
    CascadeMux I__3436 (
            .O(N__24401),
            .I(\pid_alt.N_304_cascade_ ));
    CascadeMux I__3435 (
            .O(N__24398),
            .I(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_ ));
    InMux I__3434 (
            .O(N__24395),
            .I(N__24392));
    LocalMux I__3433 (
            .O(N__24392),
            .I(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ));
    InMux I__3432 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__3431 (
            .O(N__24386),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ));
    CascadeMux I__3430 (
            .O(N__24383),
            .I(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ));
    InMux I__3429 (
            .O(N__24380),
            .I(N__24374));
    InMux I__3428 (
            .O(N__24379),
            .I(N__24374));
    LocalMux I__3427 (
            .O(N__24374),
            .I(N__24370));
    InMux I__3426 (
            .O(N__24373),
            .I(N__24367));
    Span4Mux_h I__3425 (
            .O(N__24370),
            .I(N__24364));
    LocalMux I__3424 (
            .O(N__24367),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    Odrv4 I__3423 (
            .O(N__24364),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ));
    InMux I__3422 (
            .O(N__24359),
            .I(N__24355));
    CascadeMux I__3421 (
            .O(N__24358),
            .I(N__24352));
    LocalMux I__3420 (
            .O(N__24355),
            .I(N__24349));
    InMux I__3419 (
            .O(N__24352),
            .I(N__24346));
    Odrv4 I__3418 (
            .O(N__24349),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    LocalMux I__3417 (
            .O(N__24346),
            .I(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ));
    InMux I__3416 (
            .O(N__24341),
            .I(N__24338));
    LocalMux I__3415 (
            .O(N__24338),
            .I(N__24334));
    InMux I__3414 (
            .O(N__24337),
            .I(N__24331));
    Span4Mux_v I__3413 (
            .O(N__24334),
            .I(N__24328));
    LocalMux I__3412 (
            .O(N__24331),
            .I(N__24325));
    Span4Mux_h I__3411 (
            .O(N__24328),
            .I(N__24322));
    Odrv12 I__3410 (
            .O(N__24325),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    Odrv4 I__3409 (
            .O(N__24322),
            .I(\pid_alt.error_p_regZ0Z_8 ));
    InMux I__3408 (
            .O(N__24317),
            .I(N__24314));
    LocalMux I__3407 (
            .O(N__24314),
            .I(N__24311));
    Span4Mux_h I__3406 (
            .O(N__24311),
            .I(N__24307));
    InMux I__3405 (
            .O(N__24310),
            .I(N__24304));
    Span4Mux_v I__3404 (
            .O(N__24307),
            .I(N__24301));
    LocalMux I__3403 (
            .O(N__24304),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    Odrv4 I__3402 (
            .O(N__24301),
            .I(\pid_alt.error_d_reg_prevZ0Z_8 ));
    InMux I__3401 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__3400 (
            .O(N__24293),
            .I(N__24288));
    InMux I__3399 (
            .O(N__24292),
            .I(N__24283));
    InMux I__3398 (
            .O(N__24291),
            .I(N__24283));
    Span4Mux_v I__3397 (
            .O(N__24288),
            .I(N__24280));
    LocalMux I__3396 (
            .O(N__24283),
            .I(N__24277));
    Span4Mux_v I__3395 (
            .O(N__24280),
            .I(N__24274));
    Span12Mux_v I__3394 (
            .O(N__24277),
            .I(N__24271));
    Span4Mux_v I__3393 (
            .O(N__24274),
            .I(N__24268));
    Odrv12 I__3392 (
            .O(N__24271),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    Odrv4 I__3391 (
            .O(N__24268),
            .I(\pid_alt.error_d_regZ0Z_8 ));
    InMux I__3390 (
            .O(N__24263),
            .I(N__24257));
    InMux I__3389 (
            .O(N__24262),
            .I(N__24257));
    LocalMux I__3388 (
            .O(N__24257),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ));
    InMux I__3387 (
            .O(N__24254),
            .I(N__24251));
    LocalMux I__3386 (
            .O(N__24251),
            .I(N__24248));
    Span4Mux_v I__3385 (
            .O(N__24248),
            .I(N__24243));
    InMux I__3384 (
            .O(N__24247),
            .I(N__24240));
    CascadeMux I__3383 (
            .O(N__24246),
            .I(N__24237));
    Span4Mux_v I__3382 (
            .O(N__24243),
            .I(N__24232));
    LocalMux I__3381 (
            .O(N__24240),
            .I(N__24232));
    InMux I__3380 (
            .O(N__24237),
            .I(N__24229));
    Odrv4 I__3379 (
            .O(N__24232),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    LocalMux I__3378 (
            .O(N__24229),
            .I(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ));
    InMux I__3377 (
            .O(N__24224),
            .I(N__24221));
    LocalMux I__3376 (
            .O(N__24221),
            .I(N__24216));
    InMux I__3375 (
            .O(N__24220),
            .I(N__24211));
    InMux I__3374 (
            .O(N__24219),
            .I(N__24211));
    Span4Mux_h I__3373 (
            .O(N__24216),
            .I(N__24208));
    LocalMux I__3372 (
            .O(N__24211),
            .I(N__24205));
    Odrv4 I__3371 (
            .O(N__24208),
            .I(\pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12 ));
    Odrv4 I__3370 (
            .O(N__24205),
            .I(\pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12 ));
    InMux I__3369 (
            .O(N__24200),
            .I(N__24196));
    CascadeMux I__3368 (
            .O(N__24199),
            .I(N__24193));
    LocalMux I__3367 (
            .O(N__24196),
            .I(N__24190));
    InMux I__3366 (
            .O(N__24193),
            .I(N__24187));
    Odrv4 I__3365 (
            .O(N__24190),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    LocalMux I__3364 (
            .O(N__24187),
            .I(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ));
    InMux I__3363 (
            .O(N__24182),
            .I(N__24179));
    LocalMux I__3362 (
            .O(N__24179),
            .I(N__24174));
    InMux I__3361 (
            .O(N__24178),
            .I(N__24171));
    CascadeMux I__3360 (
            .O(N__24177),
            .I(N__24168));
    Span4Mux_v I__3359 (
            .O(N__24174),
            .I(N__24163));
    LocalMux I__3358 (
            .O(N__24171),
            .I(N__24163));
    InMux I__3357 (
            .O(N__24168),
            .I(N__24160));
    Odrv4 I__3356 (
            .O(N__24163),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    LocalMux I__3355 (
            .O(N__24160),
            .I(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ));
    InMux I__3354 (
            .O(N__24155),
            .I(N__24152));
    LocalMux I__3353 (
            .O(N__24152),
            .I(N__24147));
    InMux I__3352 (
            .O(N__24151),
            .I(N__24142));
    InMux I__3351 (
            .O(N__24150),
            .I(N__24142));
    Span4Mux_h I__3350 (
            .O(N__24147),
            .I(N__24139));
    LocalMux I__3349 (
            .O(N__24142),
            .I(N__24136));
    Odrv4 I__3348 (
            .O(N__24139),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    Odrv4 I__3347 (
            .O(N__24136),
            .I(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ));
    InMux I__3346 (
            .O(N__24131),
            .I(N__24128));
    LocalMux I__3345 (
            .O(N__24128),
            .I(N__24124));
    InMux I__3344 (
            .O(N__24127),
            .I(N__24121));
    Span4Mux_h I__3343 (
            .O(N__24124),
            .I(N__24117));
    LocalMux I__3342 (
            .O(N__24121),
            .I(N__24114));
    InMux I__3341 (
            .O(N__24120),
            .I(N__24111));
    Odrv4 I__3340 (
            .O(N__24117),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    Odrv4 I__3339 (
            .O(N__24114),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    LocalMux I__3338 (
            .O(N__24111),
            .I(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ));
    InMux I__3337 (
            .O(N__24104),
            .I(N__24101));
    LocalMux I__3336 (
            .O(N__24101),
            .I(N__24096));
    InMux I__3335 (
            .O(N__24100),
            .I(N__24093));
    InMux I__3334 (
            .O(N__24099),
            .I(N__24090));
    Span4Mux_h I__3333 (
            .O(N__24096),
            .I(N__24087));
    LocalMux I__3332 (
            .O(N__24093),
            .I(\pid_alt.error_i_acumm7lto12 ));
    LocalMux I__3331 (
            .O(N__24090),
            .I(\pid_alt.error_i_acumm7lto12 ));
    Odrv4 I__3330 (
            .O(N__24087),
            .I(\pid_alt.error_i_acumm7lto12 ));
    InMux I__3329 (
            .O(N__24080),
            .I(N__24077));
    LocalMux I__3328 (
            .O(N__24077),
            .I(N__24074));
    Odrv4 I__3327 (
            .O(N__24074),
            .I(\pid_alt.error_i_acummZ0Z_12 ));
    InMux I__3326 (
            .O(N__24071),
            .I(N__24068));
    LocalMux I__3325 (
            .O(N__24068),
            .I(N__24064));
    InMux I__3324 (
            .O(N__24067),
            .I(N__24061));
    Odrv4 I__3323 (
            .O(N__24064),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    LocalMux I__3322 (
            .O(N__24061),
            .I(\pid_alt.error_i_acumm_preregZ0Z_3 ));
    InMux I__3321 (
            .O(N__24056),
            .I(N__24052));
    InMux I__3320 (
            .O(N__24055),
            .I(N__24049));
    LocalMux I__3319 (
            .O(N__24052),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    LocalMux I__3318 (
            .O(N__24049),
            .I(\pid_alt.error_i_acumm_preregZ0Z_1 ));
    CascadeMux I__3317 (
            .O(N__24044),
            .I(N__24040));
    InMux I__3316 (
            .O(N__24043),
            .I(N__24037));
    InMux I__3315 (
            .O(N__24040),
            .I(N__24034));
    LocalMux I__3314 (
            .O(N__24037),
            .I(N__24031));
    LocalMux I__3313 (
            .O(N__24034),
            .I(N__24027));
    Span12Mux_s11_v I__3312 (
            .O(N__24031),
            .I(N__24024));
    InMux I__3311 (
            .O(N__24030),
            .I(N__24021));
    Span4Mux_h I__3310 (
            .O(N__24027),
            .I(N__24018));
    Odrv12 I__3309 (
            .O(N__24024),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    LocalMux I__3308 (
            .O(N__24021),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    Odrv4 I__3307 (
            .O(N__24018),
            .I(\pid_alt.error_i_acumm_preregZ0Z_7 ));
    InMux I__3306 (
            .O(N__24011),
            .I(N__24008));
    LocalMux I__3305 (
            .O(N__24008),
            .I(N__24004));
    InMux I__3304 (
            .O(N__24007),
            .I(N__24001));
    Odrv4 I__3303 (
            .O(N__24004),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    LocalMux I__3302 (
            .O(N__24001),
            .I(\pid_alt.error_i_acumm_preregZ0Z_2 ));
    CascadeMux I__3301 (
            .O(N__23996),
            .I(\pid_alt.un1_reset_1_i_a5_0_7_cascade_ ));
    CascadeMux I__3300 (
            .O(N__23993),
            .I(N__23990));
    InMux I__3299 (
            .O(N__23990),
            .I(N__23984));
    InMux I__3298 (
            .O(N__23989),
            .I(N__23984));
    LocalMux I__3297 (
            .O(N__23984),
            .I(\pid_alt.error_d_reg_prevZ0Z_12 ));
    CascadeMux I__3296 (
            .O(N__23981),
            .I(N__23978));
    InMux I__3295 (
            .O(N__23978),
            .I(N__23974));
    CascadeMux I__3294 (
            .O(N__23977),
            .I(N__23971));
    LocalMux I__3293 (
            .O(N__23974),
            .I(N__23968));
    InMux I__3292 (
            .O(N__23971),
            .I(N__23965));
    Span4Mux_v I__3291 (
            .O(N__23968),
            .I(N__23962));
    LocalMux I__3290 (
            .O(N__23965),
            .I(N__23959));
    Odrv4 I__3289 (
            .O(N__23962),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    Odrv12 I__3288 (
            .O(N__23959),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ));
    InMux I__3287 (
            .O(N__23954),
            .I(N__23951));
    LocalMux I__3286 (
            .O(N__23951),
            .I(N__23948));
    Span4Mux_v I__3285 (
            .O(N__23948),
            .I(N__23945));
    Odrv4 I__3284 (
            .O(N__23945),
            .I(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ));
    InMux I__3283 (
            .O(N__23942),
            .I(N__23939));
    LocalMux I__3282 (
            .O(N__23939),
            .I(N__23936));
    Span4Mux_v I__3281 (
            .O(N__23936),
            .I(N__23932));
    InMux I__3280 (
            .O(N__23935),
            .I(N__23929));
    Span4Mux_h I__3279 (
            .O(N__23932),
            .I(N__23924));
    LocalMux I__3278 (
            .O(N__23929),
            .I(N__23924));
    Span4Mux_v I__3277 (
            .O(N__23924),
            .I(N__23921));
    Span4Mux_v I__3276 (
            .O(N__23921),
            .I(N__23918));
    Odrv4 I__3275 (
            .O(N__23918),
            .I(\pid_alt.error_p_regZ0Z_10 ));
    InMux I__3274 (
            .O(N__23915),
            .I(N__23911));
    InMux I__3273 (
            .O(N__23914),
            .I(N__23908));
    LocalMux I__3272 (
            .O(N__23911),
            .I(N__23905));
    LocalMux I__3271 (
            .O(N__23908),
            .I(N__23902));
    Span4Mux_h I__3270 (
            .O(N__23905),
            .I(N__23899));
    Span4Mux_v I__3269 (
            .O(N__23902),
            .I(N__23896));
    Odrv4 I__3268 (
            .O(N__23899),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    Odrv4 I__3267 (
            .O(N__23896),
            .I(\pid_alt.error_d_reg_prevZ0Z_10 ));
    InMux I__3266 (
            .O(N__23891),
            .I(N__23886));
    InMux I__3265 (
            .O(N__23890),
            .I(N__23883));
    InMux I__3264 (
            .O(N__23889),
            .I(N__23880));
    LocalMux I__3263 (
            .O(N__23886),
            .I(N__23877));
    LocalMux I__3262 (
            .O(N__23883),
            .I(N__23874));
    LocalMux I__3261 (
            .O(N__23880),
            .I(N__23867));
    Span4Mux_h I__3260 (
            .O(N__23877),
            .I(N__23867));
    Span4Mux_v I__3259 (
            .O(N__23874),
            .I(N__23867));
    Span4Mux_v I__3258 (
            .O(N__23867),
            .I(N__23864));
    Odrv4 I__3257 (
            .O(N__23864),
            .I(\pid_alt.error_d_regZ0Z_10 ));
    InMux I__3256 (
            .O(N__23861),
            .I(N__23858));
    LocalMux I__3255 (
            .O(N__23858),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ));
    CascadeMux I__3254 (
            .O(N__23855),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ));
    CascadeMux I__3253 (
            .O(N__23852),
            .I(N__23849));
    InMux I__3252 (
            .O(N__23849),
            .I(N__23846));
    LocalMux I__3251 (
            .O(N__23846),
            .I(N__23842));
    InMux I__3250 (
            .O(N__23845),
            .I(N__23839));
    Span4Mux_h I__3249 (
            .O(N__23842),
            .I(N__23836));
    LocalMux I__3248 (
            .O(N__23839),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    Odrv4 I__3247 (
            .O(N__23836),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ));
    InMux I__3246 (
            .O(N__23831),
            .I(N__23825));
    InMux I__3245 (
            .O(N__23830),
            .I(N__23825));
    LocalMux I__3244 (
            .O(N__23825),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ));
    InMux I__3243 (
            .O(N__23822),
            .I(N__23813));
    InMux I__3242 (
            .O(N__23821),
            .I(N__23813));
    InMux I__3241 (
            .O(N__23820),
            .I(N__23813));
    LocalMux I__3240 (
            .O(N__23813),
            .I(N__23810));
    Span4Mux_v I__3239 (
            .O(N__23810),
            .I(N__23807));
    Span4Mux_v I__3238 (
            .O(N__23807),
            .I(N__23804));
    Odrv4 I__3237 (
            .O(N__23804),
            .I(\pid_alt.error_d_regZ0Z_11 ));
    CascadeMux I__3236 (
            .O(N__23801),
            .I(N__23798));
    InMux I__3235 (
            .O(N__23798),
            .I(N__23792));
    InMux I__3234 (
            .O(N__23797),
            .I(N__23792));
    LocalMux I__3233 (
            .O(N__23792),
            .I(\pid_alt.error_d_reg_prevZ0Z_11 ));
    InMux I__3232 (
            .O(N__23789),
            .I(N__23783));
    InMux I__3231 (
            .O(N__23788),
            .I(N__23783));
    LocalMux I__3230 (
            .O(N__23783),
            .I(N__23780));
    Span12Mux_v I__3229 (
            .O(N__23780),
            .I(N__23777));
    Odrv12 I__3228 (
            .O(N__23777),
            .I(\pid_alt.error_p_regZ0Z_11 ));
    InMux I__3227 (
            .O(N__23774),
            .I(N__23768));
    InMux I__3226 (
            .O(N__23773),
            .I(N__23768));
    LocalMux I__3225 (
            .O(N__23768),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ));
    InMux I__3224 (
            .O(N__23765),
            .I(N__23756));
    InMux I__3223 (
            .O(N__23764),
            .I(N__23756));
    InMux I__3222 (
            .O(N__23763),
            .I(N__23756));
    LocalMux I__3221 (
            .O(N__23756),
            .I(N__23753));
    Span4Mux_v I__3220 (
            .O(N__23753),
            .I(N__23750));
    Odrv4 I__3219 (
            .O(N__23750),
            .I(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ));
    InMux I__3218 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__3217 (
            .O(N__23744),
            .I(N__23741));
    Span4Mux_v I__3216 (
            .O(N__23741),
            .I(N__23737));
    CascadeMux I__3215 (
            .O(N__23740),
            .I(N__23733));
    Span4Mux_v I__3214 (
            .O(N__23737),
            .I(N__23730));
    InMux I__3213 (
            .O(N__23736),
            .I(N__23725));
    InMux I__3212 (
            .O(N__23733),
            .I(N__23725));
    Span4Mux_v I__3211 (
            .O(N__23730),
            .I(N__23720));
    LocalMux I__3210 (
            .O(N__23725),
            .I(N__23720));
    Odrv4 I__3209 (
            .O(N__23720),
            .I(\pid_alt.error_i_acumm_preregZ0Z_11 ));
    InMux I__3208 (
            .O(N__23717),
            .I(N__23714));
    LocalMux I__3207 (
            .O(N__23714),
            .I(N__23710));
    InMux I__3206 (
            .O(N__23713),
            .I(N__23706));
    Span4Mux_v I__3205 (
            .O(N__23710),
            .I(N__23701));
    InMux I__3204 (
            .O(N__23709),
            .I(N__23698));
    LocalMux I__3203 (
            .O(N__23706),
            .I(N__23695));
    InMux I__3202 (
            .O(N__23705),
            .I(N__23690));
    InMux I__3201 (
            .O(N__23704),
            .I(N__23690));
    Odrv4 I__3200 (
            .O(N__23701),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    LocalMux I__3199 (
            .O(N__23698),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    Odrv4 I__3198 (
            .O(N__23695),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    LocalMux I__3197 (
            .O(N__23690),
            .I(\pid_alt.error_d_regZ0Z_0 ));
    InMux I__3196 (
            .O(N__23681),
            .I(N__23678));
    LocalMux I__3195 (
            .O(N__23678),
            .I(N__23675));
    Span4Mux_v I__3194 (
            .O(N__23675),
            .I(N__23672));
    Odrv4 I__3193 (
            .O(N__23672),
            .I(\pid_alt.error_d_reg_prevZ0Z_0 ));
    CascadeMux I__3192 (
            .O(N__23669),
            .I(N__23666));
    InMux I__3191 (
            .O(N__23666),
            .I(N__23663));
    LocalMux I__3190 (
            .O(N__23663),
            .I(N__23660));
    Odrv4 I__3189 (
            .O(N__23660),
            .I(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ));
    InMux I__3188 (
            .O(N__23657),
            .I(N__23652));
    InMux I__3187 (
            .O(N__23656),
            .I(N__23647));
    InMux I__3186 (
            .O(N__23655),
            .I(N__23644));
    LocalMux I__3185 (
            .O(N__23652),
            .I(N__23641));
    InMux I__3184 (
            .O(N__23651),
            .I(N__23638));
    InMux I__3183 (
            .O(N__23650),
            .I(N__23635));
    LocalMux I__3182 (
            .O(N__23647),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__3181 (
            .O(N__23644),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    Odrv4 I__3180 (
            .O(N__23641),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__3179 (
            .O(N__23638),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    LocalMux I__3178 (
            .O(N__23635),
            .I(\Commands_frame_decoder.stateZ0Z_1 ));
    CascadeMux I__3177 (
            .O(N__23624),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ));
    InMux I__3176 (
            .O(N__23621),
            .I(N__23618));
    LocalMux I__3175 (
            .O(N__23618),
            .I(N__23615));
    Odrv4 I__3174 (
            .O(N__23615),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_3_2 ));
    InMux I__3173 (
            .O(N__23612),
            .I(N__23608));
    InMux I__3172 (
            .O(N__23611),
            .I(N__23605));
    LocalMux I__3171 (
            .O(N__23608),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    LocalMux I__3170 (
            .O(N__23605),
            .I(\Commands_frame_decoder.stateZ0Z_5 ));
    CascadeMux I__3169 (
            .O(N__23600),
            .I(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ));
    InMux I__3168 (
            .O(N__23597),
            .I(N__23594));
    LocalMux I__3167 (
            .O(N__23594),
            .I(N__23589));
    InMux I__3166 (
            .O(N__23593),
            .I(N__23584));
    InMux I__3165 (
            .O(N__23592),
            .I(N__23584));
    Span4Mux_h I__3164 (
            .O(N__23589),
            .I(N__23579));
    LocalMux I__3163 (
            .O(N__23584),
            .I(N__23579));
    Span4Mux_h I__3162 (
            .O(N__23579),
            .I(N__23576));
    Span4Mux_v I__3161 (
            .O(N__23576),
            .I(N__23573));
    Odrv4 I__3160 (
            .O(N__23573),
            .I(\pid_alt.error_d_regZ0Z_12 ));
    InMux I__3159 (
            .O(N__23570),
            .I(N__23567));
    LocalMux I__3158 (
            .O(N__23567),
            .I(N__23564));
    Odrv4 I__3157 (
            .O(N__23564),
            .I(\Commands_frame_decoder.N_418 ));
    InMux I__3156 (
            .O(N__23561),
            .I(N__23555));
    InMux I__3155 (
            .O(N__23560),
            .I(N__23555));
    LocalMux I__3154 (
            .O(N__23555),
            .I(\Commands_frame_decoder.N_382_2 ));
    CascadeMux I__3153 (
            .O(N__23552),
            .I(\Commands_frame_decoder.N_383_cascade_ ));
    CascadeMux I__3152 (
            .O(N__23549),
            .I(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ));
    InMux I__3151 (
            .O(N__23546),
            .I(N__23542));
    InMux I__3150 (
            .O(N__23545),
            .I(N__23539));
    LocalMux I__3149 (
            .O(N__23542),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    LocalMux I__3148 (
            .O(N__23539),
            .I(\Commands_frame_decoder.stateZ0Z_0 ));
    InMux I__3147 (
            .O(N__23534),
            .I(N__23530));
    InMux I__3146 (
            .O(N__23533),
            .I(N__23526));
    LocalMux I__3145 (
            .O(N__23530),
            .I(N__23523));
    InMux I__3144 (
            .O(N__23529),
            .I(N__23520));
    LocalMux I__3143 (
            .O(N__23526),
            .I(N__23515));
    Span4Mux_h I__3142 (
            .O(N__23523),
            .I(N__23515));
    LocalMux I__3141 (
            .O(N__23520),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    Odrv4 I__3140 (
            .O(N__23515),
            .I(\Commands_frame_decoder.stateZ0Z_11 ));
    InMux I__3139 (
            .O(N__23510),
            .I(N__23506));
    InMux I__3138 (
            .O(N__23509),
            .I(N__23503));
    LocalMux I__3137 (
            .O(N__23506),
            .I(N__23498));
    LocalMux I__3136 (
            .O(N__23503),
            .I(N__23498));
    Odrv4 I__3135 (
            .O(N__23498),
            .I(frame_decoder_CH4data_7));
    InMux I__3134 (
            .O(N__23495),
            .I(N__23492));
    LocalMux I__3133 (
            .O(N__23492),
            .I(N__23489));
    Span4Mux_v I__3132 (
            .O(N__23489),
            .I(N__23486));
    Span4Mux_h I__3131 (
            .O(N__23486),
            .I(N__23483));
    Odrv4 I__3130 (
            .O(N__23483),
            .I(\pid_side.error_8 ));
    InMux I__3129 (
            .O(N__23480),
            .I(bfn_4_22_0_));
    InMux I__3128 (
            .O(N__23477),
            .I(N__23474));
    LocalMux I__3127 (
            .O(N__23474),
            .I(N__23471));
    Odrv4 I__3126 (
            .O(N__23471),
            .I(drone_H_disp_side_i_9));
    InMux I__3125 (
            .O(N__23468),
            .I(N__23465));
    LocalMux I__3124 (
            .O(N__23465),
            .I(N__23462));
    Span4Mux_v I__3123 (
            .O(N__23462),
            .I(N__23459));
    Span4Mux_h I__3122 (
            .O(N__23459),
            .I(N__23456));
    Odrv4 I__3121 (
            .O(N__23456),
            .I(\pid_side.error_9 ));
    InMux I__3120 (
            .O(N__23453),
            .I(\pid_side.error_cry_4 ));
    CascadeMux I__3119 (
            .O(N__23450),
            .I(N__23447));
    InMux I__3118 (
            .O(N__23447),
            .I(N__23444));
    LocalMux I__3117 (
            .O(N__23444),
            .I(N__23441));
    Odrv4 I__3116 (
            .O(N__23441),
            .I(drone_H_disp_side_i_10));
    InMux I__3115 (
            .O(N__23438),
            .I(N__23435));
    LocalMux I__3114 (
            .O(N__23435),
            .I(N__23432));
    Span4Mux_h I__3113 (
            .O(N__23432),
            .I(N__23429));
    Span4Mux_v I__3112 (
            .O(N__23429),
            .I(N__23426));
    Odrv4 I__3111 (
            .O(N__23426),
            .I(\pid_side.error_10 ));
    InMux I__3110 (
            .O(N__23423),
            .I(\pid_side.error_cry_5 ));
    InMux I__3109 (
            .O(N__23420),
            .I(N__23417));
    LocalMux I__3108 (
            .O(N__23417),
            .I(N__23414));
    Span4Mux_h I__3107 (
            .O(N__23414),
            .I(N__23411));
    Span4Mux_v I__3106 (
            .O(N__23411),
            .I(N__23408));
    Odrv4 I__3105 (
            .O(N__23408),
            .I(\pid_side.error_11 ));
    InMux I__3104 (
            .O(N__23405),
            .I(\pid_side.error_cry_6 ));
    InMux I__3103 (
            .O(N__23402),
            .I(N__23399));
    LocalMux I__3102 (
            .O(N__23399),
            .I(N__23396));
    Span4Mux_h I__3101 (
            .O(N__23396),
            .I(N__23393));
    Span4Mux_v I__3100 (
            .O(N__23393),
            .I(N__23390));
    Odrv4 I__3099 (
            .O(N__23390),
            .I(\pid_side.error_12 ));
    InMux I__3098 (
            .O(N__23387),
            .I(\pid_side.error_cry_7 ));
    InMux I__3097 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__3096 (
            .O(N__23381),
            .I(N__23378));
    Span4Mux_h I__3095 (
            .O(N__23378),
            .I(N__23375));
    Span4Mux_v I__3094 (
            .O(N__23375),
            .I(N__23372));
    Odrv4 I__3093 (
            .O(N__23372),
            .I(\pid_side.error_13 ));
    InMux I__3092 (
            .O(N__23369),
            .I(\pid_side.error_cry_8 ));
    InMux I__3091 (
            .O(N__23366),
            .I(N__23363));
    LocalMux I__3090 (
            .O(N__23363),
            .I(N__23360));
    Span4Mux_h I__3089 (
            .O(N__23360),
            .I(N__23357));
    Span4Mux_v I__3088 (
            .O(N__23357),
            .I(N__23354));
    Odrv4 I__3087 (
            .O(N__23354),
            .I(\pid_side.error_14 ));
    InMux I__3086 (
            .O(N__23351),
            .I(\pid_side.error_cry_9 ));
    InMux I__3085 (
            .O(N__23348),
            .I(\pid_side.error_cry_10 ));
    InMux I__3084 (
            .O(N__23345),
            .I(N__23342));
    LocalMux I__3083 (
            .O(N__23342),
            .I(N__23339));
    Span12Mux_s4_h I__3082 (
            .O(N__23339),
            .I(N__23336));
    Odrv12 I__3081 (
            .O(N__23336),
            .I(\pid_side.error_15 ));
    InMux I__3080 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3079 (
            .O(N__23330),
            .I(N__23327));
    Span4Mux_h I__3078 (
            .O(N__23327),
            .I(N__23324));
    Odrv4 I__3077 (
            .O(N__23324),
            .I(alt_kp_0));
    InMux I__3076 (
            .O(N__23321),
            .I(N__23318));
    LocalMux I__3075 (
            .O(N__23318),
            .I(\pid_side.error_axb_0 ));
    InMux I__3074 (
            .O(N__23315),
            .I(N__23312));
    LocalMux I__3073 (
            .O(N__23312),
            .I(N__23309));
    Span4Mux_s2_h I__3072 (
            .O(N__23309),
            .I(N__23306));
    Span4Mux_v I__3071 (
            .O(N__23306),
            .I(N__23303));
    Odrv4 I__3070 (
            .O(N__23303),
            .I(\pid_side.error_1 ));
    InMux I__3069 (
            .O(N__23300),
            .I(\pid_side.error_cry_0 ));
    InMux I__3068 (
            .O(N__23297),
            .I(N__23294));
    LocalMux I__3067 (
            .O(N__23294),
            .I(N__23291));
    Span4Mux_h I__3066 (
            .O(N__23291),
            .I(N__23288));
    Odrv4 I__3065 (
            .O(N__23288),
            .I(\pid_side.error_2 ));
    InMux I__3064 (
            .O(N__23285),
            .I(\pid_side.error_cry_1 ));
    InMux I__3063 (
            .O(N__23282),
            .I(N__23279));
    LocalMux I__3062 (
            .O(N__23279),
            .I(N__23276));
    Span4Mux_s1_h I__3061 (
            .O(N__23276),
            .I(N__23273));
    Span4Mux_h I__3060 (
            .O(N__23273),
            .I(N__23270));
    Odrv4 I__3059 (
            .O(N__23270),
            .I(\pid_side.error_3 ));
    InMux I__3058 (
            .O(N__23267),
            .I(\pid_side.error_cry_2 ));
    InMux I__3057 (
            .O(N__23264),
            .I(N__23261));
    LocalMux I__3056 (
            .O(N__23261),
            .I(N__23258));
    Span4Mux_h I__3055 (
            .O(N__23258),
            .I(N__23255));
    Odrv4 I__3054 (
            .O(N__23255),
            .I(\pid_side.error_4 ));
    InMux I__3053 (
            .O(N__23252),
            .I(\pid_side.error_cry_3 ));
    InMux I__3052 (
            .O(N__23249),
            .I(N__23246));
    LocalMux I__3051 (
            .O(N__23246),
            .I(N__23243));
    Span4Mux_h I__3050 (
            .O(N__23243),
            .I(N__23240));
    Odrv4 I__3049 (
            .O(N__23240),
            .I(\pid_side.error_5 ));
    InMux I__3048 (
            .O(N__23237),
            .I(\pid_side.error_cry_0_0 ));
    InMux I__3047 (
            .O(N__23234),
            .I(N__23231));
    LocalMux I__3046 (
            .O(N__23231),
            .I(N__23228));
    Span4Mux_s1_h I__3045 (
            .O(N__23228),
            .I(N__23225));
    Span4Mux_v I__3044 (
            .O(N__23225),
            .I(N__23222));
    Odrv4 I__3043 (
            .O(N__23222),
            .I(\pid_side.error_6 ));
    InMux I__3042 (
            .O(N__23219),
            .I(\pid_side.error_cry_1_0 ));
    InMux I__3041 (
            .O(N__23216),
            .I(N__23213));
    LocalMux I__3040 (
            .O(N__23213),
            .I(N__23210));
    Span4Mux_s1_h I__3039 (
            .O(N__23210),
            .I(N__23207));
    Span4Mux_v I__3038 (
            .O(N__23207),
            .I(N__23204));
    Odrv4 I__3037 (
            .O(N__23204),
            .I(\pid_side.error_7 ));
    InMux I__3036 (
            .O(N__23201),
            .I(\pid_side.error_cry_2_0 ));
    InMux I__3035 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__3034 (
            .O(N__23195),
            .I(N__23192));
    Odrv4 I__3033 (
            .O(N__23192),
            .I(drone_H_disp_side_i_8));
    CascadeMux I__3032 (
            .O(N__23189),
            .I(N__23186));
    InMux I__3031 (
            .O(N__23186),
            .I(N__23182));
    InMux I__3030 (
            .O(N__23185),
            .I(N__23179));
    LocalMux I__3029 (
            .O(N__23182),
            .I(N__23176));
    LocalMux I__3028 (
            .O(N__23179),
            .I(N__23173));
    Span4Mux_v I__3027 (
            .O(N__23176),
            .I(N__23170));
    Span4Mux_v I__3026 (
            .O(N__23173),
            .I(N__23167));
    Odrv4 I__3025 (
            .O(N__23170),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    Odrv4 I__3024 (
            .O(N__23167),
            .I(\pid_alt.error_d_reg_prev_i_0 ));
    InMux I__3023 (
            .O(N__23162),
            .I(N__23159));
    LocalMux I__3022 (
            .O(N__23159),
            .I(\dron_frame_decoder_1.drone_H_disp_side_8 ));
    InMux I__3021 (
            .O(N__23156),
            .I(N__23153));
    LocalMux I__3020 (
            .O(N__23153),
            .I(\dron_frame_decoder_1.drone_H_disp_side_9 ));
    InMux I__3019 (
            .O(N__23150),
            .I(N__23147));
    LocalMux I__3018 (
            .O(N__23147),
            .I(\dron_frame_decoder_1.drone_H_disp_side_10 ));
    InMux I__3017 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__3016 (
            .O(N__23141),
            .I(\pid_alt.error_axbZ0Z_1 ));
    InMux I__3015 (
            .O(N__23138),
            .I(N__23135));
    LocalMux I__3014 (
            .O(N__23135),
            .I(N__23132));
    Odrv4 I__3013 (
            .O(N__23132),
            .I(drone_altitude_12));
    CascadeMux I__3012 (
            .O(N__23129),
            .I(N__23126));
    InMux I__3011 (
            .O(N__23126),
            .I(N__23123));
    LocalMux I__3010 (
            .O(N__23123),
            .I(\pid_alt.error_axbZ0Z_12 ));
    InMux I__3009 (
            .O(N__23120),
            .I(N__23117));
    LocalMux I__3008 (
            .O(N__23117),
            .I(N__23114));
    Span4Mux_h I__3007 (
            .O(N__23114),
            .I(N__23111));
    Odrv4 I__3006 (
            .O(N__23111),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ));
    InMux I__3005 (
            .O(N__23108),
            .I(\pid_alt.un1_pid_prereg_0_cry_21 ));
    CascadeMux I__3004 (
            .O(N__23105),
            .I(N__23101));
    InMux I__3003 (
            .O(N__23104),
            .I(N__23098));
    InMux I__3002 (
            .O(N__23101),
            .I(N__23095));
    LocalMux I__3001 (
            .O(N__23098),
            .I(N__23092));
    LocalMux I__3000 (
            .O(N__23095),
            .I(N__23089));
    Span4Mux_v I__2999 (
            .O(N__23092),
            .I(N__23086));
    Span4Mux_h I__2998 (
            .O(N__23089),
            .I(N__23083));
    Odrv4 I__2997 (
            .O(N__23086),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ));
    Odrv4 I__2996 (
            .O(N__23083),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ));
    CascadeMux I__2995 (
            .O(N__23078),
            .I(N__23075));
    InMux I__2994 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__2993 (
            .O(N__23072),
            .I(N__23069));
    Span4Mux_v I__2992 (
            .O(N__23069),
            .I(N__23066));
    Odrv4 I__2991 (
            .O(N__23066),
            .I(\pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ));
    InMux I__2990 (
            .O(N__23063),
            .I(bfn_4_18_0_));
    InMux I__2989 (
            .O(N__23060),
            .I(\pid_alt.un1_pid_prereg_0_cry_23 ));
    InMux I__2988 (
            .O(N__23057),
            .I(N__23054));
    LocalMux I__2987 (
            .O(N__23054),
            .I(\pid_alt.error_axbZ0Z_13 ));
    InMux I__2986 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__2985 (
            .O(N__23048),
            .I(drone_altitude_13));
    InMux I__2984 (
            .O(N__23045),
            .I(N__23042));
    LocalMux I__2983 (
            .O(N__23042),
            .I(\pid_alt.error_axbZ0Z_14 ));
    InMux I__2982 (
            .O(N__23039),
            .I(N__23036));
    LocalMux I__2981 (
            .O(N__23036),
            .I(drone_altitude_14));
    InMux I__2980 (
            .O(N__23033),
            .I(N__23030));
    LocalMux I__2979 (
            .O(N__23030),
            .I(\pid_alt.error_axbZ0Z_2 ));
    InMux I__2978 (
            .O(N__23027),
            .I(N__23024));
    LocalMux I__2977 (
            .O(N__23024),
            .I(\pid_alt.error_axbZ0Z_3 ));
    InMux I__2976 (
            .O(N__23021),
            .I(N__23017));
    InMux I__2975 (
            .O(N__23020),
            .I(N__23014));
    LocalMux I__2974 (
            .O(N__23017),
            .I(N__23011));
    LocalMux I__2973 (
            .O(N__23014),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    Odrv12 I__2972 (
            .O(N__23011),
            .I(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ));
    CascadeMux I__2971 (
            .O(N__23006),
            .I(N__23003));
    InMux I__2970 (
            .O(N__23003),
            .I(N__23000));
    LocalMux I__2969 (
            .O(N__23000),
            .I(N__22997));
    Odrv4 I__2968 (
            .O(N__22997),
            .I(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ));
    InMux I__2967 (
            .O(N__22994),
            .I(\pid_alt.un1_pid_prereg_0_cry_13 ));
    InMux I__2966 (
            .O(N__22991),
            .I(N__22988));
    LocalMux I__2965 (
            .O(N__22988),
            .I(N__22985));
    Odrv4 I__2964 (
            .O(N__22985),
            .I(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ));
    CascadeMux I__2963 (
            .O(N__22982),
            .I(N__22978));
    CascadeMux I__2962 (
            .O(N__22981),
            .I(N__22975));
    InMux I__2961 (
            .O(N__22978),
            .I(N__22972));
    InMux I__2960 (
            .O(N__22975),
            .I(N__22969));
    LocalMux I__2959 (
            .O(N__22972),
            .I(N__22966));
    LocalMux I__2958 (
            .O(N__22969),
            .I(N__22963));
    Span4Mux_h I__2957 (
            .O(N__22966),
            .I(N__22958));
    Span4Mux_v I__2956 (
            .O(N__22963),
            .I(N__22958));
    Odrv4 I__2955 (
            .O(N__22958),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ));
    InMux I__2954 (
            .O(N__22955),
            .I(bfn_4_17_0_));
    InMux I__2953 (
            .O(N__22952),
            .I(N__22949));
    LocalMux I__2952 (
            .O(N__22949),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ));
    CascadeMux I__2951 (
            .O(N__22946),
            .I(N__22942));
    InMux I__2950 (
            .O(N__22945),
            .I(N__22939));
    InMux I__2949 (
            .O(N__22942),
            .I(N__22936));
    LocalMux I__2948 (
            .O(N__22939),
            .I(N__22931));
    LocalMux I__2947 (
            .O(N__22936),
            .I(N__22931));
    Span4Mux_v I__2946 (
            .O(N__22931),
            .I(N__22928));
    Odrv4 I__2945 (
            .O(N__22928),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ));
    InMux I__2944 (
            .O(N__22925),
            .I(\pid_alt.un1_pid_prereg_0_cry_15 ));
    InMux I__2943 (
            .O(N__22922),
            .I(N__22919));
    LocalMux I__2942 (
            .O(N__22919),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ));
    CascadeMux I__2941 (
            .O(N__22916),
            .I(N__22912));
    CascadeMux I__2940 (
            .O(N__22915),
            .I(N__22909));
    InMux I__2939 (
            .O(N__22912),
            .I(N__22906));
    InMux I__2938 (
            .O(N__22909),
            .I(N__22903));
    LocalMux I__2937 (
            .O(N__22906),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    LocalMux I__2936 (
            .O(N__22903),
            .I(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ));
    InMux I__2935 (
            .O(N__22898),
            .I(\pid_alt.un1_pid_prereg_0_cry_16 ));
    InMux I__2934 (
            .O(N__22895),
            .I(N__22892));
    LocalMux I__2933 (
            .O(N__22892),
            .I(N__22889));
    Odrv4 I__2932 (
            .O(N__22889),
            .I(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ));
    CascadeMux I__2931 (
            .O(N__22886),
            .I(N__22882));
    InMux I__2930 (
            .O(N__22885),
            .I(N__22879));
    InMux I__2929 (
            .O(N__22882),
            .I(N__22876));
    LocalMux I__2928 (
            .O(N__22879),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    LocalMux I__2927 (
            .O(N__22876),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ));
    InMux I__2926 (
            .O(N__22871),
            .I(\pid_alt.un1_pid_prereg_0_cry_17 ));
    InMux I__2925 (
            .O(N__22868),
            .I(N__22865));
    LocalMux I__2924 (
            .O(N__22865),
            .I(N__22862));
    Odrv4 I__2923 (
            .O(N__22862),
            .I(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ));
    CascadeMux I__2922 (
            .O(N__22859),
            .I(N__22855));
    CascadeMux I__2921 (
            .O(N__22858),
            .I(N__22852));
    InMux I__2920 (
            .O(N__22855),
            .I(N__22849));
    InMux I__2919 (
            .O(N__22852),
            .I(N__22846));
    LocalMux I__2918 (
            .O(N__22849),
            .I(N__22843));
    LocalMux I__2917 (
            .O(N__22846),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    Odrv12 I__2916 (
            .O(N__22843),
            .I(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ));
    InMux I__2915 (
            .O(N__22838),
            .I(\pid_alt.un1_pid_prereg_0_cry_18 ));
    InMux I__2914 (
            .O(N__22835),
            .I(\pid_alt.un1_pid_prereg_0_cry_19 ));
    InMux I__2913 (
            .O(N__22832),
            .I(\pid_alt.un1_pid_prereg_0_cry_20 ));
    InMux I__2912 (
            .O(N__22829),
            .I(\pid_alt.un1_pid_prereg_0_cry_4 ));
    InMux I__2911 (
            .O(N__22826),
            .I(N__22823));
    LocalMux I__2910 (
            .O(N__22823),
            .I(N__22820));
    Span4Mux_h I__2909 (
            .O(N__22820),
            .I(N__22817));
    Odrv4 I__2908 (
            .O(N__22817),
            .I(\pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5 ));
    CascadeMux I__2907 (
            .O(N__22814),
            .I(N__22810));
    CascadeMux I__2906 (
            .O(N__22813),
            .I(N__22807));
    InMux I__2905 (
            .O(N__22810),
            .I(N__22804));
    InMux I__2904 (
            .O(N__22807),
            .I(N__22801));
    LocalMux I__2903 (
            .O(N__22804),
            .I(N__22798));
    LocalMux I__2902 (
            .O(N__22801),
            .I(N__22795));
    Span4Mux_h I__2901 (
            .O(N__22798),
            .I(N__22792));
    Span4Mux_h I__2900 (
            .O(N__22795),
            .I(N__22789));
    Odrv4 I__2899 (
            .O(N__22792),
            .I(\pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4 ));
    Odrv4 I__2898 (
            .O(N__22789),
            .I(\pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4 ));
    InMux I__2897 (
            .O(N__22784),
            .I(\pid_alt.un1_pid_prereg_0_cry_5 ));
    InMux I__2896 (
            .O(N__22781),
            .I(bfn_4_16_0_));
    InMux I__2895 (
            .O(N__22778),
            .I(\pid_alt.un1_pid_prereg_0_cry_7 ));
    InMux I__2894 (
            .O(N__22775),
            .I(N__22772));
    LocalMux I__2893 (
            .O(N__22772),
            .I(N__22769));
    Odrv4 I__2892 (
            .O(N__22769),
            .I(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ));
    InMux I__2891 (
            .O(N__22766),
            .I(\pid_alt.un1_pid_prereg_0_cry_8 ));
    InMux I__2890 (
            .O(N__22763),
            .I(N__22760));
    LocalMux I__2889 (
            .O(N__22760),
            .I(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ));
    CascadeMux I__2888 (
            .O(N__22757),
            .I(N__22754));
    InMux I__2887 (
            .O(N__22754),
            .I(N__22750));
    InMux I__2886 (
            .O(N__22753),
            .I(N__22747));
    LocalMux I__2885 (
            .O(N__22750),
            .I(N__22744));
    LocalMux I__2884 (
            .O(N__22747),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    Odrv4 I__2883 (
            .O(N__22744),
            .I(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ));
    InMux I__2882 (
            .O(N__22739),
            .I(\pid_alt.un1_pid_prereg_0_cry_9 ));
    InMux I__2881 (
            .O(N__22736),
            .I(\pid_alt.un1_pid_prereg_0_cry_10 ));
    InMux I__2880 (
            .O(N__22733),
            .I(N__22730));
    LocalMux I__2879 (
            .O(N__22730),
            .I(N__22727));
    Odrv12 I__2878 (
            .O(N__22727),
            .I(\pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11 ));
    InMux I__2877 (
            .O(N__22724),
            .I(\pid_alt.un1_pid_prereg_0_cry_11 ));
    InMux I__2876 (
            .O(N__22721),
            .I(N__22718));
    LocalMux I__2875 (
            .O(N__22718),
            .I(N__22715));
    Odrv12 I__2874 (
            .O(N__22715),
            .I(\pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12 ));
    CascadeMux I__2873 (
            .O(N__22712),
            .I(N__22709));
    InMux I__2872 (
            .O(N__22709),
            .I(N__22705));
    CascadeMux I__2871 (
            .O(N__22708),
            .I(N__22702));
    LocalMux I__2870 (
            .O(N__22705),
            .I(N__22699));
    InMux I__2869 (
            .O(N__22702),
            .I(N__22696));
    Span4Mux_v I__2868 (
            .O(N__22699),
            .I(N__22693));
    LocalMux I__2867 (
            .O(N__22696),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11 ));
    Odrv4 I__2866 (
            .O(N__22693),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11 ));
    InMux I__2865 (
            .O(N__22688),
            .I(\pid_alt.un1_pid_prereg_0_cry_12 ));
    CascadeMux I__2864 (
            .O(N__22685),
            .I(\pid_alt.N_294_cascade_ ));
    CascadeMux I__2863 (
            .O(N__22682),
            .I(N__22677));
    InMux I__2862 (
            .O(N__22681),
            .I(N__22667));
    InMux I__2861 (
            .O(N__22680),
            .I(N__22667));
    InMux I__2860 (
            .O(N__22677),
            .I(N__22667));
    InMux I__2859 (
            .O(N__22676),
            .I(N__22667));
    LocalMux I__2858 (
            .O(N__22667),
            .I(\pid_alt.N_294 ));
    CascadeMux I__2857 (
            .O(N__22664),
            .I(N__22661));
    InMux I__2856 (
            .O(N__22661),
            .I(N__22655));
    InMux I__2855 (
            .O(N__22660),
            .I(N__22655));
    LocalMux I__2854 (
            .O(N__22655),
            .I(N__22652));
    Span4Mux_v I__2853 (
            .O(N__22652),
            .I(N__22644));
    InMux I__2852 (
            .O(N__22651),
            .I(N__22635));
    InMux I__2851 (
            .O(N__22650),
            .I(N__22635));
    InMux I__2850 (
            .O(N__22649),
            .I(N__22635));
    InMux I__2849 (
            .O(N__22648),
            .I(N__22635));
    CascadeMux I__2848 (
            .O(N__22647),
            .I(N__22632));
    Span4Mux_v I__2847 (
            .O(N__22644),
            .I(N__22625));
    LocalMux I__2846 (
            .O(N__22635),
            .I(N__22622));
    InMux I__2845 (
            .O(N__22632),
            .I(N__22611));
    InMux I__2844 (
            .O(N__22631),
            .I(N__22611));
    InMux I__2843 (
            .O(N__22630),
            .I(N__22611));
    InMux I__2842 (
            .O(N__22629),
            .I(N__22611));
    InMux I__2841 (
            .O(N__22628),
            .I(N__22611));
    Odrv4 I__2840 (
            .O(N__22625),
            .I(\pid_alt.N_295 ));
    Odrv4 I__2839 (
            .O(N__22622),
            .I(\pid_alt.N_295 ));
    LocalMux I__2838 (
            .O(N__22611),
            .I(\pid_alt.N_295 ));
    InMux I__2837 (
            .O(N__22604),
            .I(N__22600));
    InMux I__2836 (
            .O(N__22603),
            .I(N__22597));
    LocalMux I__2835 (
            .O(N__22600),
            .I(N__22591));
    LocalMux I__2834 (
            .O(N__22597),
            .I(N__22591));
    InMux I__2833 (
            .O(N__22596),
            .I(N__22588));
    Odrv4 I__2832 (
            .O(N__22591),
            .I(\pid_alt.error_i_acumm7lto4 ));
    LocalMux I__2831 (
            .O(N__22588),
            .I(\pid_alt.error_i_acumm7lto4 ));
    InMux I__2830 (
            .O(N__22583),
            .I(N__22580));
    LocalMux I__2829 (
            .O(N__22580),
            .I(\pid_alt.error_i_acummZ0Z_4 ));
    InMux I__2828 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__2827 (
            .O(N__22574),
            .I(N__22571));
    Span4Mux_v I__2826 (
            .O(N__22571),
            .I(N__22568));
    Span4Mux_s2_h I__2825 (
            .O(N__22568),
            .I(N__22564));
    InMux I__2824 (
            .O(N__22567),
            .I(N__22561));
    Odrv4 I__2823 (
            .O(N__22564),
            .I(\pid_alt.un1_pid_prereg_0 ));
    LocalMux I__2822 (
            .O(N__22561),
            .I(\pid_alt.un1_pid_prereg_0 ));
    CascadeMux I__2821 (
            .O(N__22556),
            .I(N__22553));
    InMux I__2820 (
            .O(N__22553),
            .I(N__22550));
    LocalMux I__2819 (
            .O(N__22550),
            .I(N__22547));
    Span4Mux_v I__2818 (
            .O(N__22547),
            .I(N__22544));
    Odrv4 I__2817 (
            .O(N__22544),
            .I(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ));
    InMux I__2816 (
            .O(N__22541),
            .I(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ));
    InMux I__2815 (
            .O(N__22538),
            .I(N__22535));
    LocalMux I__2814 (
            .O(N__22535),
            .I(N__22532));
    Span4Mux_v I__2813 (
            .O(N__22532),
            .I(N__22529));
    Odrv4 I__2812 (
            .O(N__22529),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ));
    InMux I__2811 (
            .O(N__22526),
            .I(\pid_alt.un1_pid_prereg_0_cry_0 ));
    InMux I__2810 (
            .O(N__22523),
            .I(N__22520));
    LocalMux I__2809 (
            .O(N__22520),
            .I(N__22517));
    Span4Mux_h I__2808 (
            .O(N__22517),
            .I(N__22514));
    Odrv4 I__2807 (
            .O(N__22514),
            .I(\pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ));
    InMux I__2806 (
            .O(N__22511),
            .I(\pid_alt.un1_pid_prereg_0_cry_1 ));
    InMux I__2805 (
            .O(N__22508),
            .I(N__22505));
    LocalMux I__2804 (
            .O(N__22505),
            .I(N__22502));
    Span4Mux_h I__2803 (
            .O(N__22502),
            .I(N__22499));
    Odrv4 I__2802 (
            .O(N__22499),
            .I(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ));
    InMux I__2801 (
            .O(N__22496),
            .I(\pid_alt.un1_pid_prereg_0_cry_2 ));
    CascadeMux I__2800 (
            .O(N__22493),
            .I(N__22490));
    InMux I__2799 (
            .O(N__22490),
            .I(N__22486));
    InMux I__2798 (
            .O(N__22489),
            .I(N__22483));
    LocalMux I__2797 (
            .O(N__22486),
            .I(N__22478));
    LocalMux I__2796 (
            .O(N__22483),
            .I(N__22478));
    Span4Mux_h I__2795 (
            .O(N__22478),
            .I(N__22475));
    Odrv4 I__2794 (
            .O(N__22475),
            .I(\pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ));
    CascadeMux I__2793 (
            .O(N__22472),
            .I(N__22469));
    InMux I__2792 (
            .O(N__22469),
            .I(N__22466));
    LocalMux I__2791 (
            .O(N__22466),
            .I(N__22463));
    Odrv4 I__2790 (
            .O(N__22463),
            .I(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ));
    InMux I__2789 (
            .O(N__22460),
            .I(\pid_alt.un1_pid_prereg_0_cry_3 ));
    InMux I__2788 (
            .O(N__22457),
            .I(N__22454));
    LocalMux I__2787 (
            .O(N__22454),
            .I(N__22451));
    Odrv4 I__2786 (
            .O(N__22451),
            .I(\pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4 ));
    CascadeMux I__2785 (
            .O(N__22448),
            .I(N__22444));
    InMux I__2784 (
            .O(N__22447),
            .I(N__22441));
    InMux I__2783 (
            .O(N__22444),
            .I(N__22438));
    LocalMux I__2782 (
            .O(N__22441),
            .I(N__22433));
    LocalMux I__2781 (
            .O(N__22438),
            .I(N__22433));
    Odrv4 I__2780 (
            .O(N__22433),
            .I(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ));
    CascadeMux I__2779 (
            .O(N__22430),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ));
    InMux I__2778 (
            .O(N__22427),
            .I(N__22418));
    InMux I__2777 (
            .O(N__22426),
            .I(N__22418));
    InMux I__2776 (
            .O(N__22425),
            .I(N__22418));
    LocalMux I__2775 (
            .O(N__22418),
            .I(N__22415));
    Span4Mux_h I__2774 (
            .O(N__22415),
            .I(N__22412));
    Span4Mux_v I__2773 (
            .O(N__22412),
            .I(N__22409));
    Odrv4 I__2772 (
            .O(N__22409),
            .I(\pid_alt.error_d_regZ0Z_14 ));
    CascadeMux I__2771 (
            .O(N__22406),
            .I(N__22403));
    InMux I__2770 (
            .O(N__22403),
            .I(N__22397));
    InMux I__2769 (
            .O(N__22402),
            .I(N__22397));
    LocalMux I__2768 (
            .O(N__22397),
            .I(\pid_alt.error_d_reg_prevZ0Z_14 ));
    InMux I__2767 (
            .O(N__22394),
            .I(N__22388));
    InMux I__2766 (
            .O(N__22393),
            .I(N__22388));
    LocalMux I__2765 (
            .O(N__22388),
            .I(N__22385));
    Span4Mux_h I__2764 (
            .O(N__22385),
            .I(N__22382));
    Odrv4 I__2763 (
            .O(N__22382),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ));
    InMux I__2762 (
            .O(N__22379),
            .I(N__22376));
    LocalMux I__2761 (
            .O(N__22376),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ));
    CascadeMux I__2760 (
            .O(N__22373),
            .I(N__22370));
    InMux I__2759 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__2758 (
            .O(N__22367),
            .I(\pid_alt.error_i_acummZ0Z_5 ));
    CascadeMux I__2757 (
            .O(N__22364),
            .I(\pid_alt.N_295_cascade_ ));
    InMux I__2756 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__2755 (
            .O(N__22358),
            .I(\pid_alt.error_i_acummZ0Z_1 ));
    InMux I__2754 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__2753 (
            .O(N__22352),
            .I(\pid_alt.error_i_acummZ0Z_2 ));
    InMux I__2752 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__2751 (
            .O(N__22346),
            .I(\pid_alt.error_i_acummZ0Z_3 ));
    CascadeMux I__2750 (
            .O(N__22343),
            .I(N__22340));
    InMux I__2749 (
            .O(N__22340),
            .I(N__22334));
    InMux I__2748 (
            .O(N__22339),
            .I(N__22334));
    LocalMux I__2747 (
            .O(N__22334),
            .I(\pid_alt.m39_i_a2_3 ));
    CascadeMux I__2746 (
            .O(N__22331),
            .I(N__22327));
    InMux I__2745 (
            .O(N__22330),
            .I(N__22322));
    InMux I__2744 (
            .O(N__22327),
            .I(N__22322));
    LocalMux I__2743 (
            .O(N__22322),
            .I(N__22319));
    Odrv4 I__2742 (
            .O(N__22319),
            .I(\pid_alt.m39_i_a2_4 ));
    InMux I__2741 (
            .O(N__22316),
            .I(N__22309));
    InMux I__2740 (
            .O(N__22315),
            .I(N__22309));
    InMux I__2739 (
            .O(N__22314),
            .I(N__22306));
    LocalMux I__2738 (
            .O(N__22309),
            .I(\pid_alt.error_i_acumm7lto5 ));
    LocalMux I__2737 (
            .O(N__22306),
            .I(\pid_alt.error_i_acumm7lto5 ));
    InMux I__2736 (
            .O(N__22301),
            .I(N__22297));
    InMux I__2735 (
            .O(N__22300),
            .I(N__22294));
    LocalMux I__2734 (
            .O(N__22297),
            .I(N__22291));
    LocalMux I__2733 (
            .O(N__22294),
            .I(N__22288));
    Span12Mux_v I__2732 (
            .O(N__22291),
            .I(N__22285));
    Span12Mux_v I__2731 (
            .O(N__22288),
            .I(N__22282));
    Odrv12 I__2730 (
            .O(N__22285),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    Odrv12 I__2729 (
            .O(N__22282),
            .I(\pid_alt.error_p_regZ0Z_13 ));
    InMux I__2728 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__2727 (
            .O(N__22274),
            .I(N__22270));
    InMux I__2726 (
            .O(N__22273),
            .I(N__22267));
    Span4Mux_h I__2725 (
            .O(N__22270),
            .I(N__22264));
    LocalMux I__2724 (
            .O(N__22267),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    Odrv4 I__2723 (
            .O(N__22264),
            .I(\pid_alt.error_d_reg_prevZ0Z_13 ));
    InMux I__2722 (
            .O(N__22259),
            .I(N__22254));
    InMux I__2721 (
            .O(N__22258),
            .I(N__22251));
    InMux I__2720 (
            .O(N__22257),
            .I(N__22248));
    LocalMux I__2719 (
            .O(N__22254),
            .I(N__22243));
    LocalMux I__2718 (
            .O(N__22251),
            .I(N__22243));
    LocalMux I__2717 (
            .O(N__22248),
            .I(N__22240));
    Span4Mux_v I__2716 (
            .O(N__22243),
            .I(N__22235));
    Span4Mux_h I__2715 (
            .O(N__22240),
            .I(N__22235));
    Span4Mux_v I__2714 (
            .O(N__22235),
            .I(N__22232));
    Odrv4 I__2713 (
            .O(N__22232),
            .I(\pid_alt.error_d_regZ0Z_13 ));
    InMux I__2712 (
            .O(N__22229),
            .I(N__22223));
    InMux I__2711 (
            .O(N__22228),
            .I(N__22223));
    LocalMux I__2710 (
            .O(N__22223),
            .I(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ));
    InMux I__2709 (
            .O(N__22220),
            .I(N__22214));
    InMux I__2708 (
            .O(N__22219),
            .I(N__22214));
    LocalMux I__2707 (
            .O(N__22214),
            .I(N__22211));
    Span4Mux_h I__2706 (
            .O(N__22211),
            .I(N__22208));
    Span4Mux_v I__2705 (
            .O(N__22208),
            .I(N__22205));
    Span4Mux_v I__2704 (
            .O(N__22205),
            .I(N__22202));
    Odrv4 I__2703 (
            .O(N__22202),
            .I(\pid_alt.error_p_regZ0Z_12 ));
    InMux I__2702 (
            .O(N__22199),
            .I(N__22196));
    LocalMux I__2701 (
            .O(N__22196),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ));
    CascadeMux I__2700 (
            .O(N__22193),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ));
    InMux I__2699 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__2698 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__2697 (
            .O(N__22184),
            .I(N__22181));
    Odrv4 I__2696 (
            .O(N__22181),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ));
    CascadeMux I__2695 (
            .O(N__22178),
            .I(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ));
    InMux I__2694 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__2693 (
            .O(N__22172),
            .I(N__22168));
    InMux I__2692 (
            .O(N__22171),
            .I(N__22165));
    Span4Mux_h I__2691 (
            .O(N__22168),
            .I(N__22162));
    LocalMux I__2690 (
            .O(N__22165),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    Odrv4 I__2689 (
            .O(N__22162),
            .I(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ));
    InMux I__2688 (
            .O(N__22157),
            .I(N__22151));
    InMux I__2687 (
            .O(N__22156),
            .I(N__22151));
    LocalMux I__2686 (
            .O(N__22151),
            .I(N__22148));
    Span4Mux_h I__2685 (
            .O(N__22148),
            .I(N__22145));
    Span4Mux_v I__2684 (
            .O(N__22145),
            .I(N__22142));
    Span4Mux_v I__2683 (
            .O(N__22142),
            .I(N__22139));
    Odrv4 I__2682 (
            .O(N__22139),
            .I(\pid_alt.error_p_regZ0Z_14 ));
    CascadeMux I__2681 (
            .O(N__22136),
            .I(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ));
    CascadeMux I__2680 (
            .O(N__22133),
            .I(N__22130));
    InMux I__2679 (
            .O(N__22130),
            .I(N__22127));
    LocalMux I__2678 (
            .O(N__22127),
            .I(\Commands_frame_decoder.state_ns_0_a3_3_1 ));
    InMux I__2677 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__2676 (
            .O(N__22121),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ));
    CascadeMux I__2675 (
            .O(N__22118),
            .I(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ));
    InMux I__2674 (
            .O(N__22115),
            .I(N__22108));
    InMux I__2673 (
            .O(N__22114),
            .I(N__22108));
    InMux I__2672 (
            .O(N__22113),
            .I(N__22105));
    LocalMux I__2671 (
            .O(N__22108),
            .I(N__22102));
    LocalMux I__2670 (
            .O(N__22105),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    Odrv4 I__2669 (
            .O(N__22102),
            .I(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ));
    InMux I__2668 (
            .O(N__22097),
            .I(N__22094));
    LocalMux I__2667 (
            .O(N__22094),
            .I(N__22091));
    Span4Mux_v I__2666 (
            .O(N__22091),
            .I(N__22086));
    InMux I__2665 (
            .O(N__22090),
            .I(N__22083));
    InMux I__2664 (
            .O(N__22089),
            .I(N__22080));
    Span4Mux_v I__2663 (
            .O(N__22086),
            .I(N__22077));
    LocalMux I__2662 (
            .O(N__22083),
            .I(N__22074));
    LocalMux I__2661 (
            .O(N__22080),
            .I(N__22071));
    Sp12to4 I__2660 (
            .O(N__22077),
            .I(N__22068));
    Span4Mux_s3_h I__2659 (
            .O(N__22074),
            .I(N__22065));
    Span4Mux_s3_h I__2658 (
            .O(N__22071),
            .I(N__22062));
    Span12Mux_s3_h I__2657 (
            .O(N__22068),
            .I(N__22057));
    Sp12to4 I__2656 (
            .O(N__22065),
            .I(N__22057));
    Span4Mux_v I__2655 (
            .O(N__22062),
            .I(N__22054));
    Odrv12 I__2654 (
            .O(N__22057),
            .I(\pid_alt.error_14 ));
    Odrv4 I__2653 (
            .O(N__22054),
            .I(\pid_alt.error_14 ));
    InMux I__2652 (
            .O(N__22049),
            .I(\pid_alt.error_cry_13 ));
    InMux I__2651 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__2650 (
            .O(N__22043),
            .I(drone_altitude_15));
    InMux I__2649 (
            .O(N__22040),
            .I(\pid_alt.error_cry_14 ));
    InMux I__2648 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__2647 (
            .O(N__22034),
            .I(N__22029));
    InMux I__2646 (
            .O(N__22033),
            .I(N__22026));
    InMux I__2645 (
            .O(N__22032),
            .I(N__22023));
    Span12Mux_s7_v I__2644 (
            .O(N__22029),
            .I(N__22018));
    LocalMux I__2643 (
            .O(N__22026),
            .I(N__22018));
    LocalMux I__2642 (
            .O(N__22023),
            .I(N__22015));
    Span12Mux_v I__2641 (
            .O(N__22018),
            .I(N__22010));
    Span12Mux_s10_v I__2640 (
            .O(N__22015),
            .I(N__22010));
    Odrv12 I__2639 (
            .O(N__22010),
            .I(\pid_alt.error_15 ));
    InMux I__2638 (
            .O(N__22007),
            .I(N__22004));
    LocalMux I__2637 (
            .O(N__22004),
            .I(\dron_frame_decoder_1.drone_altitude_11 ));
    InMux I__2636 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__2635 (
            .O(N__21998),
            .I(drone_altitude_i_11));
    CascadeMux I__2634 (
            .O(N__21995),
            .I(N__21991));
    InMux I__2633 (
            .O(N__21994),
            .I(N__21988));
    InMux I__2632 (
            .O(N__21991),
            .I(N__21985));
    LocalMux I__2631 (
            .O(N__21988),
            .I(N__21982));
    LocalMux I__2630 (
            .O(N__21985),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    Odrv12 I__2629 (
            .O(N__21982),
            .I(\pid_alt.error_i_acummZ0Z_11 ));
    InMux I__2628 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__2627 (
            .O(N__21974),
            .I(N__21971));
    Span4Mux_h I__2626 (
            .O(N__21971),
            .I(N__21967));
    InMux I__2625 (
            .O(N__21970),
            .I(N__21964));
    Span4Mux_v I__2624 (
            .O(N__21967),
            .I(N__21961));
    LocalMux I__2623 (
            .O(N__21964),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    Odrv4 I__2622 (
            .O(N__21961),
            .I(\pid_alt.error_i_acummZ0Z_7 ));
    InMux I__2621 (
            .O(N__21956),
            .I(N__21953));
    LocalMux I__2620 (
            .O(N__21953),
            .I(N__21950));
    Span4Mux_s3_h I__2619 (
            .O(N__21950),
            .I(N__21947));
    Odrv4 I__2618 (
            .O(N__21947),
            .I(alt_kp_1));
    InMux I__2617 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__2616 (
            .O(N__21941),
            .I(N__21938));
    Span4Mux_s3_h I__2615 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__2614 (
            .O(N__21935),
            .I(alt_kp_7));
    CEMux I__2613 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2612 (
            .O(N__21929),
            .I(N__21924));
    CEMux I__2611 (
            .O(N__21928),
            .I(N__21921));
    CEMux I__2610 (
            .O(N__21927),
            .I(N__21918));
    Span4Mux_h I__2609 (
            .O(N__21924),
            .I(N__21915));
    LocalMux I__2608 (
            .O(N__21921),
            .I(N__21912));
    LocalMux I__2607 (
            .O(N__21918),
            .I(N__21909));
    Odrv4 I__2606 (
            .O(N__21915),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    Odrv4 I__2605 (
            .O(N__21912),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    Odrv12 I__2604 (
            .O(N__21909),
            .I(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ));
    CascadeMux I__2603 (
            .O(N__21902),
            .I(N__21898));
    CascadeMux I__2602 (
            .O(N__21901),
            .I(N__21895));
    InMux I__2601 (
            .O(N__21898),
            .I(N__21892));
    InMux I__2600 (
            .O(N__21895),
            .I(N__21889));
    LocalMux I__2599 (
            .O(N__21892),
            .I(alt_command_2));
    LocalMux I__2598 (
            .O(N__21889),
            .I(alt_command_2));
    InMux I__2597 (
            .O(N__21884),
            .I(N__21880));
    InMux I__2596 (
            .O(N__21883),
            .I(N__21877));
    LocalMux I__2595 (
            .O(N__21880),
            .I(N__21874));
    LocalMux I__2594 (
            .O(N__21877),
            .I(N__21870));
    Span4Mux_s3_h I__2593 (
            .O(N__21874),
            .I(N__21867));
    InMux I__2592 (
            .O(N__21873),
            .I(N__21864));
    Span4Mux_s3_h I__2591 (
            .O(N__21870),
            .I(N__21861));
    Span4Mux_v I__2590 (
            .O(N__21867),
            .I(N__21858));
    LocalMux I__2589 (
            .O(N__21864),
            .I(N__21855));
    Span4Mux_v I__2588 (
            .O(N__21861),
            .I(N__21852));
    Sp12to4 I__2587 (
            .O(N__21858),
            .I(N__21847));
    Span12Mux_s3_h I__2586 (
            .O(N__21855),
            .I(N__21847));
    Odrv4 I__2585 (
            .O(N__21852),
            .I(\pid_alt.error_6 ));
    Odrv12 I__2584 (
            .O(N__21847),
            .I(\pid_alt.error_6 ));
    InMux I__2583 (
            .O(N__21842),
            .I(\pid_alt.error_cry_5 ));
    InMux I__2582 (
            .O(N__21839),
            .I(N__21836));
    LocalMux I__2581 (
            .O(N__21836),
            .I(drone_altitude_i_7));
    CascadeMux I__2580 (
            .O(N__21833),
            .I(N__21829));
    CascadeMux I__2579 (
            .O(N__21832),
            .I(N__21826));
    InMux I__2578 (
            .O(N__21829),
            .I(N__21823));
    InMux I__2577 (
            .O(N__21826),
            .I(N__21820));
    LocalMux I__2576 (
            .O(N__21823),
            .I(alt_command_3));
    LocalMux I__2575 (
            .O(N__21820),
            .I(alt_command_3));
    InMux I__2574 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__2573 (
            .O(N__21812),
            .I(N__21807));
    InMux I__2572 (
            .O(N__21811),
            .I(N__21804));
    InMux I__2571 (
            .O(N__21810),
            .I(N__21801));
    Span12Mux_s6_v I__2570 (
            .O(N__21807),
            .I(N__21796));
    LocalMux I__2569 (
            .O(N__21804),
            .I(N__21796));
    LocalMux I__2568 (
            .O(N__21801),
            .I(N__21793));
    Span12Mux_v I__2567 (
            .O(N__21796),
            .I(N__21788));
    Span12Mux_s11_v I__2566 (
            .O(N__21793),
            .I(N__21788));
    Odrv12 I__2565 (
            .O(N__21788),
            .I(\pid_alt.error_7 ));
    InMux I__2564 (
            .O(N__21785),
            .I(\pid_alt.error_cry_6 ));
    InMux I__2563 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__2562 (
            .O(N__21779),
            .I(drone_altitude_i_8));
    CascadeMux I__2561 (
            .O(N__21776),
            .I(N__21773));
    InMux I__2560 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__2559 (
            .O(N__21770),
            .I(alt_command_4));
    InMux I__2558 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__2557 (
            .O(N__21764),
            .I(N__21760));
    InMux I__2556 (
            .O(N__21763),
            .I(N__21756));
    Span4Mux_v I__2555 (
            .O(N__21760),
            .I(N__21753));
    InMux I__2554 (
            .O(N__21759),
            .I(N__21750));
    LocalMux I__2553 (
            .O(N__21756),
            .I(N__21747));
    Span4Mux_v I__2552 (
            .O(N__21753),
            .I(N__21744));
    LocalMux I__2551 (
            .O(N__21750),
            .I(N__21741));
    Span4Mux_s3_h I__2550 (
            .O(N__21747),
            .I(N__21738));
    Span4Mux_v I__2549 (
            .O(N__21744),
            .I(N__21735));
    Span4Mux_v I__2548 (
            .O(N__21741),
            .I(N__21732));
    Span4Mux_v I__2547 (
            .O(N__21738),
            .I(N__21729));
    Span4Mux_h I__2546 (
            .O(N__21735),
            .I(N__21724));
    Span4Mux_h I__2545 (
            .O(N__21732),
            .I(N__21724));
    Odrv4 I__2544 (
            .O(N__21729),
            .I(\pid_alt.error_8 ));
    Odrv4 I__2543 (
            .O(N__21724),
            .I(\pid_alt.error_8 ));
    InMux I__2542 (
            .O(N__21719),
            .I(bfn_3_20_0_));
    InMux I__2541 (
            .O(N__21716),
            .I(N__21713));
    LocalMux I__2540 (
            .O(N__21713),
            .I(drone_altitude_i_9));
    CascadeMux I__2539 (
            .O(N__21710),
            .I(N__21707));
    InMux I__2538 (
            .O(N__21707),
            .I(N__21704));
    LocalMux I__2537 (
            .O(N__21704),
            .I(alt_command_5));
    InMux I__2536 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__2535 (
            .O(N__21698),
            .I(N__21693));
    InMux I__2534 (
            .O(N__21697),
            .I(N__21690));
    InMux I__2533 (
            .O(N__21696),
            .I(N__21687));
    Span4Mux_v I__2532 (
            .O(N__21693),
            .I(N__21684));
    LocalMux I__2531 (
            .O(N__21690),
            .I(N__21681));
    LocalMux I__2530 (
            .O(N__21687),
            .I(N__21678));
    Sp12to4 I__2529 (
            .O(N__21684),
            .I(N__21675));
    Span4Mux_s3_h I__2528 (
            .O(N__21681),
            .I(N__21672));
    Span4Mux_s3_h I__2527 (
            .O(N__21678),
            .I(N__21669));
    Span12Mux_s3_h I__2526 (
            .O(N__21675),
            .I(N__21666));
    Span4Mux_v I__2525 (
            .O(N__21672),
            .I(N__21663));
    Span4Mux_v I__2524 (
            .O(N__21669),
            .I(N__21660));
    Odrv12 I__2523 (
            .O(N__21666),
            .I(\pid_alt.error_9 ));
    Odrv4 I__2522 (
            .O(N__21663),
            .I(\pid_alt.error_9 ));
    Odrv4 I__2521 (
            .O(N__21660),
            .I(\pid_alt.error_9 ));
    InMux I__2520 (
            .O(N__21653),
            .I(\pid_alt.error_cry_8 ));
    InMux I__2519 (
            .O(N__21650),
            .I(N__21647));
    LocalMux I__2518 (
            .O(N__21647),
            .I(drone_altitude_i_10));
    CascadeMux I__2517 (
            .O(N__21644),
            .I(N__21641));
    InMux I__2516 (
            .O(N__21641),
            .I(N__21638));
    LocalMux I__2515 (
            .O(N__21638),
            .I(alt_command_6));
    InMux I__2514 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__2513 (
            .O(N__21632),
            .I(N__21627));
    InMux I__2512 (
            .O(N__21631),
            .I(N__21624));
    InMux I__2511 (
            .O(N__21630),
            .I(N__21621));
    Span4Mux_v I__2510 (
            .O(N__21627),
            .I(N__21618));
    LocalMux I__2509 (
            .O(N__21624),
            .I(N__21615));
    LocalMux I__2508 (
            .O(N__21621),
            .I(N__21612));
    Sp12to4 I__2507 (
            .O(N__21618),
            .I(N__21609));
    Span4Mux_s3_h I__2506 (
            .O(N__21615),
            .I(N__21606));
    Span4Mux_s3_h I__2505 (
            .O(N__21612),
            .I(N__21603));
    Span12Mux_s3_h I__2504 (
            .O(N__21609),
            .I(N__21600));
    Span4Mux_v I__2503 (
            .O(N__21606),
            .I(N__21597));
    Span4Mux_v I__2502 (
            .O(N__21603),
            .I(N__21594));
    Odrv12 I__2501 (
            .O(N__21600),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2500 (
            .O(N__21597),
            .I(\pid_alt.error_10 ));
    Odrv4 I__2499 (
            .O(N__21594),
            .I(\pid_alt.error_10 ));
    InMux I__2498 (
            .O(N__21587),
            .I(\pid_alt.error_cry_9 ));
    CascadeMux I__2497 (
            .O(N__21584),
            .I(N__21581));
    InMux I__2496 (
            .O(N__21581),
            .I(N__21578));
    LocalMux I__2495 (
            .O(N__21578),
            .I(alt_command_7));
    InMux I__2494 (
            .O(N__21575),
            .I(N__21570));
    InMux I__2493 (
            .O(N__21574),
            .I(N__21567));
    InMux I__2492 (
            .O(N__21573),
            .I(N__21564));
    LocalMux I__2491 (
            .O(N__21570),
            .I(N__21561));
    LocalMux I__2490 (
            .O(N__21567),
            .I(N__21558));
    LocalMux I__2489 (
            .O(N__21564),
            .I(N__21555));
    Span12Mux_s3_h I__2488 (
            .O(N__21561),
            .I(N__21552));
    Span4Mux_s3_h I__2487 (
            .O(N__21558),
            .I(N__21549));
    Span4Mux_s3_h I__2486 (
            .O(N__21555),
            .I(N__21546));
    Span12Mux_v I__2485 (
            .O(N__21552),
            .I(N__21543));
    Span4Mux_v I__2484 (
            .O(N__21549),
            .I(N__21540));
    Span4Mux_v I__2483 (
            .O(N__21546),
            .I(N__21537));
    Odrv12 I__2482 (
            .O(N__21543),
            .I(\pid_alt.error_11 ));
    Odrv4 I__2481 (
            .O(N__21540),
            .I(\pid_alt.error_11 ));
    Odrv4 I__2480 (
            .O(N__21537),
            .I(\pid_alt.error_11 ));
    InMux I__2479 (
            .O(N__21530),
            .I(\pid_alt.error_cry_10 ));
    InMux I__2478 (
            .O(N__21527),
            .I(N__21524));
    LocalMux I__2477 (
            .O(N__21524),
            .I(N__21521));
    Span4Mux_h I__2476 (
            .O(N__21521),
            .I(N__21516));
    InMux I__2475 (
            .O(N__21520),
            .I(N__21513));
    InMux I__2474 (
            .O(N__21519),
            .I(N__21510));
    Span4Mux_v I__2473 (
            .O(N__21516),
            .I(N__21507));
    LocalMux I__2472 (
            .O(N__21513),
            .I(N__21504));
    LocalMux I__2471 (
            .O(N__21510),
            .I(N__21501));
    Span4Mux_v I__2470 (
            .O(N__21507),
            .I(N__21498));
    Span4Mux_v I__2469 (
            .O(N__21504),
            .I(N__21495));
    Span12Mux_s3_h I__2468 (
            .O(N__21501),
            .I(N__21492));
    Span4Mux_v I__2467 (
            .O(N__21498),
            .I(N__21487));
    Span4Mux_h I__2466 (
            .O(N__21495),
            .I(N__21487));
    Odrv12 I__2465 (
            .O(N__21492),
            .I(\pid_alt.error_12 ));
    Odrv4 I__2464 (
            .O(N__21487),
            .I(\pid_alt.error_12 ));
    InMux I__2463 (
            .O(N__21482),
            .I(\pid_alt.error_cry_11 ));
    InMux I__2462 (
            .O(N__21479),
            .I(N__21476));
    LocalMux I__2461 (
            .O(N__21476),
            .I(N__21472));
    InMux I__2460 (
            .O(N__21475),
            .I(N__21469));
    Span4Mux_s2_h I__2459 (
            .O(N__21472),
            .I(N__21465));
    LocalMux I__2458 (
            .O(N__21469),
            .I(N__21462));
    InMux I__2457 (
            .O(N__21468),
            .I(N__21459));
    Sp12to4 I__2456 (
            .O(N__21465),
            .I(N__21456));
    Span4Mux_s3_h I__2455 (
            .O(N__21462),
            .I(N__21453));
    LocalMux I__2454 (
            .O(N__21459),
            .I(N__21450));
    Span12Mux_v I__2453 (
            .O(N__21456),
            .I(N__21447));
    Span4Mux_v I__2452 (
            .O(N__21453),
            .I(N__21444));
    Span12Mux_s3_h I__2451 (
            .O(N__21450),
            .I(N__21441));
    Odrv12 I__2450 (
            .O(N__21447),
            .I(\pid_alt.error_13 ));
    Odrv4 I__2449 (
            .O(N__21444),
            .I(\pid_alt.error_13 ));
    Odrv12 I__2448 (
            .O(N__21441),
            .I(\pid_alt.error_13 ));
    InMux I__2447 (
            .O(N__21434),
            .I(\pid_alt.error_cry_12 ));
    InMux I__2446 (
            .O(N__21431),
            .I(N__21422));
    InMux I__2445 (
            .O(N__21430),
            .I(N__21422));
    InMux I__2444 (
            .O(N__21429),
            .I(N__21422));
    LocalMux I__2443 (
            .O(N__21422),
            .I(\Commands_frame_decoder.source_CH1data8 ));
    InMux I__2442 (
            .O(N__21419),
            .I(N__21416));
    LocalMux I__2441 (
            .O(N__21416),
            .I(N__21413));
    Span4Mux_v I__2440 (
            .O(N__21413),
            .I(N__21409));
    InMux I__2439 (
            .O(N__21412),
            .I(N__21406));
    Span4Mux_v I__2438 (
            .O(N__21409),
            .I(N__21403));
    LocalMux I__2437 (
            .O(N__21406),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ));
    Odrv4 I__2436 (
            .O(N__21403),
            .I(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ));
    InMux I__2435 (
            .O(N__21398),
            .I(N__21393));
    InMux I__2434 (
            .O(N__21397),
            .I(N__21390));
    InMux I__2433 (
            .O(N__21396),
            .I(N__21387));
    LocalMux I__2432 (
            .O(N__21393),
            .I(N__21384));
    LocalMux I__2431 (
            .O(N__21390),
            .I(N__21381));
    LocalMux I__2430 (
            .O(N__21387),
            .I(N__21378));
    Span4Mux_s3_h I__2429 (
            .O(N__21384),
            .I(N__21375));
    Span4Mux_v I__2428 (
            .O(N__21381),
            .I(N__21372));
    Span4Mux_s3_h I__2427 (
            .O(N__21378),
            .I(N__21369));
    Sp12to4 I__2426 (
            .O(N__21375),
            .I(N__21366));
    Span4Mux_h I__2425 (
            .O(N__21372),
            .I(N__21363));
    Span4Mux_v I__2424 (
            .O(N__21369),
            .I(N__21360));
    Odrv12 I__2423 (
            .O(N__21366),
            .I(\pid_alt.error_1 ));
    Odrv4 I__2422 (
            .O(N__21363),
            .I(\pid_alt.error_1 ));
    Odrv4 I__2421 (
            .O(N__21360),
            .I(\pid_alt.error_1 ));
    InMux I__2420 (
            .O(N__21353),
            .I(\pid_alt.error_cry_0 ));
    InMux I__2419 (
            .O(N__21350),
            .I(N__21347));
    LocalMux I__2418 (
            .O(N__21347),
            .I(N__21344));
    Span4Mux_h I__2417 (
            .O(N__21344),
            .I(N__21339));
    InMux I__2416 (
            .O(N__21343),
            .I(N__21336));
    InMux I__2415 (
            .O(N__21342),
            .I(N__21333));
    Span4Mux_v I__2414 (
            .O(N__21339),
            .I(N__21328));
    LocalMux I__2413 (
            .O(N__21336),
            .I(N__21328));
    LocalMux I__2412 (
            .O(N__21333),
            .I(N__21325));
    Span4Mux_v I__2411 (
            .O(N__21328),
            .I(N__21322));
    Span4Mux_v I__2410 (
            .O(N__21325),
            .I(N__21319));
    Span4Mux_v I__2409 (
            .O(N__21322),
            .I(N__21314));
    Span4Mux_v I__2408 (
            .O(N__21319),
            .I(N__21314));
    Odrv4 I__2407 (
            .O(N__21314),
            .I(\pid_alt.error_2 ));
    InMux I__2406 (
            .O(N__21311),
            .I(\pid_alt.error_cry_1 ));
    InMux I__2405 (
            .O(N__21308),
            .I(N__21305));
    LocalMux I__2404 (
            .O(N__21305),
            .I(N__21300));
    InMux I__2403 (
            .O(N__21304),
            .I(N__21297));
    InMux I__2402 (
            .O(N__21303),
            .I(N__21294));
    Span4Mux_s3_h I__2401 (
            .O(N__21300),
            .I(N__21291));
    LocalMux I__2400 (
            .O(N__21297),
            .I(N__21288));
    LocalMux I__2399 (
            .O(N__21294),
            .I(N__21285));
    Span4Mux_v I__2398 (
            .O(N__21291),
            .I(N__21282));
    Span4Mux_s3_h I__2397 (
            .O(N__21288),
            .I(N__21279));
    Span4Mux_v I__2396 (
            .O(N__21285),
            .I(N__21276));
    Span4Mux_v I__2395 (
            .O(N__21282),
            .I(N__21273));
    Span4Mux_v I__2394 (
            .O(N__21279),
            .I(N__21270));
    Span4Mux_h I__2393 (
            .O(N__21276),
            .I(N__21267));
    Odrv4 I__2392 (
            .O(N__21273),
            .I(\pid_alt.error_3 ));
    Odrv4 I__2391 (
            .O(N__21270),
            .I(\pid_alt.error_3 ));
    Odrv4 I__2390 (
            .O(N__21267),
            .I(\pid_alt.error_3 ));
    InMux I__2389 (
            .O(N__21260),
            .I(\pid_alt.error_cry_2 ));
    CascadeMux I__2388 (
            .O(N__21257),
            .I(N__21253));
    CascadeMux I__2387 (
            .O(N__21256),
            .I(N__21250));
    InMux I__2386 (
            .O(N__21253),
            .I(N__21247));
    InMux I__2385 (
            .O(N__21250),
            .I(N__21244));
    LocalMux I__2384 (
            .O(N__21247),
            .I(alt_command_0));
    LocalMux I__2383 (
            .O(N__21244),
            .I(alt_command_0));
    InMux I__2382 (
            .O(N__21239),
            .I(N__21236));
    LocalMux I__2381 (
            .O(N__21236),
            .I(N__21233));
    Span4Mux_s1_h I__2380 (
            .O(N__21233),
            .I(N__21229));
    InMux I__2379 (
            .O(N__21232),
            .I(N__21226));
    Span4Mux_v I__2378 (
            .O(N__21229),
            .I(N__21220));
    LocalMux I__2377 (
            .O(N__21226),
            .I(N__21220));
    InMux I__2376 (
            .O(N__21225),
            .I(N__21217));
    Span4Mux_v I__2375 (
            .O(N__21220),
            .I(N__21214));
    LocalMux I__2374 (
            .O(N__21217),
            .I(N__21211));
    Span4Mux_v I__2373 (
            .O(N__21214),
            .I(N__21208));
    Span4Mux_s3_h I__2372 (
            .O(N__21211),
            .I(N__21205));
    Span4Mux_s1_h I__2371 (
            .O(N__21208),
            .I(N__21202));
    Span4Mux_v I__2370 (
            .O(N__21205),
            .I(N__21199));
    Odrv4 I__2369 (
            .O(N__21202),
            .I(\pid_alt.error_4 ));
    Odrv4 I__2368 (
            .O(N__21199),
            .I(\pid_alt.error_4 ));
    InMux I__2367 (
            .O(N__21194),
            .I(\pid_alt.error_cry_3 ));
    InMux I__2366 (
            .O(N__21191),
            .I(N__21188));
    LocalMux I__2365 (
            .O(N__21188),
            .I(drone_altitude_i_5));
    CascadeMux I__2364 (
            .O(N__21185),
            .I(N__21181));
    InMux I__2363 (
            .O(N__21184),
            .I(N__21178));
    InMux I__2362 (
            .O(N__21181),
            .I(N__21175));
    LocalMux I__2361 (
            .O(N__21178),
            .I(alt_command_1));
    LocalMux I__2360 (
            .O(N__21175),
            .I(alt_command_1));
    InMux I__2359 (
            .O(N__21170),
            .I(N__21166));
    InMux I__2358 (
            .O(N__21169),
            .I(N__21162));
    LocalMux I__2357 (
            .O(N__21166),
            .I(N__21159));
    InMux I__2356 (
            .O(N__21165),
            .I(N__21156));
    LocalMux I__2355 (
            .O(N__21162),
            .I(N__21153));
    Span12Mux_s2_h I__2354 (
            .O(N__21159),
            .I(N__21150));
    LocalMux I__2353 (
            .O(N__21156),
            .I(N__21147));
    Span4Mux_s3_h I__2352 (
            .O(N__21153),
            .I(N__21144));
    Span12Mux_v I__2351 (
            .O(N__21150),
            .I(N__21141));
    Span12Mux_s3_h I__2350 (
            .O(N__21147),
            .I(N__21138));
    Span4Mux_v I__2349 (
            .O(N__21144),
            .I(N__21135));
    Odrv12 I__2348 (
            .O(N__21141),
            .I(\pid_alt.error_5 ));
    Odrv12 I__2347 (
            .O(N__21138),
            .I(\pid_alt.error_5 ));
    Odrv4 I__2346 (
            .O(N__21135),
            .I(\pid_alt.error_5 ));
    InMux I__2345 (
            .O(N__21128),
            .I(\pid_alt.error_cry_4 ));
    InMux I__2344 (
            .O(N__21125),
            .I(N__21122));
    LocalMux I__2343 (
            .O(N__21122),
            .I(drone_altitude_i_6));
    InMux I__2342 (
            .O(N__21119),
            .I(N__21110));
    InMux I__2341 (
            .O(N__21118),
            .I(N__21110));
    InMux I__2340 (
            .O(N__21117),
            .I(N__21110));
    LocalMux I__2339 (
            .O(N__21110),
            .I(N__21107));
    Span12Mux_s10_h I__2338 (
            .O(N__21107),
            .I(N__21104));
    Span12Mux_v I__2337 (
            .O(N__21104),
            .I(N__21101));
    Odrv12 I__2336 (
            .O(N__21101),
            .I(\pid_alt.error_d_regZ0Z_16 ));
    CascadeMux I__2335 (
            .O(N__21098),
            .I(N__21095));
    InMux I__2334 (
            .O(N__21095),
            .I(N__21089));
    InMux I__2333 (
            .O(N__21094),
            .I(N__21089));
    LocalMux I__2332 (
            .O(N__21089),
            .I(\pid_alt.error_d_reg_prevZ0Z_16 ));
    InMux I__2331 (
            .O(N__21086),
            .I(N__21080));
    InMux I__2330 (
            .O(N__21085),
            .I(N__21080));
    LocalMux I__2329 (
            .O(N__21080),
            .I(N__21077));
    Span4Mux_h I__2328 (
            .O(N__21077),
            .I(N__21074));
    Span4Mux_v I__2327 (
            .O(N__21074),
            .I(N__21071));
    Odrv4 I__2326 (
            .O(N__21071),
            .I(\pid_alt.error_p_regZ0Z_16 ));
    InMux I__2325 (
            .O(N__21068),
            .I(N__21065));
    LocalMux I__2324 (
            .O(N__21065),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ));
    CascadeMux I__2323 (
            .O(N__21062),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ));
    CascadeMux I__2322 (
            .O(N__21059),
            .I(\Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ));
    CascadeMux I__2321 (
            .O(N__21056),
            .I(\Commands_frame_decoder.source_CH1data8_cascade_ ));
    InMux I__2320 (
            .O(N__21053),
            .I(N__21050));
    LocalMux I__2319 (
            .O(N__21050),
            .I(N__21047));
    Span4Mux_h I__2318 (
            .O(N__21047),
            .I(N__21044));
    Span4Mux_v I__2317 (
            .O(N__21044),
            .I(N__21041));
    Odrv4 I__2316 (
            .O(N__21041),
            .I(\pid_alt.error_i_regZ0Z_19 ));
    InMux I__2315 (
            .O(N__21038),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_18 ));
    InMux I__2314 (
            .O(N__21035),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_19 ));
    InMux I__2313 (
            .O(N__21032),
            .I(N__21026));
    InMux I__2312 (
            .O(N__21031),
            .I(N__21026));
    LocalMux I__2311 (
            .O(N__21026),
            .I(N__21023));
    Span4Mux_h I__2310 (
            .O(N__21023),
            .I(N__21020));
    Span4Mux_v I__2309 (
            .O(N__21020),
            .I(N__21017));
    Odrv4 I__2308 (
            .O(N__21017),
            .I(\pid_alt.error_i_regZ0Z_20 ));
    InMux I__2307 (
            .O(N__21014),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_20 ));
    InMux I__2306 (
            .O(N__21011),
            .I(N__21008));
    LocalMux I__2305 (
            .O(N__21008),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ));
    CascadeMux I__2304 (
            .O(N__21005),
            .I(N__21001));
    InMux I__2303 (
            .O(N__21004),
            .I(N__20998));
    InMux I__2302 (
            .O(N__21001),
            .I(N__20995));
    LocalMux I__2301 (
            .O(N__20998),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    LocalMux I__2300 (
            .O(N__20995),
            .I(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ));
    InMux I__2299 (
            .O(N__20990),
            .I(N__20987));
    LocalMux I__2298 (
            .O(N__20987),
            .I(N__20982));
    InMux I__2297 (
            .O(N__20986),
            .I(N__20979));
    InMux I__2296 (
            .O(N__20985),
            .I(N__20976));
    Odrv4 I__2295 (
            .O(N__20982),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__2294 (
            .O(N__20979),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    LocalMux I__2293 (
            .O(N__20976),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ));
    InMux I__2292 (
            .O(N__20969),
            .I(N__20965));
    InMux I__2291 (
            .O(N__20968),
            .I(N__20962));
    LocalMux I__2290 (
            .O(N__20965),
            .I(N__20959));
    LocalMux I__2289 (
            .O(N__20962),
            .I(N__20954));
    Span4Mux_h I__2288 (
            .O(N__20959),
            .I(N__20954));
    Span4Mux_v I__2287 (
            .O(N__20954),
            .I(N__20951));
    Odrv4 I__2286 (
            .O(N__20951),
            .I(\pid_alt.error_p_regZ0Z_17 ));
    InMux I__2285 (
            .O(N__20948),
            .I(N__20945));
    LocalMux I__2284 (
            .O(N__20945),
            .I(N__20941));
    InMux I__2283 (
            .O(N__20944),
            .I(N__20938));
    Span4Mux_h I__2282 (
            .O(N__20941),
            .I(N__20935));
    LocalMux I__2281 (
            .O(N__20938),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    Odrv4 I__2280 (
            .O(N__20935),
            .I(\pid_alt.error_d_reg_prevZ0Z_17 ));
    InMux I__2279 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__2278 (
            .O(N__20927),
            .I(N__20922));
    InMux I__2277 (
            .O(N__20926),
            .I(N__20917));
    InMux I__2276 (
            .O(N__20925),
            .I(N__20917));
    Span4Mux_v I__2275 (
            .O(N__20922),
            .I(N__20914));
    LocalMux I__2274 (
            .O(N__20917),
            .I(N__20911));
    Span4Mux_v I__2273 (
            .O(N__20914),
            .I(N__20908));
    Span12Mux_v I__2272 (
            .O(N__20911),
            .I(N__20905));
    Span4Mux_v I__2271 (
            .O(N__20908),
            .I(N__20902));
    Odrv12 I__2270 (
            .O(N__20905),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    Odrv4 I__2269 (
            .O(N__20902),
            .I(\pid_alt.error_d_regZ0Z_17 ));
    InMux I__2268 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__2267 (
            .O(N__20894),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ));
    CascadeMux I__2266 (
            .O(N__20891),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ));
    InMux I__2265 (
            .O(N__20888),
            .I(N__20882));
    InMux I__2264 (
            .O(N__20887),
            .I(N__20882));
    LocalMux I__2263 (
            .O(N__20882),
            .I(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ));
    CascadeMux I__2262 (
            .O(N__20879),
            .I(N__20876));
    InMux I__2261 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2260 (
            .O(N__20873),
            .I(N__20870));
    Span4Mux_v I__2259 (
            .O(N__20870),
            .I(N__20867));
    Odrv4 I__2258 (
            .O(N__20867),
            .I(\pid_alt.error_i_regZ0Z_11 ));
    InMux I__2257 (
            .O(N__20864),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_10 ));
    CascadeMux I__2256 (
            .O(N__20861),
            .I(N__20858));
    InMux I__2255 (
            .O(N__20858),
            .I(N__20855));
    LocalMux I__2254 (
            .O(N__20855),
            .I(N__20852));
    Span4Mux_h I__2253 (
            .O(N__20852),
            .I(N__20849));
    Span4Mux_v I__2252 (
            .O(N__20849),
            .I(N__20846));
    Odrv4 I__2251 (
            .O(N__20846),
            .I(\pid_alt.error_i_regZ0Z_12 ));
    InMux I__2250 (
            .O(N__20843),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_11 ));
    CascadeMux I__2249 (
            .O(N__20840),
            .I(N__20837));
    InMux I__2248 (
            .O(N__20837),
            .I(N__20834));
    LocalMux I__2247 (
            .O(N__20834),
            .I(N__20831));
    Span4Mux_h I__2246 (
            .O(N__20831),
            .I(N__20828));
    Span4Mux_v I__2245 (
            .O(N__20828),
            .I(N__20825));
    Odrv4 I__2244 (
            .O(N__20825),
            .I(\pid_alt.error_i_regZ0Z_13 ));
    InMux I__2243 (
            .O(N__20822),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_12 ));
    InMux I__2242 (
            .O(N__20819),
            .I(N__20816));
    LocalMux I__2241 (
            .O(N__20816),
            .I(N__20813));
    Span4Mux_v I__2240 (
            .O(N__20813),
            .I(N__20810));
    Span4Mux_v I__2239 (
            .O(N__20810),
            .I(N__20807));
    Odrv4 I__2238 (
            .O(N__20807),
            .I(\pid_alt.error_i_regZ0Z_14 ));
    InMux I__2237 (
            .O(N__20804),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_13 ));
    InMux I__2236 (
            .O(N__20801),
            .I(N__20798));
    LocalMux I__2235 (
            .O(N__20798),
            .I(N__20795));
    Span4Mux_h I__2234 (
            .O(N__20795),
            .I(N__20792));
    Span4Mux_v I__2233 (
            .O(N__20792),
            .I(N__20789));
    Odrv4 I__2232 (
            .O(N__20789),
            .I(\pid_alt.error_i_regZ0Z_15 ));
    InMux I__2231 (
            .O(N__20786),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_14 ));
    InMux I__2230 (
            .O(N__20783),
            .I(N__20780));
    LocalMux I__2229 (
            .O(N__20780),
            .I(N__20777));
    Span4Mux_h I__2228 (
            .O(N__20777),
            .I(N__20774));
    Span4Mux_v I__2227 (
            .O(N__20774),
            .I(N__20771));
    Odrv4 I__2226 (
            .O(N__20771),
            .I(\pid_alt.error_i_regZ0Z_16 ));
    InMux I__2225 (
            .O(N__20768),
            .I(bfn_3_16_0_));
    InMux I__2224 (
            .O(N__20765),
            .I(N__20762));
    LocalMux I__2223 (
            .O(N__20762),
            .I(N__20759));
    Span4Mux_v I__2222 (
            .O(N__20759),
            .I(N__20756));
    Span4Mux_v I__2221 (
            .O(N__20756),
            .I(N__20753));
    Odrv4 I__2220 (
            .O(N__20753),
            .I(\pid_alt.error_i_regZ0Z_17 ));
    InMux I__2219 (
            .O(N__20750),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_16 ));
    InMux I__2218 (
            .O(N__20747),
            .I(N__20744));
    LocalMux I__2217 (
            .O(N__20744),
            .I(N__20741));
    Span12Mux_v I__2216 (
            .O(N__20741),
            .I(N__20738));
    Odrv12 I__2215 (
            .O(N__20738),
            .I(\pid_alt.error_i_regZ0Z_18 ));
    InMux I__2214 (
            .O(N__20735),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_17 ));
    CascadeMux I__2213 (
            .O(N__20732),
            .I(N__20729));
    InMux I__2212 (
            .O(N__20729),
            .I(N__20726));
    LocalMux I__2211 (
            .O(N__20726),
            .I(N__20723));
    Span4Mux_v I__2210 (
            .O(N__20723),
            .I(N__20720));
    Odrv4 I__2209 (
            .O(N__20720),
            .I(\pid_alt.error_i_regZ0Z_3 ));
    InMux I__2208 (
            .O(N__20717),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_2 ));
    CascadeMux I__2207 (
            .O(N__20714),
            .I(N__20711));
    InMux I__2206 (
            .O(N__20711),
            .I(N__20708));
    LocalMux I__2205 (
            .O(N__20708),
            .I(N__20705));
    Span4Mux_h I__2204 (
            .O(N__20705),
            .I(N__20702));
    Span4Mux_v I__2203 (
            .O(N__20702),
            .I(N__20699));
    Odrv4 I__2202 (
            .O(N__20699),
            .I(\pid_alt.error_i_regZ0Z_4 ));
    InMux I__2201 (
            .O(N__20696),
            .I(N__20691));
    InMux I__2200 (
            .O(N__20695),
            .I(N__20686));
    InMux I__2199 (
            .O(N__20694),
            .I(N__20686));
    LocalMux I__2198 (
            .O(N__20691),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    LocalMux I__2197 (
            .O(N__20686),
            .I(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ));
    InMux I__2196 (
            .O(N__20681),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_3 ));
    InMux I__2195 (
            .O(N__20678),
            .I(N__20675));
    LocalMux I__2194 (
            .O(N__20675),
            .I(N__20672));
    Span4Mux_v I__2193 (
            .O(N__20672),
            .I(N__20669));
    Odrv4 I__2192 (
            .O(N__20669),
            .I(\pid_alt.error_i_regZ0Z_5 ));
    InMux I__2191 (
            .O(N__20666),
            .I(N__20661));
    InMux I__2190 (
            .O(N__20665),
            .I(N__20656));
    InMux I__2189 (
            .O(N__20664),
            .I(N__20656));
    LocalMux I__2188 (
            .O(N__20661),
            .I(\pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5 ));
    LocalMux I__2187 (
            .O(N__20656),
            .I(\pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5 ));
    InMux I__2186 (
            .O(N__20651),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_4 ));
    InMux I__2185 (
            .O(N__20648),
            .I(N__20644));
    InMux I__2184 (
            .O(N__20647),
            .I(N__20641));
    LocalMux I__2183 (
            .O(N__20644),
            .I(N__20638));
    LocalMux I__2182 (
            .O(N__20641),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    Odrv4 I__2181 (
            .O(N__20638),
            .I(\pid_alt.error_i_acummZ0Z_6 ));
    CascadeMux I__2180 (
            .O(N__20633),
            .I(N__20630));
    InMux I__2179 (
            .O(N__20630),
            .I(N__20627));
    LocalMux I__2178 (
            .O(N__20627),
            .I(N__20624));
    Span4Mux_v I__2177 (
            .O(N__20624),
            .I(N__20621));
    Odrv4 I__2176 (
            .O(N__20621),
            .I(\pid_alt.error_i_regZ0Z_6 ));
    InMux I__2175 (
            .O(N__20618),
            .I(N__20612));
    InMux I__2174 (
            .O(N__20617),
            .I(N__20612));
    LocalMux I__2173 (
            .O(N__20612),
            .I(N__20608));
    InMux I__2172 (
            .O(N__20611),
            .I(N__20605));
    Span4Mux_v I__2171 (
            .O(N__20608),
            .I(N__20602));
    LocalMux I__2170 (
            .O(N__20605),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    Odrv4 I__2169 (
            .O(N__20602),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ));
    InMux I__2168 (
            .O(N__20597),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_5 ));
    CascadeMux I__2167 (
            .O(N__20594),
            .I(N__20591));
    InMux I__2166 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__2165 (
            .O(N__20588),
            .I(N__20585));
    Span4Mux_v I__2164 (
            .O(N__20585),
            .I(N__20582));
    Odrv4 I__2163 (
            .O(N__20582),
            .I(\pid_alt.error_i_regZ0Z_7 ));
    InMux I__2162 (
            .O(N__20579),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_6 ));
    InMux I__2161 (
            .O(N__20576),
            .I(N__20572));
    InMux I__2160 (
            .O(N__20575),
            .I(N__20569));
    LocalMux I__2159 (
            .O(N__20572),
            .I(N__20566));
    LocalMux I__2158 (
            .O(N__20569),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    Odrv4 I__2157 (
            .O(N__20566),
            .I(\pid_alt.error_i_acummZ0Z_8 ));
    CascadeMux I__2156 (
            .O(N__20561),
            .I(N__20558));
    InMux I__2155 (
            .O(N__20558),
            .I(N__20555));
    LocalMux I__2154 (
            .O(N__20555),
            .I(N__20552));
    Span4Mux_h I__2153 (
            .O(N__20552),
            .I(N__20549));
    Span4Mux_v I__2152 (
            .O(N__20549),
            .I(N__20546));
    Odrv4 I__2151 (
            .O(N__20546),
            .I(\pid_alt.error_i_regZ0Z_8 ));
    InMux I__2150 (
            .O(N__20543),
            .I(bfn_3_15_0_));
    InMux I__2149 (
            .O(N__20540),
            .I(N__20536));
    InMux I__2148 (
            .O(N__20539),
            .I(N__20533));
    LocalMux I__2147 (
            .O(N__20536),
            .I(N__20530));
    LocalMux I__2146 (
            .O(N__20533),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    Odrv4 I__2145 (
            .O(N__20530),
            .I(\pid_alt.error_i_acummZ0Z_9 ));
    CascadeMux I__2144 (
            .O(N__20525),
            .I(N__20522));
    InMux I__2143 (
            .O(N__20522),
            .I(N__20519));
    LocalMux I__2142 (
            .O(N__20519),
            .I(N__20516));
    Span4Mux_h I__2141 (
            .O(N__20516),
            .I(N__20513));
    Span4Mux_v I__2140 (
            .O(N__20513),
            .I(N__20510));
    Odrv4 I__2139 (
            .O(N__20510),
            .I(\pid_alt.error_i_regZ0Z_9 ));
    InMux I__2138 (
            .O(N__20507),
            .I(N__20502));
    InMux I__2137 (
            .O(N__20506),
            .I(N__20497));
    InMux I__2136 (
            .O(N__20505),
            .I(N__20497));
    LocalMux I__2135 (
            .O(N__20502),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    LocalMux I__2134 (
            .O(N__20497),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ));
    InMux I__2133 (
            .O(N__20492),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_8 ));
    InMux I__2132 (
            .O(N__20489),
            .I(N__20485));
    InMux I__2131 (
            .O(N__20488),
            .I(N__20482));
    LocalMux I__2130 (
            .O(N__20485),
            .I(N__20479));
    LocalMux I__2129 (
            .O(N__20482),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    Odrv12 I__2128 (
            .O(N__20479),
            .I(\pid_alt.error_i_acummZ0Z_10 ));
    CascadeMux I__2127 (
            .O(N__20474),
            .I(N__20471));
    InMux I__2126 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__2125 (
            .O(N__20468),
            .I(N__20465));
    Span4Mux_v I__2124 (
            .O(N__20465),
            .I(N__20462));
    Odrv4 I__2123 (
            .O(N__20462),
            .I(\pid_alt.error_i_regZ0Z_10 ));
    InMux I__2122 (
            .O(N__20459),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_9 ));
    InMux I__2121 (
            .O(N__20456),
            .I(N__20451));
    InMux I__2120 (
            .O(N__20455),
            .I(N__20446));
    InMux I__2119 (
            .O(N__20454),
            .I(N__20446));
    LocalMux I__2118 (
            .O(N__20451),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    LocalMux I__2117 (
            .O(N__20446),
            .I(\pid_alt.error_i_acumm_preregZ0Z_6 ));
    InMux I__2116 (
            .O(N__20441),
            .I(N__20436));
    CascadeMux I__2115 (
            .O(N__20440),
            .I(N__20433));
    CascadeMux I__2114 (
            .O(N__20439),
            .I(N__20430));
    LocalMux I__2113 (
            .O(N__20436),
            .I(N__20427));
    InMux I__2112 (
            .O(N__20433),
            .I(N__20422));
    InMux I__2111 (
            .O(N__20430),
            .I(N__20422));
    Odrv4 I__2110 (
            .O(N__20427),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    LocalMux I__2109 (
            .O(N__20422),
            .I(\pid_alt.error_i_acumm_preregZ0Z_10 ));
    CascadeMux I__2108 (
            .O(N__20417),
            .I(N__20414));
    InMux I__2107 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__2106 (
            .O(N__20411),
            .I(N__20406));
    InMux I__2105 (
            .O(N__20410),
            .I(N__20403));
    InMux I__2104 (
            .O(N__20409),
            .I(N__20400));
    Odrv4 I__2103 (
            .O(N__20406),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__2102 (
            .O(N__20403),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    LocalMux I__2101 (
            .O(N__20400),
            .I(\pid_alt.error_i_acumm_preregZ0Z_9 ));
    InMux I__2100 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__2099 (
            .O(N__20390),
            .I(N__20385));
    InMux I__2098 (
            .O(N__20389),
            .I(N__20382));
    InMux I__2097 (
            .O(N__20388),
            .I(N__20379));
    Odrv4 I__2096 (
            .O(N__20385),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__2095 (
            .O(N__20382),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    LocalMux I__2094 (
            .O(N__20379),
            .I(\pid_alt.error_i_acumm_preregZ0Z_8 ));
    CascadeMux I__2093 (
            .O(N__20372),
            .I(N__20369));
    InMux I__2092 (
            .O(N__20369),
            .I(N__20366));
    LocalMux I__2091 (
            .O(N__20366),
            .I(N__20363));
    Odrv4 I__2090 (
            .O(N__20363),
            .I(\pid_alt.error_i_regZ0Z_1 ));
    InMux I__2089 (
            .O(N__20360),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_0 ));
    CascadeMux I__2088 (
            .O(N__20357),
            .I(N__20354));
    InMux I__2087 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2086 (
            .O(N__20351),
            .I(N__20348));
    Span4Mux_v I__2085 (
            .O(N__20348),
            .I(N__20345));
    Odrv4 I__2084 (
            .O(N__20345),
            .I(\pid_alt.error_i_regZ0Z_2 ));
    InMux I__2083 (
            .O(N__20342),
            .I(\pid_alt.un1_error_i_acumm_prereg_cry_1 ));
    InMux I__2082 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__2081 (
            .O(N__20336),
            .I(N__20333));
    Odrv12 I__2080 (
            .O(N__20333),
            .I(\pid_alt.O_2_6 ));
    CEMux I__2079 (
            .O(N__20330),
            .I(N__20279));
    CEMux I__2078 (
            .O(N__20329),
            .I(N__20279));
    CEMux I__2077 (
            .O(N__20328),
            .I(N__20279));
    CEMux I__2076 (
            .O(N__20327),
            .I(N__20279));
    CEMux I__2075 (
            .O(N__20326),
            .I(N__20279));
    CEMux I__2074 (
            .O(N__20325),
            .I(N__20279));
    CEMux I__2073 (
            .O(N__20324),
            .I(N__20279));
    CEMux I__2072 (
            .O(N__20323),
            .I(N__20279));
    CEMux I__2071 (
            .O(N__20322),
            .I(N__20279));
    CEMux I__2070 (
            .O(N__20321),
            .I(N__20279));
    CEMux I__2069 (
            .O(N__20320),
            .I(N__20279));
    CEMux I__2068 (
            .O(N__20319),
            .I(N__20279));
    CEMux I__2067 (
            .O(N__20318),
            .I(N__20279));
    CEMux I__2066 (
            .O(N__20317),
            .I(N__20279));
    CEMux I__2065 (
            .O(N__20316),
            .I(N__20279));
    CEMux I__2064 (
            .O(N__20315),
            .I(N__20279));
    CEMux I__2063 (
            .O(N__20314),
            .I(N__20279));
    GlobalMux I__2062 (
            .O(N__20279),
            .I(N__20276));
    gio2CtrlBuf I__2061 (
            .O(N__20276),
            .I(\pid_alt.N_850_0_g ));
    InMux I__2060 (
            .O(N__20273),
            .I(N__20270));
    LocalMux I__2059 (
            .O(N__20270),
            .I(N__20267));
    Span4Mux_s2_h I__2058 (
            .O(N__20267),
            .I(N__20264));
    Odrv4 I__2057 (
            .O(N__20264),
            .I(alt_kp_2));
    InMux I__2056 (
            .O(N__20261),
            .I(N__20258));
    LocalMux I__2055 (
            .O(N__20258),
            .I(N__20255));
    Span4Mux_v I__2054 (
            .O(N__20255),
            .I(N__20252));
    Sp12to4 I__2053 (
            .O(N__20252),
            .I(N__20249));
    Odrv12 I__2052 (
            .O(N__20249),
            .I(alt_kp_3));
    InMux I__2051 (
            .O(N__20246),
            .I(N__20243));
    LocalMux I__2050 (
            .O(N__20243),
            .I(N__20240));
    Span4Mux_s3_h I__2049 (
            .O(N__20240),
            .I(N__20237));
    Odrv4 I__2048 (
            .O(N__20237),
            .I(alt_kp_5));
    InMux I__2047 (
            .O(N__20234),
            .I(N__20231));
    LocalMux I__2046 (
            .O(N__20231),
            .I(N__20228));
    Span4Mux_s2_h I__2045 (
            .O(N__20228),
            .I(N__20225));
    Odrv4 I__2044 (
            .O(N__20225),
            .I(alt_kp_6));
    InMux I__2043 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__2042 (
            .O(N__20219),
            .I(N__20216));
    Span4Mux_h I__2041 (
            .O(N__20216),
            .I(N__20213));
    Odrv4 I__2040 (
            .O(N__20213),
            .I(alt_kd_3));
    InMux I__2039 (
            .O(N__20210),
            .I(N__20207));
    LocalMux I__2038 (
            .O(N__20207),
            .I(N__20204));
    Span4Mux_s3_h I__2037 (
            .O(N__20204),
            .I(N__20201));
    Odrv4 I__2036 (
            .O(N__20201),
            .I(alt_kd_0));
    InMux I__2035 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__2034 (
            .O(N__20195),
            .I(N__20192));
    Span4Mux_s3_h I__2033 (
            .O(N__20192),
            .I(N__20189));
    Odrv4 I__2032 (
            .O(N__20189),
            .I(alt_kd_4));
    InMux I__2031 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__2030 (
            .O(N__20183),
            .I(\dron_frame_decoder_1.drone_altitude_10 ));
    InMux I__2029 (
            .O(N__20180),
            .I(N__20177));
    LocalMux I__2028 (
            .O(N__20177),
            .I(\dron_frame_decoder_1.drone_altitude_8 ));
    InMux I__2027 (
            .O(N__20174),
            .I(N__20171));
    LocalMux I__2026 (
            .O(N__20171),
            .I(\dron_frame_decoder_1.drone_altitude_9 ));
    InMux I__2025 (
            .O(N__20168),
            .I(N__20162));
    InMux I__2024 (
            .O(N__20167),
            .I(N__20162));
    LocalMux I__2023 (
            .O(N__20162),
            .I(N__20159));
    Span4Mux_v I__2022 (
            .O(N__20159),
            .I(N__20156));
    Odrv4 I__2021 (
            .O(N__20156),
            .I(\pid_alt.error_p_regZ0Z_5 ));
    InMux I__2020 (
            .O(N__20153),
            .I(N__20147));
    InMux I__2019 (
            .O(N__20152),
            .I(N__20147));
    LocalMux I__2018 (
            .O(N__20147),
            .I(\pid_alt.error_d_reg_prevZ0Z_5 ));
    InMux I__2017 (
            .O(N__20144),
            .I(N__20135));
    InMux I__2016 (
            .O(N__20143),
            .I(N__20135));
    InMux I__2015 (
            .O(N__20142),
            .I(N__20135));
    LocalMux I__2014 (
            .O(N__20135),
            .I(N__20132));
    Span12Mux_v I__2013 (
            .O(N__20132),
            .I(N__20129));
    Odrv12 I__2012 (
            .O(N__20129),
            .I(\pid_alt.error_d_regZ0Z_5 ));
    CascadeMux I__2011 (
            .O(N__20126),
            .I(N__20123));
    InMux I__2010 (
            .O(N__20123),
            .I(N__20117));
    InMux I__2009 (
            .O(N__20122),
            .I(N__20117));
    LocalMux I__2008 (
            .O(N__20117),
            .I(N__20114));
    Odrv4 I__2007 (
            .O(N__20114),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ));
    InMux I__2006 (
            .O(N__20111),
            .I(N__20105));
    InMux I__2005 (
            .O(N__20110),
            .I(N__20105));
    LocalMux I__2004 (
            .O(N__20105),
            .I(N__20102));
    Span4Mux_v I__2003 (
            .O(N__20102),
            .I(N__20099));
    Odrv4 I__2002 (
            .O(N__20099),
            .I(\pid_alt.error_p_regZ0Z_6 ));
    InMux I__2001 (
            .O(N__20096),
            .I(N__20090));
    InMux I__2000 (
            .O(N__20095),
            .I(N__20090));
    LocalMux I__1999 (
            .O(N__20090),
            .I(\pid_alt.error_d_reg_prevZ0Z_6 ));
    InMux I__1998 (
            .O(N__20087),
            .I(N__20078));
    InMux I__1997 (
            .O(N__20086),
            .I(N__20078));
    InMux I__1996 (
            .O(N__20085),
            .I(N__20078));
    LocalMux I__1995 (
            .O(N__20078),
            .I(N__20075));
    Span12Mux_v I__1994 (
            .O(N__20075),
            .I(N__20072));
    Odrv12 I__1993 (
            .O(N__20072),
            .I(\pid_alt.error_d_regZ0Z_6 ));
    InMux I__1992 (
            .O(N__20069),
            .I(N__20066));
    LocalMux I__1991 (
            .O(N__20066),
            .I(N__20063));
    Span4Mux_h I__1990 (
            .O(N__20063),
            .I(N__20060));
    Odrv4 I__1989 (
            .O(N__20060),
            .I(\pid_side.O_0_24 ));
    InMux I__1988 (
            .O(N__20057),
            .I(N__20054));
    LocalMux I__1987 (
            .O(N__20054),
            .I(N__20051));
    Span4Mux_h I__1986 (
            .O(N__20051),
            .I(N__20048));
    Odrv4 I__1985 (
            .O(N__20048),
            .I(\pid_side.O_0_13 ));
    InMux I__1984 (
            .O(N__20045),
            .I(N__20039));
    InMux I__1983 (
            .O(N__20044),
            .I(N__20039));
    LocalMux I__1982 (
            .O(N__20039),
            .I(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ));
    InMux I__1981 (
            .O(N__20036),
            .I(N__20027));
    InMux I__1980 (
            .O(N__20035),
            .I(N__20027));
    InMux I__1979 (
            .O(N__20034),
            .I(N__20027));
    LocalMux I__1978 (
            .O(N__20027),
            .I(N__20024));
    Span4Mux_v I__1977 (
            .O(N__20024),
            .I(N__20021));
    Span4Mux_v I__1976 (
            .O(N__20021),
            .I(N__20018));
    Span4Mux_v I__1975 (
            .O(N__20018),
            .I(N__20015));
    Odrv4 I__1974 (
            .O(N__20015),
            .I(\pid_alt.error_d_regZ0Z_18 ));
    CascadeMux I__1973 (
            .O(N__20012),
            .I(N__20009));
    InMux I__1972 (
            .O(N__20009),
            .I(N__20003));
    InMux I__1971 (
            .O(N__20008),
            .I(N__20003));
    LocalMux I__1970 (
            .O(N__20003),
            .I(\pid_alt.error_d_reg_prevZ0Z_18 ));
    InMux I__1969 (
            .O(N__20000),
            .I(N__19994));
    InMux I__1968 (
            .O(N__19999),
            .I(N__19994));
    LocalMux I__1967 (
            .O(N__19994),
            .I(N__19991));
    Span4Mux_v I__1966 (
            .O(N__19991),
            .I(N__19988));
    Odrv4 I__1965 (
            .O(N__19988),
            .I(\pid_alt.error_p_regZ0Z_18 ));
    InMux I__1964 (
            .O(N__19985),
            .I(N__19982));
    LocalMux I__1963 (
            .O(N__19982),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ));
    InMux I__1962 (
            .O(N__19979),
            .I(N__19973));
    InMux I__1961 (
            .O(N__19978),
            .I(N__19973));
    LocalMux I__1960 (
            .O(N__19973),
            .I(N__19970));
    Odrv4 I__1959 (
            .O(N__19970),
            .I(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ));
    CascadeMux I__1958 (
            .O(N__19967),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ));
    InMux I__1957 (
            .O(N__19964),
            .I(N__19961));
    LocalMux I__1956 (
            .O(N__19961),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ));
    CascadeMux I__1955 (
            .O(N__19958),
            .I(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ));
    InMux I__1954 (
            .O(N__19955),
            .I(N__19949));
    InMux I__1953 (
            .O(N__19954),
            .I(N__19949));
    LocalMux I__1952 (
            .O(N__19949),
            .I(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ));
    CascadeMux I__1951 (
            .O(N__19946),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ));
    InMux I__1950 (
            .O(N__19943),
            .I(N__19934));
    InMux I__1949 (
            .O(N__19942),
            .I(N__19934));
    InMux I__1948 (
            .O(N__19941),
            .I(N__19934));
    LocalMux I__1947 (
            .O(N__19934),
            .I(N__19931));
    Span4Mux_v I__1946 (
            .O(N__19931),
            .I(N__19928));
    Span4Mux_v I__1945 (
            .O(N__19928),
            .I(N__19925));
    Odrv4 I__1944 (
            .O(N__19925),
            .I(\pid_alt.error_d_regZ0Z_9 ));
    CascadeMux I__1943 (
            .O(N__19922),
            .I(N__19919));
    InMux I__1942 (
            .O(N__19919),
            .I(N__19913));
    InMux I__1941 (
            .O(N__19918),
            .I(N__19913));
    LocalMux I__1940 (
            .O(N__19913),
            .I(\pid_alt.error_d_reg_prevZ0Z_9 ));
    InMux I__1939 (
            .O(N__19910),
            .I(N__19904));
    InMux I__1938 (
            .O(N__19909),
            .I(N__19904));
    LocalMux I__1937 (
            .O(N__19904),
            .I(N__19901));
    Span4Mux_h I__1936 (
            .O(N__19901),
            .I(N__19898));
    Span4Mux_v I__1935 (
            .O(N__19898),
            .I(N__19895));
    Odrv4 I__1934 (
            .O(N__19895),
            .I(\pid_alt.error_p_regZ0Z_9 ));
    InMux I__1933 (
            .O(N__19892),
            .I(N__19889));
    LocalMux I__1932 (
            .O(N__19889),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ));
    InMux I__1931 (
            .O(N__19886),
            .I(N__19880));
    InMux I__1930 (
            .O(N__19885),
            .I(N__19880));
    LocalMux I__1929 (
            .O(N__19880),
            .I(N__19877));
    Span4Mux_h I__1928 (
            .O(N__19877),
            .I(N__19874));
    Odrv4 I__1927 (
            .O(N__19874),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ));
    CascadeMux I__1926 (
            .O(N__19871),
            .I(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ));
    InMux I__1925 (
            .O(N__19868),
            .I(N__19865));
    LocalMux I__1924 (
            .O(N__19865),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ));
    CascadeMux I__1923 (
            .O(N__19862),
            .I(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ));
    InMux I__1922 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__1921 (
            .O(N__19856),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ));
    InMux I__1920 (
            .O(N__19853),
            .I(N__19847));
    InMux I__1919 (
            .O(N__19852),
            .I(N__19847));
    LocalMux I__1918 (
            .O(N__19847),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ));
    CascadeMux I__1917 (
            .O(N__19844),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ));
    InMux I__1916 (
            .O(N__19841),
            .I(N__19835));
    InMux I__1915 (
            .O(N__19840),
            .I(N__19835));
    LocalMux I__1914 (
            .O(N__19835),
            .I(N__19832));
    Span4Mux_v I__1913 (
            .O(N__19832),
            .I(N__19829));
    Span4Mux_v I__1912 (
            .O(N__19829),
            .I(N__19826));
    Odrv4 I__1911 (
            .O(N__19826),
            .I(\pid_alt.error_p_regZ0Z_4 ));
    InMux I__1910 (
            .O(N__19823),
            .I(N__19817));
    InMux I__1909 (
            .O(N__19822),
            .I(N__19817));
    LocalMux I__1908 (
            .O(N__19817),
            .I(N__19814));
    Odrv4 I__1907 (
            .O(N__19814),
            .I(\pid_alt.error_d_reg_prevZ0Z_4 ));
    InMux I__1906 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__1905 (
            .O(N__19808),
            .I(N__19803));
    InMux I__1904 (
            .O(N__19807),
            .I(N__19798));
    InMux I__1903 (
            .O(N__19806),
            .I(N__19798));
    Sp12to4 I__1902 (
            .O(N__19803),
            .I(N__19793));
    LocalMux I__1901 (
            .O(N__19798),
            .I(N__19793));
    Odrv12 I__1900 (
            .O(N__19793),
            .I(\pid_alt.error_d_regZ0Z_4 ));
    CascadeMux I__1899 (
            .O(N__19790),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ));
    InMux I__1898 (
            .O(N__19787),
            .I(N__19784));
    LocalMux I__1897 (
            .O(N__19784),
            .I(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ));
    InMux I__1896 (
            .O(N__19781),
            .I(N__19778));
    LocalMux I__1895 (
            .O(N__19778),
            .I(N__19775));
    Span4Mux_s2_h I__1894 (
            .O(N__19775),
            .I(N__19772));
    Odrv4 I__1893 (
            .O(N__19772),
            .I(alt_ki_5));
    InMux I__1892 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__1891 (
            .O(N__19766),
            .I(N__19763));
    Span4Mux_h I__1890 (
            .O(N__19763),
            .I(N__19760));
    Odrv4 I__1889 (
            .O(N__19760),
            .I(\pid_alt.O_2_5 ));
    InMux I__1888 (
            .O(N__19757),
            .I(N__19754));
    LocalMux I__1887 (
            .O(N__19754),
            .I(N__19751));
    Span4Mux_h I__1886 (
            .O(N__19751),
            .I(N__19748));
    Odrv4 I__1885 (
            .O(N__19748),
            .I(\pid_alt.O_2_4 ));
    InMux I__1884 (
            .O(N__19745),
            .I(N__19742));
    LocalMux I__1883 (
            .O(N__19742),
            .I(N__19739));
    Span4Mux_s2_h I__1882 (
            .O(N__19739),
            .I(N__19736));
    Odrv4 I__1881 (
            .O(N__19736),
            .I(alt_kd_5));
    InMux I__1880 (
            .O(N__19733),
            .I(N__19730));
    LocalMux I__1879 (
            .O(N__19730),
            .I(N__19727));
    Span4Mux_s2_h I__1878 (
            .O(N__19727),
            .I(N__19724));
    Odrv4 I__1877 (
            .O(N__19724),
            .I(alt_kd_1));
    InMux I__1876 (
            .O(N__19721),
            .I(N__19718));
    LocalMux I__1875 (
            .O(N__19718),
            .I(N__19715));
    Span4Mux_h I__1874 (
            .O(N__19715),
            .I(N__19712));
    Odrv4 I__1873 (
            .O(N__19712),
            .I(\pid_alt.O_1_9 ));
    InMux I__1872 (
            .O(N__19709),
            .I(N__19706));
    LocalMux I__1871 (
            .O(N__19706),
            .I(N__19703));
    Span4Mux_v I__1870 (
            .O(N__19703),
            .I(N__19700));
    Odrv4 I__1869 (
            .O(N__19700),
            .I(alt_ki_0));
    InMux I__1868 (
            .O(N__19697),
            .I(N__19694));
    LocalMux I__1867 (
            .O(N__19694),
            .I(N__19691));
    Span4Mux_s2_h I__1866 (
            .O(N__19691),
            .I(N__19688));
    Odrv4 I__1865 (
            .O(N__19688),
            .I(alt_ki_4));
    InMux I__1864 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__1863 (
            .O(N__19682),
            .I(N__19679));
    Span4Mux_v I__1862 (
            .O(N__19679),
            .I(N__19676));
    Odrv4 I__1861 (
            .O(N__19676),
            .I(alt_ki_1));
    InMux I__1860 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__1859 (
            .O(N__19670),
            .I(N__19667));
    Span4Mux_v I__1858 (
            .O(N__19667),
            .I(N__19664));
    Odrv4 I__1857 (
            .O(N__19664),
            .I(alt_ki_2));
    InMux I__1856 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__1855 (
            .O(N__19658),
            .I(N__19655));
    Span4Mux_s2_h I__1854 (
            .O(N__19655),
            .I(N__19652));
    Odrv4 I__1853 (
            .O(N__19652),
            .I(alt_ki_3));
    InMux I__1852 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__1851 (
            .O(N__19646),
            .I(\pid_alt.O_3_9 ));
    InMux I__1850 (
            .O(N__19643),
            .I(N__19640));
    LocalMux I__1849 (
            .O(N__19640),
            .I(\pid_alt.O_3_10 ));
    InMux I__1848 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__1847 (
            .O(N__19634),
            .I(\pid_alt.O_3_11 ));
    InMux I__1846 (
            .O(N__19631),
            .I(N__19628));
    LocalMux I__1845 (
            .O(N__19628),
            .I(\pid_alt.O_3_13 ));
    InMux I__1844 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__1843 (
            .O(N__19622),
            .I(N__19619));
    Span4Mux_v I__1842 (
            .O(N__19619),
            .I(N__19616));
    Odrv4 I__1841 (
            .O(N__19616),
            .I(\pid_alt.O_1_8 ));
    InMux I__1840 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__1839 (
            .O(N__19610),
            .I(N__19607));
    Span4Mux_h I__1838 (
            .O(N__19607),
            .I(N__19604));
    Odrv4 I__1837 (
            .O(N__19604),
            .I(\pid_alt.O_1_11 ));
    InMux I__1836 (
            .O(N__19601),
            .I(N__19598));
    LocalMux I__1835 (
            .O(N__19598),
            .I(N__19595));
    Odrv4 I__1834 (
            .O(N__19595),
            .I(alt_kd_6));
    InMux I__1833 (
            .O(N__19592),
            .I(N__19589));
    LocalMux I__1832 (
            .O(N__19589),
            .I(N__19586));
    Odrv4 I__1831 (
            .O(N__19586),
            .I(alt_kd_2));
    InMux I__1830 (
            .O(N__19583),
            .I(N__19580));
    LocalMux I__1829 (
            .O(N__19580),
            .I(N__19577));
    Span4Mux_s2_h I__1828 (
            .O(N__19577),
            .I(N__19574));
    Odrv4 I__1827 (
            .O(N__19574),
            .I(alt_kd_7));
    InMux I__1826 (
            .O(N__19571),
            .I(N__19568));
    LocalMux I__1825 (
            .O(N__19568),
            .I(N__19565));
    Span4Mux_h I__1824 (
            .O(N__19565),
            .I(N__19562));
    Odrv4 I__1823 (
            .O(N__19562),
            .I(\pid_alt.O_3_24 ));
    InMux I__1822 (
            .O(N__19559),
            .I(N__19556));
    LocalMux I__1821 (
            .O(N__19556),
            .I(N__19553));
    Odrv4 I__1820 (
            .O(N__19553),
            .I(\pid_alt.O_3_20 ));
    InMux I__1819 (
            .O(N__19550),
            .I(N__19547));
    LocalMux I__1818 (
            .O(N__19547),
            .I(N__19544));
    Odrv4 I__1817 (
            .O(N__19544),
            .I(\pid_alt.O_3_21 ));
    InMux I__1816 (
            .O(N__19541),
            .I(N__19538));
    LocalMux I__1815 (
            .O(N__19538),
            .I(N__19535));
    Odrv4 I__1814 (
            .O(N__19535),
            .I(\pid_alt.O_3_22 ));
    InMux I__1813 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__1812 (
            .O(N__19529),
            .I(N__19526));
    Odrv4 I__1811 (
            .O(N__19526),
            .I(\pid_alt.O_3_23 ));
    InMux I__1810 (
            .O(N__19523),
            .I(N__19520));
    LocalMux I__1809 (
            .O(N__19520),
            .I(N__19517));
    Odrv4 I__1808 (
            .O(N__19517),
            .I(\pid_alt.O_3_15 ));
    InMux I__1807 (
            .O(N__19514),
            .I(N__19511));
    LocalMux I__1806 (
            .O(N__19511),
            .I(N__19508));
    Odrv4 I__1805 (
            .O(N__19508),
            .I(\pid_alt.O_3_19 ));
    InMux I__1804 (
            .O(N__19505),
            .I(N__19502));
    LocalMux I__1803 (
            .O(N__19502),
            .I(\pid_alt.O_3_14 ));
    InMux I__1802 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1801 (
            .O(N__19496),
            .I(\pid_alt.O_3_8 ));
    InMux I__1800 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__1799 (
            .O(N__19490),
            .I(N__19487));
    Odrv4 I__1798 (
            .O(N__19487),
            .I(\pid_alt.O_3_6 ));
    CascadeMux I__1797 (
            .O(N__19484),
            .I(N__19480));
    InMux I__1796 (
            .O(N__19483),
            .I(N__19476));
    InMux I__1795 (
            .O(N__19480),
            .I(N__19469));
    InMux I__1794 (
            .O(N__19479),
            .I(N__19469));
    LocalMux I__1793 (
            .O(N__19476),
            .I(N__19466));
    InMux I__1792 (
            .O(N__19475),
            .I(N__19461));
    InMux I__1791 (
            .O(N__19474),
            .I(N__19461));
    LocalMux I__1790 (
            .O(N__19469),
            .I(N__19458));
    Span4Mux_v I__1789 (
            .O(N__19466),
            .I(N__19453));
    LocalMux I__1788 (
            .O(N__19461),
            .I(N__19453));
    Odrv4 I__1787 (
            .O(N__19458),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    Odrv4 I__1786 (
            .O(N__19453),
            .I(\pid_alt.error_p_regZ0Z_2 ));
    InMux I__1785 (
            .O(N__19448),
            .I(N__19445));
    LocalMux I__1784 (
            .O(N__19445),
            .I(\pid_alt.O_3_7 ));
    InMux I__1783 (
            .O(N__19442),
            .I(N__19438));
    InMux I__1782 (
            .O(N__19441),
            .I(N__19434));
    LocalMux I__1781 (
            .O(N__19438),
            .I(N__19431));
    InMux I__1780 (
            .O(N__19437),
            .I(N__19428));
    LocalMux I__1779 (
            .O(N__19434),
            .I(N__19425));
    Span4Mux_v I__1778 (
            .O(N__19431),
            .I(N__19420));
    LocalMux I__1777 (
            .O(N__19428),
            .I(N__19420));
    Odrv12 I__1776 (
            .O(N__19425),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    Odrv4 I__1775 (
            .O(N__19420),
            .I(\pid_alt.error_p_regZ0Z_3 ));
    InMux I__1774 (
            .O(N__19415),
            .I(N__19412));
    LocalMux I__1773 (
            .O(N__19412),
            .I(\pid_alt.O_3_5 ));
    InMux I__1772 (
            .O(N__19409),
            .I(N__19399));
    InMux I__1771 (
            .O(N__19408),
            .I(N__19399));
    InMux I__1770 (
            .O(N__19407),
            .I(N__19394));
    InMux I__1769 (
            .O(N__19406),
            .I(N__19394));
    InMux I__1768 (
            .O(N__19405),
            .I(N__19389));
    InMux I__1767 (
            .O(N__19404),
            .I(N__19389));
    LocalMux I__1766 (
            .O(N__19399),
            .I(N__19382));
    LocalMux I__1765 (
            .O(N__19394),
            .I(N__19382));
    LocalMux I__1764 (
            .O(N__19389),
            .I(N__19382));
    Odrv12 I__1763 (
            .O(N__19382),
            .I(\pid_alt.error_p_regZ0Z_1 ));
    InMux I__1762 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__1761 (
            .O(N__19376),
            .I(N__19373));
    Odrv4 I__1760 (
            .O(N__19373),
            .I(\pid_alt.O_3_12 ));
    InMux I__1759 (
            .O(N__19370),
            .I(N__19367));
    LocalMux I__1758 (
            .O(N__19367),
            .I(N__19364));
    Odrv4 I__1757 (
            .O(N__19364),
            .I(\pid_alt.O_3_16 ));
    InMux I__1756 (
            .O(N__19361),
            .I(N__19358));
    LocalMux I__1755 (
            .O(N__19358),
            .I(N__19355));
    Odrv4 I__1754 (
            .O(N__19355),
            .I(\pid_alt.O_3_17 ));
    InMux I__1753 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__1752 (
            .O(N__19349),
            .I(N__19346));
    Odrv4 I__1751 (
            .O(N__19346),
            .I(\pid_alt.O_3_18 ));
    InMux I__1750 (
            .O(N__19343),
            .I(N__19340));
    LocalMux I__1749 (
            .O(N__19340),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ));
    CascadeMux I__1748 (
            .O(N__19337),
            .I(N__19332));
    InMux I__1747 (
            .O(N__19336),
            .I(N__19324));
    InMux I__1746 (
            .O(N__19335),
            .I(N__19324));
    InMux I__1745 (
            .O(N__19332),
            .I(N__19319));
    InMux I__1744 (
            .O(N__19331),
            .I(N__19319));
    InMux I__1743 (
            .O(N__19330),
            .I(N__19314));
    InMux I__1742 (
            .O(N__19329),
            .I(N__19314));
    LocalMux I__1741 (
            .O(N__19324),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__1740 (
            .O(N__19319),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    LocalMux I__1739 (
            .O(N__19314),
            .I(\pid_alt.error_d_reg_prevZ0Z_1 ));
    InMux I__1738 (
            .O(N__19307),
            .I(N__19296));
    InMux I__1737 (
            .O(N__19306),
            .I(N__19296));
    InMux I__1736 (
            .O(N__19305),
            .I(N__19289));
    InMux I__1735 (
            .O(N__19304),
            .I(N__19289));
    InMux I__1734 (
            .O(N__19303),
            .I(N__19289));
    InMux I__1733 (
            .O(N__19302),
            .I(N__19284));
    InMux I__1732 (
            .O(N__19301),
            .I(N__19284));
    LocalMux I__1731 (
            .O(N__19296),
            .I(N__19277));
    LocalMux I__1730 (
            .O(N__19289),
            .I(N__19277));
    LocalMux I__1729 (
            .O(N__19284),
            .I(N__19277));
    Odrv12 I__1728 (
            .O(N__19277),
            .I(\pid_alt.error_d_regZ0Z_1 ));
    InMux I__1727 (
            .O(N__19274),
            .I(N__19271));
    LocalMux I__1726 (
            .O(N__19271),
            .I(\pid_alt.N_3_1 ));
    InMux I__1725 (
            .O(N__19268),
            .I(N__19265));
    LocalMux I__1724 (
            .O(N__19265),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ));
    InMux I__1723 (
            .O(N__19262),
            .I(N__19254));
    InMux I__1722 (
            .O(N__19261),
            .I(N__19249));
    InMux I__1721 (
            .O(N__19260),
            .I(N__19249));
    InMux I__1720 (
            .O(N__19259),
            .I(N__19242));
    InMux I__1719 (
            .O(N__19258),
            .I(N__19242));
    InMux I__1718 (
            .O(N__19257),
            .I(N__19242));
    LocalMux I__1717 (
            .O(N__19254),
            .I(N__19235));
    LocalMux I__1716 (
            .O(N__19249),
            .I(N__19235));
    LocalMux I__1715 (
            .O(N__19242),
            .I(N__19235));
    Odrv12 I__1714 (
            .O(N__19235),
            .I(\pid_alt.error_d_regZ0Z_2 ));
    InMux I__1713 (
            .O(N__19232),
            .I(N__19229));
    LocalMux I__1712 (
            .O(N__19229),
            .I(N__19222));
    InMux I__1711 (
            .O(N__19228),
            .I(N__19217));
    InMux I__1710 (
            .O(N__19227),
            .I(N__19217));
    InMux I__1709 (
            .O(N__19226),
            .I(N__19212));
    InMux I__1708 (
            .O(N__19225),
            .I(N__19212));
    Odrv4 I__1707 (
            .O(N__19222),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__1706 (
            .O(N__19217),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    LocalMux I__1705 (
            .O(N__19212),
            .I(\pid_alt.error_d_reg_prevZ0Z_2 ));
    InMux I__1704 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__1703 (
            .O(N__19202),
            .I(N__19199));
    Odrv4 I__1702 (
            .O(N__19199),
            .I(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ));
    InMux I__1701 (
            .O(N__19196),
            .I(N__19193));
    LocalMux I__1700 (
            .O(N__19193),
            .I(N__19190));
    Span4Mux_v I__1699 (
            .O(N__19190),
            .I(N__19185));
    InMux I__1698 (
            .O(N__19189),
            .I(N__19180));
    InMux I__1697 (
            .O(N__19188),
            .I(N__19180));
    Odrv4 I__1696 (
            .O(N__19185),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    LocalMux I__1695 (
            .O(N__19180),
            .I(\pid_alt.error_d_reg_prevZ0Z_3 ));
    InMux I__1694 (
            .O(N__19175),
            .I(N__19165));
    InMux I__1693 (
            .O(N__19174),
            .I(N__19165));
    InMux I__1692 (
            .O(N__19173),
            .I(N__19165));
    InMux I__1691 (
            .O(N__19172),
            .I(N__19162));
    LocalMux I__1690 (
            .O(N__19165),
            .I(N__19159));
    LocalMux I__1689 (
            .O(N__19162),
            .I(N__19154));
    Span12Mux_v I__1688 (
            .O(N__19159),
            .I(N__19154));
    Odrv12 I__1687 (
            .O(N__19154),
            .I(\pid_alt.error_d_regZ0Z_3 ));
    InMux I__1686 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__1685 (
            .O(N__19148),
            .I(N__19145));
    Odrv4 I__1684 (
            .O(N__19145),
            .I(\pid_alt.g0_4_0 ));
    InMux I__1683 (
            .O(N__19142),
            .I(N__19139));
    LocalMux I__1682 (
            .O(N__19139),
            .I(\pid_alt.N_1505_i_0 ));
    InMux I__1681 (
            .O(N__19136),
            .I(N__19133));
    LocalMux I__1680 (
            .O(N__19133),
            .I(\pid_alt.N_3_0 ));
    CascadeMux I__1679 (
            .O(N__19130),
            .I(N__19127));
    InMux I__1678 (
            .O(N__19127),
            .I(N__19124));
    LocalMux I__1677 (
            .O(N__19124),
            .I(\pid_alt.N_1507_0 ));
    InMux I__1676 (
            .O(N__19121),
            .I(N__19118));
    LocalMux I__1675 (
            .O(N__19118),
            .I(\pid_alt.N_5 ));
    InMux I__1674 (
            .O(N__19115),
            .I(N__19112));
    LocalMux I__1673 (
            .O(N__19112),
            .I(\pid_alt.N_1511_0 ));
    CascadeMux I__1672 (
            .O(N__19109),
            .I(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ));
    InMux I__1671 (
            .O(N__19106),
            .I(N__19102));
    InMux I__1670 (
            .O(N__19105),
            .I(N__19097));
    LocalMux I__1669 (
            .O(N__19102),
            .I(N__19094));
    InMux I__1668 (
            .O(N__19101),
            .I(N__19089));
    InMux I__1667 (
            .O(N__19100),
            .I(N__19089));
    LocalMux I__1666 (
            .O(N__19097),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    Odrv4 I__1665 (
            .O(N__19094),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    LocalMux I__1664 (
            .O(N__19089),
            .I(\pid_alt.error_p_regZ0Z_0 ));
    InMux I__1663 (
            .O(N__19082),
            .I(N__19079));
    LocalMux I__1662 (
            .O(N__19079),
            .I(\pid_alt.N_1505_i_1 ));
    CascadeMux I__1661 (
            .O(N__19076),
            .I(N__19073));
    InMux I__1660 (
            .O(N__19073),
            .I(N__19070));
    LocalMux I__1659 (
            .O(N__19070),
            .I(\pid_alt.N_1507_1 ));
    CascadeMux I__1658 (
            .O(N__19067),
            .I(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ));
    InMux I__1657 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__1656 (
            .O(N__19061),
            .I(N__19058));
    Span12Mux_s4_h I__1655 (
            .O(N__19058),
            .I(N__19055));
    Span12Mux_v I__1654 (
            .O(N__19055),
            .I(N__19052));
    Odrv12 I__1653 (
            .O(N__19052),
            .I(\pid_alt.O_1_4 ));
    InMux I__1652 (
            .O(N__19049),
            .I(N__19046));
    LocalMux I__1651 (
            .O(N__19046),
            .I(N__19043));
    Span4Mux_v I__1650 (
            .O(N__19043),
            .I(N__19040));
    Span4Mux_s1_h I__1649 (
            .O(N__19040),
            .I(N__19037));
    Odrv4 I__1648 (
            .O(N__19037),
            .I(\pid_alt.O_3_4 ));
    CascadeMux I__1647 (
            .O(N__19034),
            .I(N__19031));
    InMux I__1646 (
            .O(N__19031),
            .I(N__19028));
    LocalMux I__1645 (
            .O(N__19028),
            .I(\pid_alt.N_1505_i ));
    CascadeMux I__1644 (
            .O(N__19025),
            .I(\pid_alt.N_1505_i_cascade_ ));
    InMux I__1643 (
            .O(N__19022),
            .I(N__19019));
    LocalMux I__1642 (
            .O(N__19019),
            .I(\pid_alt.un1_pid_prereg_0_axb_2_1 ));
    CascadeMux I__1641 (
            .O(N__19016),
            .I(\pid_alt.N_1513_0_cascade_ ));
    InMux I__1640 (
            .O(N__19013),
            .I(N__19010));
    LocalMux I__1639 (
            .O(N__19010),
            .I(\pid_side.O_0_11 ));
    InMux I__1638 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__1637 (
            .O(N__19004),
            .I(\pid_side.O_0_6 ));
    InMux I__1636 (
            .O(N__19001),
            .I(N__18998));
    LocalMux I__1635 (
            .O(N__18998),
            .I(\pid_side.O_0_17 ));
    InMux I__1634 (
            .O(N__18995),
            .I(N__18992));
    LocalMux I__1633 (
            .O(N__18992),
            .I(\pid_side.O_0_16 ));
    InMux I__1632 (
            .O(N__18989),
            .I(N__18986));
    LocalMux I__1631 (
            .O(N__18986),
            .I(\pid_side.O_0_12 ));
    InMux I__1630 (
            .O(N__18983),
            .I(N__18980));
    LocalMux I__1629 (
            .O(N__18980),
            .I(\pid_side.O_0_20 ));
    InMux I__1628 (
            .O(N__18977),
            .I(N__18974));
    LocalMux I__1627 (
            .O(N__18974),
            .I(\pid_side.O_0_21 ));
    InMux I__1626 (
            .O(N__18971),
            .I(N__18968));
    LocalMux I__1625 (
            .O(N__18968),
            .I(\pid_side.O_0_22 ));
    InMux I__1624 (
            .O(N__18965),
            .I(N__18962));
    LocalMux I__1623 (
            .O(N__18962),
            .I(\pid_side.O_0_9 ));
    InMux I__1622 (
            .O(N__18959),
            .I(N__18956));
    LocalMux I__1621 (
            .O(N__18956),
            .I(N__18953));
    Odrv4 I__1620 (
            .O(N__18953),
            .I(\pid_side.O_0_19 ));
    InMux I__1619 (
            .O(N__18950),
            .I(N__18947));
    LocalMux I__1618 (
            .O(N__18947),
            .I(\pid_side.O_0_14 ));
    InMux I__1617 (
            .O(N__18944),
            .I(N__18941));
    LocalMux I__1616 (
            .O(N__18941),
            .I(\pid_side.O_0_8 ));
    InMux I__1615 (
            .O(N__18938),
            .I(N__18935));
    LocalMux I__1614 (
            .O(N__18935),
            .I(\pid_side.O_0_10 ));
    InMux I__1613 (
            .O(N__18932),
            .I(N__18929));
    LocalMux I__1612 (
            .O(N__18929),
            .I(N__18926));
    Odrv4 I__1611 (
            .O(N__18926),
            .I(\pid_side.O_0_23 ));
    InMux I__1610 (
            .O(N__18923),
            .I(N__18920));
    LocalMux I__1609 (
            .O(N__18920),
            .I(N__18917));
    Odrv4 I__1608 (
            .O(N__18917),
            .I(\pid_side.O_0_15 ));
    InMux I__1607 (
            .O(N__18914),
            .I(N__18911));
    LocalMux I__1606 (
            .O(N__18911),
            .I(N__18908));
    Odrv4 I__1605 (
            .O(N__18908),
            .I(\pid_side.O_0_18 ));
    InMux I__1604 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__1603 (
            .O(N__18902),
            .I(\pid_alt.O_2_17 ));
    InMux I__1602 (
            .O(N__18899),
            .I(N__18896));
    LocalMux I__1601 (
            .O(N__18896),
            .I(N__18893));
    Span4Mux_v I__1600 (
            .O(N__18893),
            .I(N__18890));
    Odrv4 I__1599 (
            .O(N__18890),
            .I(\pid_alt.O_1_6 ));
    InMux I__1598 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__1597 (
            .O(N__18884),
            .I(\pid_alt.O_2_12 ));
    InMux I__1596 (
            .O(N__18881),
            .I(N__18878));
    LocalMux I__1595 (
            .O(N__18878),
            .I(\pid_alt.O_2_19 ));
    InMux I__1594 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__1593 (
            .O(N__18872),
            .I(\pid_alt.O_2_14 ));
    InMux I__1592 (
            .O(N__18869),
            .I(N__18866));
    LocalMux I__1591 (
            .O(N__18866),
            .I(\pid_alt.O_2_15 ));
    InMux I__1590 (
            .O(N__18863),
            .I(N__18860));
    LocalMux I__1589 (
            .O(N__18860),
            .I(N__18857));
    Span4Mux_h I__1588 (
            .O(N__18857),
            .I(N__18854));
    Span4Mux_v I__1587 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__1586 (
            .O(N__18851),
            .I(\pid_alt.O_1_5 ));
    InMux I__1585 (
            .O(N__18848),
            .I(N__18845));
    LocalMux I__1584 (
            .O(N__18845),
            .I(N__18842));
    Span4Mux_h I__1583 (
            .O(N__18842),
            .I(N__18839));
    Odrv4 I__1582 (
            .O(N__18839),
            .I(\pid_alt.O_2_22 ));
    InMux I__1581 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__1580 (
            .O(N__18833),
            .I(\pid_alt.O_2_11 ));
    InMux I__1579 (
            .O(N__18830),
            .I(N__18827));
    LocalMux I__1578 (
            .O(N__18827),
            .I(N__18824));
    Odrv4 I__1577 (
            .O(N__18824),
            .I(\pid_alt.O_2_24 ));
    InMux I__1576 (
            .O(N__18821),
            .I(N__18818));
    LocalMux I__1575 (
            .O(N__18818),
            .I(\pid_alt.O_2_7 ));
    InMux I__1574 (
            .O(N__18815),
            .I(N__18812));
    LocalMux I__1573 (
            .O(N__18812),
            .I(\pid_alt.O_2_8 ));
    InMux I__1572 (
            .O(N__18809),
            .I(N__18806));
    LocalMux I__1571 (
            .O(N__18806),
            .I(N__18803));
    Odrv4 I__1570 (
            .O(N__18803),
            .I(\pid_alt.O_2_23 ));
    InMux I__1569 (
            .O(N__18800),
            .I(N__18797));
    LocalMux I__1568 (
            .O(N__18797),
            .I(\pid_alt.O_2_10 ));
    InMux I__1567 (
            .O(N__18794),
            .I(N__18791));
    LocalMux I__1566 (
            .O(N__18791),
            .I(\pid_alt.O_2_9 ));
    InMux I__1565 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__1564 (
            .O(N__18785),
            .I(N__18782));
    Odrv4 I__1563 (
            .O(N__18782),
            .I(\pid_alt.O_2_16 ));
    InMux I__1562 (
            .O(N__18779),
            .I(N__18776));
    LocalMux I__1561 (
            .O(N__18776),
            .I(N__18773));
    Odrv4 I__1560 (
            .O(N__18773),
            .I(\pid_alt.O_1_24 ));
    InMux I__1559 (
            .O(N__18770),
            .I(N__18767));
    LocalMux I__1558 (
            .O(N__18767),
            .I(\pid_alt.O_1_13 ));
    InMux I__1557 (
            .O(N__18764),
            .I(N__18761));
    LocalMux I__1556 (
            .O(N__18761),
            .I(\pid_alt.O_1_14 ));
    InMux I__1555 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__1554 (
            .O(N__18755),
            .I(\pid_alt.O_1_10 ));
    InMux I__1553 (
            .O(N__18752),
            .I(N__18749));
    LocalMux I__1552 (
            .O(N__18749),
            .I(\pid_alt.O_1_21 ));
    InMux I__1551 (
            .O(N__18746),
            .I(N__18743));
    LocalMux I__1550 (
            .O(N__18743),
            .I(N__18740));
    Odrv4 I__1549 (
            .O(N__18740),
            .I(\pid_alt.O_2_13 ));
    InMux I__1548 (
            .O(N__18737),
            .I(N__18734));
    LocalMux I__1547 (
            .O(N__18734),
            .I(N__18731));
    Odrv4 I__1546 (
            .O(N__18731),
            .I(\pid_alt.O_2_21 ));
    InMux I__1545 (
            .O(N__18728),
            .I(N__18725));
    LocalMux I__1544 (
            .O(N__18725),
            .I(N__18722));
    Odrv4 I__1543 (
            .O(N__18722),
            .I(\pid_alt.O_2_18 ));
    InMux I__1542 (
            .O(N__18719),
            .I(N__18716));
    LocalMux I__1541 (
            .O(N__18716),
            .I(N__18713));
    Odrv4 I__1540 (
            .O(N__18713),
            .I(\pid_alt.O_2_20 ));
    InMux I__1539 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1538 (
            .O(N__18707),
            .I(\pid_alt.O_1_15 ));
    InMux I__1537 (
            .O(N__18704),
            .I(N__18701));
    LocalMux I__1536 (
            .O(N__18701),
            .I(N__18698));
    Odrv4 I__1535 (
            .O(N__18698),
            .I(\pid_alt.O_1_16 ));
    InMux I__1534 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__1533 (
            .O(N__18692),
            .I(N__18689));
    Odrv4 I__1532 (
            .O(N__18689),
            .I(\pid_alt.O_1_17 ));
    InMux I__1531 (
            .O(N__18686),
            .I(N__18683));
    LocalMux I__1530 (
            .O(N__18683),
            .I(N__18680));
    Odrv4 I__1529 (
            .O(N__18680),
            .I(\pid_alt.O_1_19 ));
    InMux I__1528 (
            .O(N__18677),
            .I(N__18674));
    LocalMux I__1527 (
            .O(N__18674),
            .I(N__18671));
    Odrv4 I__1526 (
            .O(N__18671),
            .I(\pid_alt.O_1_20 ));
    InMux I__1525 (
            .O(N__18668),
            .I(N__18665));
    LocalMux I__1524 (
            .O(N__18665),
            .I(\pid_alt.O_1_7 ));
    InMux I__1523 (
            .O(N__18662),
            .I(N__18659));
    LocalMux I__1522 (
            .O(N__18659),
            .I(\pid_alt.O_1_22 ));
    InMux I__1521 (
            .O(N__18656),
            .I(N__18653));
    LocalMux I__1520 (
            .O(N__18653),
            .I(\pid_alt.O_1_23 ));
    InMux I__1519 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__1518 (
            .O(N__18647),
            .I(\pid_alt.O_1_18 ));
    InMux I__1517 (
            .O(N__18644),
            .I(N__18641));
    LocalMux I__1516 (
            .O(N__18641),
            .I(\pid_alt.O_1_12 ));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\scaler_4.un3_source_data_0_cry_7 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\scaler_4.un2_source_data_0_cry_8 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\reset_module_System.count_1_cry_8 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\reset_module_System.count_1_cry_16 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(\ppm_encoder_1.un1_throttle_cry_7 ),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\ppm_encoder_1.un1_rudder_cry_13 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\ppm_encoder_1.un1_elevator_cry_7 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\ppm_encoder_1.un1_aileron_cry_7 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_cry_8 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\pid_side.un1_pid_prereg_cry_16 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_cry_8 ),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\pid_front.un1_pid_prereg_cry_16 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\pid_alt.error_cry_7 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_4_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_21_0_));
    defparam IN_MUX_bfv_4_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_22_0_ (
            .carryinitin(\pid_side.error_cry_3_0 ),
            .carryinitout(bfn_4_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(\pid_front.error_cry_3_0 ),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .carryinitout(bfn_8_8_0_));
    ICE_GB \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0  (
            .USERSIGNALTOGLOBALBUFFER(N__42143),
            .GLOBALBUFFEROUTPUT(\ppm_encoder_1.N_661_g ));
    ICE_GB \pid_alt.state_RNICP2N1_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__25910),
            .GLOBALBUFFEROUTPUT(\pid_alt.N_850_0_g ));
    ICE_GB \reset_module_System.reset_RNITC69_0  (
            .USERSIGNALTOGLOBALBUFFER(N__48314),
            .GLOBALBUFFEROUTPUT(N_851_g));
    ICE_GB \reset_module_System.reset_RNITC69  (
            .USERSIGNALTOGLOBALBUFFER(N__49034),
            .GLOBALBUFFEROUTPUT(reset_system_g));
    ICE_GB \pid_alt.state_RNIH1EN_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__31118),
            .GLOBALBUFFEROUTPUT(\pid_alt.state_0_g_0 ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_8_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_8_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18644),
            .lcout(\pid_alt.error_d_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_11_LC_1_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_11_LC_1_5_2  (
            .in0(N__18710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_12_LC_1_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_12_LC_1_5_3  (
            .in0(N__18704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_13_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_13_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18695),
            .lcout(\pid_alt.error_d_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_15_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_15_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18686),
            .lcout(\pid_alt.error_d_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_16_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_16_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18677),
            .lcout(\pid_alt.error_d_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51542),
            .ce(N__20330),
            .sr(N__50717));
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_3_LC_1_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_esr_3_LC_1_6_0  (
            .in0(N__18668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_18_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_18_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18662),
            .lcout(\pid_alt.error_d_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_19_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_19_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18656),
            .lcout(\pid_alt.error_d_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_14_LC_1_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_14_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18650),
            .lcout(\pid_alt.error_d_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_20_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_20_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18779),
            .lcout(\pid_alt.error_d_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_9_LC_1_6_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_9_LC_1_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_9_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18770),
            .lcout(\pid_alt.error_d_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_10_LC_1_6_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_10_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_10_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18764),
            .lcout(\pid_alt.error_d_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_6_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_6_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18758),
            .lcout(\pid_alt.error_d_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51540),
            .ce(N__20328),
            .sr(N__50715));
    defparam \pid_alt.error_d_reg_esr_17_LC_1_7_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_7_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_17_LC_1_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_17_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18752),
            .lcout(\pid_alt.error_d_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51537),
            .ce(N__20327),
            .sr(N__50714));
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_9_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_9_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18746),
            .lcout(\pid_alt.error_i_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51531),
            .ce(N__20325),
            .sr(N__50712));
    defparam \pid_alt.error_i_reg_esr_17_LC_1_9_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_17_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_17_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18737),
            .lcout(\pid_alt.error_i_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51531),
            .ce(N__20325),
            .sr(N__50712));
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_14_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_14_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18728),
            .lcout(\pid_alt.error_i_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51531),
            .ce(N__20325),
            .sr(N__50712));
    defparam \pid_alt.error_i_reg_esr_16_LC_1_9_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_16_LC_1_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_16_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18719),
            .lcout(\pid_alt.error_i_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51531),
            .ce(N__20325),
            .sr(N__50712));
    defparam \pid_alt.error_i_reg_esr_18_LC_1_9_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_18_LC_1_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_18_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(\pid_alt.error_i_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51531),
            .ce(N__20325),
            .sr(N__50712));
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_7_LC_1_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_7_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18836),
            .lcout(\pid_alt.error_i_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_20_LC_1_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_20_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18830),
            .lcout(\pid_alt.error_i_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_3_LC_1_10_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_3_LC_1_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_3_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18821),
            .lcout(\pid_alt.error_i_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_4_LC_1_10_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_4_LC_1_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_4_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18815),
            .lcout(\pid_alt.error_i_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_19_LC_1_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_19_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18809),
            .lcout(\pid_alt.error_i_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_6_LC_1_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_6_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18800),
            .lcout(\pid_alt.error_i_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_5_LC_1_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_5_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18794),
            .lcout(\pid_alt.error_i_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_12_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_12_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18788),
            .lcout(\pid_alt.error_i_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51527),
            .ce(N__20324),
            .sr(N__50711));
    defparam \pid_alt.error_i_reg_esr_13_LC_1_11_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_13_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_13_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18905),
            .lcout(\pid_alt.error_i_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_2_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_2_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18899),
            .lcout(\pid_alt.error_d_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_8_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_8_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18887),
            .lcout(\pid_alt.error_i_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_15_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_15_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18881),
            .lcout(\pid_alt.error_i_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_i_reg_esr_10_LC_1_11_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_10_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_10_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18875),
            .lcout(\pid_alt.error_i_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_11_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_11_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18869),
            .lcout(\pid_alt.error_i_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51522),
            .ce(N__20323),
            .sr(N__50710));
    defparam \pid_alt.error_d_reg_esr_1_LC_1_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_1_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_1_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18863),
            .lcout(\pid_alt.error_d_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51517),
            .ce(N__20321),
            .sr(N__50708));
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_1_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_13_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_13_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22259),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51511),
            .ce(N__25564),
            .sr(N__49537));
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_4_LC_1_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_4_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19811),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51511),
            .ce(N__25564),
            .sr(N__49537));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_1_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_1_14_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_1_14_1  (
            .in0(N__19441),
            .in1(N__19196),
            .in2(_gnd_net_),
            .in3(N__19172),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_6  (
            .in0(N__22301),
            .in1(N__22273),
            .in2(_gnd_net_),
            .in3(N__22258),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_5_LC_1_15_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_5_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_5_LC_1_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_5_LC_1_15_0  (
            .in0(N__50204),
            .in1(N__30853),
            .in2(_gnd_net_),
            .in3(N__18965),
            .lcout(\pid_side.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_15_LC_1_15_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_15_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_15_LC_1_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_side.error_p_reg_15_LC_1_15_1  (
            .in0(N__18959),
            .in1(N__50206),
            .in2(_gnd_net_),
            .in3(N__28260),
            .lcout(\pid_side.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_10_LC_1_15_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_10_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_10_LC_1_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_10_LC_1_15_2  (
            .in0(N__50202),
            .in1(N__29391),
            .in2(_gnd_net_),
            .in3(N__18950),
            .lcout(\pid_side.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_4_LC_1_15_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_4_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_4_LC_1_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_4_LC_1_15_3  (
            .in0(N__28368),
            .in1(N__50208),
            .in2(_gnd_net_),
            .in3(N__18944),
            .lcout(\pid_side.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_6_LC_1_15_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_6_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_6_LC_1_15_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \pid_side.error_p_reg_6_LC_1_15_4  (
            .in0(N__18938),
            .in1(_gnd_net_),
            .in2(N__50226),
            .in3(N__28336),
            .lcout(\pid_side.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_19_LC_1_15_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_19_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_19_LC_1_15_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_19_LC_1_15_5  (
            .in0(N__28293),
            .in1(N__50207),
            .in2(_gnd_net_),
            .in3(N__18932),
            .lcout(\pid_side.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_11_LC_1_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_11_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_11_LC_1_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_11_LC_1_15_6  (
            .in0(N__50203),
            .in1(N__28408),
            .in2(_gnd_net_),
            .in3(N__18923),
            .lcout(\pid_side.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_14_LC_1_15_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_14_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_14_LC_1_15_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_14_LC_1_15_7  (
            .in0(N__28219),
            .in1(N__50205),
            .in2(_gnd_net_),
            .in3(N__18914),
            .lcout(\pid_side.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51494),
            .ce(),
            .sr(N__50705));
    defparam \pid_side.error_p_reg_7_LC_1_16_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_7_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_7_LC_1_16_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_7_LC_1_16_0  (
            .in0(N__30354),
            .in1(N__50217),
            .in2(_gnd_net_),
            .in3(N__19013),
            .lcout(\pid_side.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_2_LC_1_16_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_2_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_2_LC_1_16_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \pid_side.error_p_reg_2_LC_1_16_1  (
            .in0(N__19007),
            .in1(_gnd_net_),
            .in2(N__50227),
            .in3(N__34701),
            .lcout(\pid_side.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_13_LC_1_16_2 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_13_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_13_LC_1_16_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_13_LC_1_16_2  (
            .in0(N__30825),
            .in1(N__50215),
            .in2(_gnd_net_),
            .in3(N__19001),
            .lcout(\pid_side.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_12_LC_1_16_3 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_12_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_12_LC_1_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_12_LC_1_16_3  (
            .in0(N__50212),
            .in1(N__28695),
            .in2(_gnd_net_),
            .in3(N__18995),
            .lcout(\pid_side.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_8_LC_1_16_4 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_8_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_8_LC_1_16_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_8_LC_1_16_4  (
            .in0(N__28438),
            .in1(N__50218),
            .in2(_gnd_net_),
            .in3(N__18989),
            .lcout(\pid_side.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_16_LC_1_16_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_16_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_16_LC_1_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_16_LC_1_16_5  (
            .in0(N__50213),
            .in1(N__30909),
            .in2(_gnd_net_),
            .in3(N__18983),
            .lcout(\pid_side.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_17_LC_1_16_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_17_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_17_LC_1_16_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_17_LC_1_16_6  (
            .in0(N__28176),
            .in1(N__50216),
            .in2(_gnd_net_),
            .in3(N__18977),
            .lcout(\pid_side.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_side.error_p_reg_18_LC_1_16_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_18_LC_1_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_18_LC_1_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_18_LC_1_16_7  (
            .in0(N__50214),
            .in1(N__28645),
            .in2(_gnd_net_),
            .in3(N__18971),
            .lcout(\pid_side.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51485),
            .ce(),
            .sr(N__50704));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_1_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_1_17_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_1_17_0  (
            .in0(N__19483),
            .in1(N__19232),
            .in2(_gnd_net_),
            .in3(N__19262),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_1_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_1_17_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__24182),
            .in2(N__19067),
            .in3(N__19022),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_17_2  (
            .in0(N__22577),
            .in1(N__19101),
            .in2(_gnd_net_),
            .in3(N__23705),
            .lcout(\pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_1_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_1_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_1_17_3  (
            .in0(N__19336),
            .in1(N__19409),
            .in2(N__19034),
            .in3(N__19307),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_0_LC_1_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_0_LC_1_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_0_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19064),
            .lcout(\pid_alt.error_d_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51472),
            .ce(N__20318),
            .sr(N__50703));
    defparam \pid_alt.error_p_reg_esr_0_LC_1_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_0_LC_1_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_0_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19049),
            .lcout(\pid_alt.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51472),
            .ce(N__20318),
            .sr(N__50703));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_17_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__19100),
            .in2(_gnd_net_),
            .in3(N__23704),
            .lcout(\pid_alt.N_1505_i ),
            .ltout(\pid_alt.N_1505_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_1_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_1_17_7 .LUT_INIT=16'b0010010010110010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_1_17_7  (
            .in0(N__19335),
            .in1(N__19408),
            .in2(N__19025),
            .in3(N__19306),
            .lcout(\pid_alt.un1_pid_prereg_0_axb_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_18_0 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_18_0  (
            .in0(N__19142),
            .in1(N__19121),
            .in2(N__19130),
            .in3(N__19136),
            .lcout(),
            .ltout(\pid_alt.N_1513_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_18_1 .LUT_INIT=16'b1110100011010100;
    LogicCell40 \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_18_1  (
            .in0(N__19151),
            .in1(N__19115),
            .in2(N__19016),
            .in3(N__19442),
            .lcout(\pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_18_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__19105),
            .in2(_gnd_net_),
            .in3(N__23709),
            .lcout(\pid_alt.N_1505_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_18_3  (
            .in0(N__19406),
            .in1(N__19331),
            .in2(_gnd_net_),
            .in3(N__19303),
            .lcout(\pid_alt.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_18_4 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_18_4  (
            .in0(N__19304),
            .in1(_gnd_net_),
            .in2(N__19337),
            .in3(N__19407),
            .lcout(\pid_alt.N_1507_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_18_5  (
            .in0(N__19227),
            .in1(N__19479),
            .in2(_gnd_net_),
            .in3(N__19260),
            .lcout(\pid_alt.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_18_6 .LUT_INIT=16'b1010000011111010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_18_6  (
            .in0(N__19261),
            .in1(_gnd_net_),
            .in2(N__19484),
            .in3(N__19228),
            .lcout(\pid_alt.N_1511_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_18_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_1_LC_1_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_1_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19305),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51459),
            .ce(N__25575),
            .sr(N__49579));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_19_0 .LUT_INIT=16'b0011000001110001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_19_0  (
            .in0(N__19082),
            .in1(N__19343),
            .in2(N__19076),
            .in3(N__19274),
            .lcout(),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_19_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_19_1  (
            .in0(N__24254),
            .in1(N__19205),
            .in2(N__19109),
            .in3(N__19268),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_19_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__19106),
            .in2(_gnd_net_),
            .in3(N__23713),
            .lcout(\pid_alt.N_1505_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_19_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_19_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_19_3  (
            .in0(N__19405),
            .in1(N__19330),
            .in2(_gnd_net_),
            .in3(N__19302),
            .lcout(\pid_alt.N_1507_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_19_4  (
            .in0(N__19474),
            .in1(N__19225),
            .in2(_gnd_net_),
            .in3(N__19257),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_19_5  (
            .in0(N__19404),
            .in1(N__19329),
            .in2(_gnd_net_),
            .in3(N__19301),
            .lcout(\pid_alt.N_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_19_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_19_6  (
            .in0(N__19475),
            .in1(N__19226),
            .in2(_gnd_net_),
            .in3(N__19258),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_19_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_2_LC_1_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_2_LC_1_19_7  (
            .in0(N__19259),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51442),
            .ce(N__25576),
            .sr(N__49587));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_20_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_20_0  (
            .in0(N__20968),
            .in1(N__20944),
            .in2(_gnd_net_),
            .in3(N__20925),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_1_20_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_1_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_17_LC_1_20_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_17_LC_1_20_1  (
            .in0(N__20926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51428),
            .ce(N__25577),
            .sr(N__49596));
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_1_20_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_1_20_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_1_20_2  (
            .in0(N__19437),
            .in1(N__19188),
            .in2(_gnd_net_),
            .in3(N__19173),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_1_20_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_3_LC_1_20_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_3_LC_1_20_3  (
            .in0(N__19175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51428),
            .ce(N__25577),
            .sr(N__49596));
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_1_20_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_1_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__19189),
            .in2(_gnd_net_),
            .in3(N__19174),
            .lcout(\pid_alt.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_5  (
            .in0(N__24337),
            .in1(N__24310),
            .in2(_gnd_net_),
            .in3(N__24291),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_8_LC_1_20_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_8_LC_1_20_6  (
            .in0(N__24292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51428),
            .ce(N__25577),
            .sr(N__49596));
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_2_LC_1_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_2_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19493),
            .lcout(\pid_alt.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51414),
            .ce(N__20317),
            .sr(N__50701));
    defparam \pid_alt.error_p_reg_esr_3_LC_1_22_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_3_LC_1_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_3_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19448),
            .lcout(\pid_alt.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_1_LC_1_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_1_LC_1_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_1_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19415),
            .lcout(\pid_alt.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_8_LC_1_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_8_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(\pid_alt.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_12_LC_1_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_12_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19370),
            .lcout(\pid_alt.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_13_LC_1_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_13_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19361),
            .lcout(\pid_alt.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_14_LC_1_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_14_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19352),
            .lcout(\pid_alt.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_20_LC_1_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_20_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19571),
            .lcout(\pid_alt.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51400),
            .ce(N__20316),
            .sr(N__50700));
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_16_LC_1_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_16_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19559),
            .lcout(\pid_alt.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_17_LC_1_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_17_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19550),
            .lcout(\pid_alt.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_18_LC_1_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_18_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19541),
            .lcout(\pid_alt.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_3 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_19_LC_1_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_19_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19532),
            .lcout(\pid_alt.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_11_LC_1_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_11_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19523),
            .lcout(\pid_alt.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_5 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_15_LC_1_23_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_p_reg_esr_15_LC_1_23_5  (
            .in0(N__19514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_6 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_10_LC_1_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_10_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19505),
            .lcout(\pid_alt.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_7 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_4_LC_1_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_4_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19499),
            .lcout(\pid_alt.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51385),
            .ce(N__20315),
            .sr(N__50699));
    defparam \pid_alt.error_p_reg_esr_5_LC_1_24_0 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_24_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_5_LC_1_24_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pid_alt.error_p_reg_esr_5_LC_1_24_0  (
            .in0(_gnd_net_),
            .in1(N__19649),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51374),
            .ce(N__20314),
            .sr(N__50698));
    defparam \pid_alt.error_p_reg_esr_6_LC_1_24_1 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_6_LC_1_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_6_LC_1_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19643),
            .lcout(\pid_alt.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51374),
            .ce(N__20314),
            .sr(N__50698));
    defparam \pid_alt.error_p_reg_esr_7_LC_1_24_2 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_24_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_7_LC_1_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_7_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19637),
            .lcout(\pid_alt.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51374),
            .ce(N__20314),
            .sr(N__50698));
    defparam \pid_alt.error_p_reg_esr_9_LC_1_24_4 .C_ON=1'b0;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_p_reg_esr_9_LC_1_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_p_reg_esr_9_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19631),
            .lcout(\pid_alt.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51374),
            .ce(N__20314),
            .sr(N__50698));
    defparam \pid_alt.error_d_reg_esr_4_LC_2_5_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_4_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_4_LC_2_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_4_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19625),
            .lcout(\pid_alt.error_d_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51541),
            .ce(N__20329),
            .sr(N__50716));
    defparam \pid_alt.error_d_reg_esr_7_LC_2_5_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_7_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_7_LC_2_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_7_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19613),
            .lcout(\pid_alt.error_d_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51541),
            .ce(N__20329),
            .sr(N__50716));
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_6_LC_2_6_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_6_LC_2_6_1  (
            .in0(N__50824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40110),
            .lcout(alt_kd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51538),
            .ce(N__21927),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_6_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_2_LC_2_6_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_2_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__39500),
            .in2(_gnd_net_),
            .in3(N__50823),
            .lcout(alt_kd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51538),
            .ce(N__21927),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_7_LC_2_6_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_7_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__40012),
            .in2(_gnd_net_),
            .in3(N__50825),
            .lcout(alt_kd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51538),
            .ce(N__21927),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_5_LC_2_7_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_5_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__40273),
            .in2(_gnd_net_),
            .in3(N__50819),
            .lcout(alt_kd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51535),
            .ce(N__21932),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_1_LC_2_7_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_1_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__39626),
            .in2(_gnd_net_),
            .in3(N__50818),
            .lcout(alt_kd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51535),
            .ce(N__21932),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_esr_5_LC_2_8_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_esr_5_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_esr_5_LC_2_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_esr_5_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19721),
            .lcout(\pid_alt.error_d_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51532),
            .ce(N__20326),
            .sr(N__50713));
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_0_LC_2_9_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_0_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__39749),
            .in2(_gnd_net_),
            .in3(N__50817),
            .lcout(alt_ki_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51528),
            .ce(N__38841),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_4_LC_2_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_4_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__40395),
            .in2(_gnd_net_),
            .in3(N__50815),
            .lcout(alt_ki_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51523),
            .ce(N__38832),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_2_10_2 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_2_10_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__25393),
            .in2(_gnd_net_),
            .in3(N__23509),
            .lcout(\scaler_4.un3_source_data_0_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_1_LC_2_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_1_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__39625),
            .in2(_gnd_net_),
            .in3(N__50812),
            .lcout(alt_ki_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51523),
            .ce(N__38832),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_2_LC_2_10_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_2_LC_2_10_5  (
            .in0(N__50813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39488),
            .lcout(alt_ki_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51523),
            .ce(N__38832),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_10_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_3_LC_2_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_3_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__39362),
            .in2(_gnd_net_),
            .in3(N__50814),
            .lcout(alt_ki_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51523),
            .ce(N__38832),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_5_LC_2_10_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_5_LC_2_10_7  (
            .in0(N__50816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40262),
            .lcout(alt_ki_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51523),
            .ce(N__38832),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_11_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_10_LC_2_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_10_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23889),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51518),
            .ce(N__25557),
            .sr(N__49518));
    defparam \pid_alt.error_i_reg_esr_1_LC_2_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_1_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_1_LC_2_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_1_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19769),
            .lcout(\pid_alt.error_i_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51512),
            .ce(N__20320),
            .sr(N__50707));
    defparam \pid_alt.error_i_reg_esr_0_LC_2_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_0_LC_2_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_0_LC_2_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_0_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19757),
            .lcout(\pid_alt.error_i_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51505),
            .ce(N__20319),
            .sr(N__50706));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HDV_8_LC_2_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HDV_8_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HDV_8_LC_2_14_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI8HDV_8_LC_2_14_0  (
            .in0(N__33313),
            .in1(N__20389),
            .in2(N__33377),
            .in3(N__20410),
            .lcout(\pid_alt.m39_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_2_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_8_LC_2_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_8_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24373),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51495),
            .ce(N__25565),
            .sr(N__49538));
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_2_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_9_LC_2_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_9_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20507),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51495),
            .ce(N__25565),
            .sr(N__49538));
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_2_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_13_LC_2_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_13_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22113),
            .lcout(\pid_alt.error_i_acumm7lto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51495),
            .ce(N__25565),
            .sr(N__49538));
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_21_LC_2_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_21_LC_2_14_4  (
            .in0(N__24731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51495),
            .ce(N__25565),
            .sr(N__49538));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_2_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_2_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_2_14_5  (
            .in0(N__24801),
            .in1(N__24762),
            .in2(_gnd_net_),
            .in3(N__24728),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_2_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_2_14_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_2_14_6  (
            .in0(N__24730),
            .in1(_gnd_net_),
            .in2(N__24767),
            .in3(N__24803),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_2_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_2_14_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_2_14_7  (
            .in0(N__24802),
            .in1(N__24763),
            .in2(_gnd_net_),
            .in3(N__24729),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_15_0  (
            .in0(N__19859),
            .in1(N__19852),
            .in2(N__22493),
            .in3(N__20694),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_15_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_15_1  (
            .in0(N__19840),
            .in1(N__19822),
            .in2(_gnd_net_),
            .in3(N__19806),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_15_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__19853),
            .in2(N__19844),
            .in3(N__20695),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_2_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_2_15_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_2_15_3  (
            .in0(N__23935),
            .in1(N__23914),
            .in2(_gnd_net_),
            .in3(N__23890),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_2_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_2_15_5 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_2_15_5  (
            .in0(N__19841),
            .in1(N__19823),
            .in2(_gnd_net_),
            .in3(N__19807),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FQN6_4_LC_2_15_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FQN6_4_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FQN6_4_LC_2_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1FQN6_4_LC_2_15_6  (
            .in0(N__22447),
            .in1(N__20122),
            .in2(N__19790),
            .in3(N__20664),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNILSTB3_4_LC_2_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNILSTB3_4_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNILSTB3_4_LC_2_15_7 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNILSTB3_4_LC_2_15_7  (
            .in0(N__20665),
            .in1(_gnd_net_),
            .in2(N__20126),
            .in3(N__19787),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_2_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_2_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_2_16_1  (
            .in0(N__19909),
            .in1(N__19918),
            .in2(_gnd_net_),
            .in3(N__19941),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_2_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_2_16_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__21004),
            .in2(N__19946),
            .in3(N__20986),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_2_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_9_LC_2_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_9_LC_2_16_4  (
            .in0(N__19943),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51473),
            .ce(N__25569),
            .sr(N__49550));
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_2_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_2_16_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_2_16_5  (
            .in0(N__19892),
            .in1(N__19886),
            .in2(_gnd_net_),
            .in3(N__20506),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_2_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_2_16_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_2_16_6  (
            .in0(N__19942),
            .in1(_gnd_net_),
            .in2(N__19922),
            .in3(N__19910),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_2_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_2_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_2_16_7  (
            .in0(N__24359),
            .in1(N__19885),
            .in2(N__19871),
            .in3(N__20505),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_17_0  (
            .in0(N__20044),
            .in1(N__19868),
            .in2(N__22858),
            .in3(N__25713),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_17_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_17_1  (
            .in0(N__19999),
            .in1(N__20008),
            .in2(_gnd_net_),
            .in3(N__20034),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_17_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_17_2  (
            .in0(N__20045),
            .in1(_gnd_net_),
            .in2(N__19862),
            .in3(N__25714),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_17_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_17_3  (
            .in0(N__24466),
            .in1(N__24890),
            .in2(_gnd_net_),
            .in3(N__24910),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_18_LC_2_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_18_LC_2_17_4  (
            .in0(N__20036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51461),
            .ce(N__25572),
            .sr(N__49560));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_17_5  (
            .in0(N__19985),
            .in1(N__19979),
            .in2(_gnd_net_),
            .in3(N__25684),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_17_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_17_6  (
            .in0(N__20035),
            .in1(_gnd_net_),
            .in2(N__20012),
            .in3(N__20000),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_2_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_2_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_2_17_7  (
            .in0(N__22885),
            .in1(N__19978),
            .in2(N__19967),
            .in3(N__25683),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIA5V86_5_LC_2_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIA5V86_5_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIA5V86_5_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIA5V86_5_LC_2_18_0  (
            .in0(N__19954),
            .in1(N__19964),
            .in2(N__22814),
            .in3(N__20617),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_18_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_18_1  (
            .in0(N__20110),
            .in1(N__20095),
            .in2(_gnd_net_),
            .in3(N__20085),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_18_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_18_2  (
            .in0(N__19955),
            .in1(_gnd_net_),
            .in2(N__19958),
            .in3(N__20618),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_18_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_18_3  (
            .in0(N__20168),
            .in1(N__20153),
            .in2(_gnd_net_),
            .in3(N__20143),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_5_LC_2_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_5_LC_2_18_4  (
            .in0(N__20144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51443),
            .ce(N__25573),
            .sr(N__49568));
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_18_5  (
            .in0(N__20167),
            .in1(N__20152),
            .in2(_gnd_net_),
            .in3(N__20142),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_6_LC_2_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_6_LC_2_18_6  (
            .in0(N__20087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51443),
            .ce(N__25573),
            .sr(N__49568));
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_18_7 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_18_7  (
            .in0(N__20111),
            .in1(N__20096),
            .in2(_gnd_net_),
            .in3(N__20086),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_20_LC_2_19_0 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_20_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_20_LC_2_19_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pid_side.error_p_reg_20_LC_2_19_0  (
            .in0(N__28137),
            .in1(_gnd_net_),
            .in2(N__50228),
            .in3(N__20069),
            .lcout(\pid_side.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51429),
            .ce(),
            .sr(N__50702));
    defparam \pid_side.error_p_reg_9_LC_2_19_1 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_9_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_9_LC_2_19_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_side.error_p_reg_9_LC_2_19_1  (
            .in0(N__27894),
            .in1(N__50222),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\pid_side.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51429),
            .ce(),
            .sr(N__50702));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25160),
            .lcout(drone_altitude_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25151),
            .lcout(drone_altitude_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_2_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_2_19_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(N__25796),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20180),
            .lcout(drone_altitude_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20174),
            .lcout(drone_altitude_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_19_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_19_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_19_7  (
            .in0(_gnd_net_),
            .in1(N__20186),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_altitude_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_2_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_2_20_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_10_LC_2_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_10_LC_2_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37130),
            .lcout(\dron_frame_decoder_1.drone_altitude_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_2_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_11_LC_2_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_11_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37052),
            .lcout(\dron_frame_decoder_1.drone_altitude_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_2_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_12_LC_2_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_12_LC_2_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36946),
            .lcout(drone_altitude_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_2_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_15_LC_2_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_15_LC_2_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36632),
            .lcout(drone_altitude_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_2_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_2_20_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_8_LC_2_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_8_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42611),
            .lcout(\dron_frame_decoder_1.drone_altitude_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36808),
            .lcout(\dron_frame_decoder_1.drone_altitude_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51417),
            .ce(N__25823),
            .sr(N__49588));
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_21_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_21_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_4_LC_2_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_4_LC_2_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40396),
            .lcout(alt_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51402),
            .ce(N__25880),
            .sr(N__49597));
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_21_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_5_LC_2_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_5_LC_2_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40250),
            .lcout(alt_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51402),
            .ce(N__25880),
            .sr(N__49597));
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_21_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_21_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_6_LC_2_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_6_LC_2_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40142),
            .lcout(alt_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51402),
            .ce(N__25880),
            .sr(N__49597));
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_21_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_21_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_esr_7_LC_2_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_esr_7_LC_2_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40011),
            .lcout(alt_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51402),
            .ce(N__25880),
            .sr(N__49597));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_23_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_23_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_23_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_23_1  (
            .in0(N__50806),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39527),
            .lcout(alt_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51376),
            .ce(N__25952),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_5  (
            .in0(N__50807),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39380),
            .lcout(alt_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51376),
            .ce(N__25952),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_2_23_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_2_23_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_2_23_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_2_23_6  (
            .in0(_gnd_net_),
            .in1(N__40272),
            .in2(_gnd_net_),
            .in3(N__50805),
            .lcout(alt_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51376),
            .ce(N__25952),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_23_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_23_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_23_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_23_7  (
            .in0(N__50808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40141),
            .lcout(alt_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51376),
            .ce(N__25952),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_3_5_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_3_5_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_3_LC_3_5_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_3_LC_3_5_0  (
            .in0(N__50821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39334),
            .lcout(alt_kd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51539),
            .ce(N__21928),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_5_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_5_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_0_LC_3_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_0_LC_3_5_1  (
            .in0(_gnd_net_),
            .in1(N__39769),
            .in2(_gnd_net_),
            .in3(N__50820),
            .lcout(alt_kd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51539),
            .ce(N__21928),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_3_5_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_3_5_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kd_4_LC_3_5_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kd_4_LC_3_5_7  (
            .in0(_gnd_net_),
            .in1(N__40379),
            .in2(_gnd_net_),
            .in3(N__50822),
            .lcout(alt_kd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51539),
            .ce(N__21928),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_3_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_2_0_LC_3_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_2_0_LC_3_8_4  (
            .in0(N__39742),
            .in1(N__23651),
            .in2(N__39497),
            .in3(N__21419),
            .lcout(\Commands_frame_decoder.N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_2_LC_3_10_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_reg_esr_2_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_reg_esr_2_LC_3_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_reg_esr_2_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20339),
            .lcout(\pid_alt.error_i_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51519),
            .ce(N__20322),
            .sr(N__50709));
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_3_11_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_6_LC_3_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_6_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40122),
            .lcout(frame_decoder_OFF4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51513),
            .ce(N__26963),
            .sr(N__49515));
    defparam \pid_alt.error_i_acumm_10_LC_3_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_10_LC_3_12_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_10_LC_3_12_0 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \pid_alt.error_i_acumm_10_LC_3_12_0  (
            .in0(N__20441),
            .in1(N__20488),
            .in2(N__31948),
            .in3(N__22648),
            .lcout(\pid_alt.error_i_acummZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51506),
            .ce(),
            .sr(N__33225));
    defparam \pid_alt.error_i_acumm_6_LC_3_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_6_LC_3_12_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_6_LC_3_12_2 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \pid_alt.error_i_acumm_6_LC_3_12_2  (
            .in0(N__20456),
            .in1(N__20647),
            .in2(N__31949),
            .in3(N__22649),
            .lcout(\pid_alt.error_i_acummZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51506),
            .ce(),
            .sr(N__33225));
    defparam \pid_alt.error_i_acumm_8_LC_3_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_8_LC_3_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_8_LC_3_12_4 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \pid_alt.error_i_acumm_8_LC_3_12_4  (
            .in0(N__20393),
            .in1(N__20575),
            .in2(N__31950),
            .in3(N__22650),
            .lcout(\pid_alt.error_i_acummZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51506),
            .ce(),
            .sr(N__33225));
    defparam \pid_alt.error_i_acumm_9_LC_3_12_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_9_LC_3_12_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_9_LC_3_12_5 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \pid_alt.error_i_acumm_9_LC_3_12_5  (
            .in0(N__22651),
            .in1(N__31910),
            .in2(N__20417),
            .in3(N__20539),
            .lcout(\pid_alt.error_i_acummZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51506),
            .ce(),
            .sr(N__33225));
    defparam \pid_alt.pid_prereg_esr_RNIL6HQ_3_LC_3_12_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIL6HQ_3_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIL6HQ_3_LC_3_12_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIL6HQ_3_LC_3_12_6  (
            .in0(_gnd_net_),
            .in1(N__31466),
            .in2(_gnd_net_),
            .in3(N__31892),
            .lcout(\pid_alt.N_306_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI08CV_10_LC_3_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI08CV_10_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI08CV_10_LC_3_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI08CV_10_LC_3_13_0  (
            .in0(N__20455),
            .in1(N__23736),
            .in2(N__20440),
            .in3(N__24030),
            .lcout(\pid_alt.m39_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20611),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51496),
            .ce(N__25561),
            .sr(N__49523));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGERC1_10_LC_3_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGERC1_10_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIGERC1_10_LC_3_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIGERC1_10_LC_3_13_2  (
            .in0(N__20454),
            .in1(N__22314),
            .in2(N__20439),
            .in3(N__22596),
            .lcout(\pid_alt.un1_reset_1_i_a5_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20696),
            .lcout(\pid_alt.error_i_acumm7lto4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51496),
            .ce(N__25561),
            .sr(N__49523));
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20666),
            .lcout(\pid_alt.error_i_acumm7lto5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51496),
            .ce(N__25561),
            .sr(N__49523));
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_10_LC_3_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_10_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51496),
            .ce(N__25561),
            .sr(N__49523));
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24544),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51496),
            .ce(N__25561),
            .sr(N__49523));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6ECV_11_LC_3_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6ECV_11_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI6ECV_11_LC_3_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI6ECV_11_LC_3_13_7  (
            .in0(N__20409),
            .in1(N__20388),
            .in2(N__23740),
            .in3(N__24104),
            .lcout(\pid_alt.un1_reset_1_i_a5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0  (
            .in0(_gnd_net_),
            .in1(N__24988),
            .in2(N__25015),
            .in3(_gnd_net_),
            .lcout(\pid_alt.un1_pid_prereg_0 ),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__22361),
            .in2(N__20372),
            .in3(N__20360),
            .lcout(\pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_0 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2  (
            .in0(_gnd_net_),
            .in1(N__22355),
            .in2(N__20357),
            .in3(N__20342),
            .lcout(\pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_1 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__22349),
            .in2(N__20732),
            .in3(N__20717),
            .lcout(\pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_2 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(N__22583),
            .in2(N__20714),
            .in3(N__20681),
            .lcout(\pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_3 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNI67I91_5_LC_3_14_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNI67I91_5_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNI67I91_5_LC_3_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNI67I91_5_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__20678),
            .in2(N__22373),
            .in3(N__20651),
            .lcout(\pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_4 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6  (
            .in0(_gnd_net_),
            .in1(N__20648),
            .in2(N__20633),
            .in3(N__20597),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_5 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(N__21977),
            .in2(N__20594),
            .in3(N__20579),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_6 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__20576),
            .in2(N__20561),
            .in3(N__20543),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__20540),
            .in2(N__20525),
            .in3(N__20492),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_8 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__20489),
            .in2(N__20474),
            .in3(N__20459),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_9 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__21994),
            .in2(N__20879),
            .in3(N__20864),
            .lcout(\pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_10 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIG2KM_12_LC_3_15_4 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIG2KM_12_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIG2KM_12_LC_3_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIG2KM_12_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__24080),
            .in2(N__20861),
            .in3(N__20843),
            .lcout(\pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_11 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .C_ON=1'b1;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__33281),
            .in2(N__20840),
            .in3(N__20822),
            .lcout(\pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_12 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__20819),
            .in2(_gnd_net_),
            .in3(N__20804),
            .lcout(\pid_alt.error_i_reg_esr_RNI15KJZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_13 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__20801),
            .in2(_gnd_net_),
            .in3(N__20786),
            .lcout(\pid_alt.error_i_reg_esr_RNI38LJZ0Z_15 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_14 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__20783),
            .in2(_gnd_net_),
            .in3(N__20768),
            .lcout(\pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__20765),
            .in2(_gnd_net_),
            .in3(N__20750),
            .lcout(\pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_16 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__20747),
            .in2(_gnd_net_),
            .in3(N__20735),
            .lcout(\pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_17 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .C_ON=1'b1;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(N__21053),
            .in2(_gnd_net_),
            .in3(N__21038),
            .lcout(\pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_18 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .C_ON=1'b1;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__21031),
            .in2(_gnd_net_),
            .in3(N__21035),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ ),
            .ltout(),
            .carryin(\pid_alt.un1_error_i_acumm_prereg_cry_19 ),
            .carryout(\pid_alt.un1_error_i_acumm_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .C_ON=1'b0;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5  (
            .in0(N__21032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21014),
            .lcout(\pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_16_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_16_6  (
            .in0(N__21011),
            .in1(N__22753),
            .in2(N__21005),
            .in3(N__20985),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_7  (
            .in0(N__22175),
            .in1(N__22190),
            .in2(N__22982),
            .in3(N__24120),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_17_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_17_0  (
            .in0(N__20897),
            .in1(N__25659),
            .in2(N__22916),
            .in3(N__20887),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_17_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_17_1 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_17_1  (
            .in0(N__20969),
            .in1(N__20948),
            .in2(_gnd_net_),
            .in3(N__20930),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_17_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_17_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__25660),
            .in2(N__20891),
            .in3(N__20888),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_17_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_17_3 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_17_3  (
            .in0(N__21085),
            .in1(N__21094),
            .in2(_gnd_net_),
            .in3(N__21117),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_17_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_16_LC_3_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_16_LC_3_17_4  (
            .in0(N__21119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51444),
            .ce(N__25570),
            .sr(N__49551));
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_17_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_17_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_17_5  (
            .in0(N__21068),
            .in1(N__25597),
            .in2(_gnd_net_),
            .in3(N__28538),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_17_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_17_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_17_6  (
            .in0(N__21118),
            .in1(_gnd_net_),
            .in2(N__21098),
            .in3(N__21086),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_17_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_17_7  (
            .in0(N__22945),
            .in1(N__25596),
            .in2(N__21062),
            .in3(N__28537),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_18_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto3_LC_3_18_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto3_LC_3_18_0  (
            .in0(N__39498),
            .in1(N__39364),
            .in2(_gnd_net_),
            .in3(N__39633),
            .lcout(),
            .ltout(\Commands_frame_decoder.source_CH1data8lt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_18_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_LC_3_18_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_LC_3_18_1  (
            .in0(N__40138),
            .in1(N__40400),
            .in2(N__21059),
            .in3(N__21412),
            .lcout(\Commands_frame_decoder.source_CH1data8 ),
            .ltout(\Commands_frame_decoder.source_CH1data8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_18_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_1_LC_3_18_2 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \Commands_frame_decoder.source_CH1data_1_LC_3_18_2  (
            .in0(N__25497),
            .in1(N__21184),
            .in2(N__21056),
            .in3(N__39634),
            .lcout(alt_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51430),
            .ce(),
            .sr(N__49561));
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_18_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_18_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_2_LC_3_18_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_2_LC_3_18_3  (
            .in0(N__21430),
            .in1(N__39499),
            .in2(N__21902),
            .in3(N__25498),
            .lcout(alt_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51430),
            .ce(),
            .sr(N__49561));
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_18_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_3_LC_3_18_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_3_LC_3_18_4  (
            .in0(N__25499),
            .in1(N__39365),
            .in2(N__21833),
            .in3(N__21431),
            .lcout(alt_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51430),
            .ce(),
            .sr(N__49561));
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_18_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH1data_0_LC_3_18_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Commands_frame_decoder.source_CH1data_0_LC_3_18_5  (
            .in0(N__21429),
            .in1(N__39770),
            .in2(N__21257),
            .in3(N__25496),
            .lcout(alt_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51430),
            .ce(),
            .sr(N__49561));
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_3_18_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_CH1data8lto7_1_LC_3_18_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.source_CH1data8lto7_1_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__39994),
            .in2(_gnd_net_),
            .in3(N__40257),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_LC_3_19_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_LC_3_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.error_cry_0_c_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\pid_alt.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_3_19_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_RNI1N2F_LC_3_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_0_c_RNI1N2F_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__23144),
            .in2(_gnd_net_),
            .in3(N__21353),
            .lcout(\pid_alt.error_1 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_0 ),
            .carryout(\pid_alt.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_3_19_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_1_c_RNI3Q3F_LC_3_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_1_c_RNI3Q3F_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__23033),
            .in2(_gnd_net_),
            .in3(N__21311),
            .lcout(\pid_alt.error_2 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_1 ),
            .carryout(\pid_alt.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_3_19_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_2_c_RNI5T4F_LC_3_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_2_c_RNI5T4F_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__23027),
            .in2(_gnd_net_),
            .in3(N__21260),
            .lcout(\pid_alt.error_3 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_2 ),
            .carryout(\pid_alt.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_3_19_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_3_c_RNIKE1T_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_3_c_RNIKE1T_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__25034),
            .in2(N__21256),
            .in3(N__21194),
            .lcout(\pid_alt.error_4 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_3 ),
            .carryout(\pid_alt.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_3_19_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_4_c_RNINI2T_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_4_c_RNINI2T_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__21191),
            .in2(N__21185),
            .in3(N__21128),
            .lcout(\pid_alt.error_5 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_4 ),
            .carryout(\pid_alt.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_3_19_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_5_c_RNIQM3T_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_5_c_RNIQM3T_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__21125),
            .in2(N__21901),
            .in3(N__21842),
            .lcout(\pid_alt.error_6 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_5 ),
            .carryout(\pid_alt.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_3_19_7 .C_ON=1'b1;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_6_c_RNITQ4T_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_6_c_RNITQ4T_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__21839),
            .in2(N__21832),
            .in3(N__21785),
            .lcout(\pid_alt.error_7 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_6 ),
            .carryout(\pid_alt.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_3_20_0 .C_ON=1'b1;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_7_c_RNI9LEM_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_7_c_RNI9LEM_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__21782),
            .in2(N__21776),
            .in3(N__21719),
            .lcout(\pid_alt.error_8 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\pid_alt.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_3_20_1 .C_ON=1'b1;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_8_c_RNICPFM_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_8_c_RNICPFM_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__21716),
            .in2(N__21710),
            .in3(N__21653),
            .lcout(\pid_alt.error_9 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_8 ),
            .carryout(\pid_alt.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_3_20_2 .C_ON=1'b1;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_9_c_RNIMMUJ_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_9_c_RNIMMUJ_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__21650),
            .in2(N__21644),
            .in3(N__21587),
            .lcout(\pid_alt.error_10 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_9 ),
            .carryout(\pid_alt.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_3_20_3 .C_ON=1'b1;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_10_c_RNI0SDO_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_cry_10_c_RNI0SDO_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__22001),
            .in2(N__21584),
            .in3(N__21530),
            .lcout(\pid_alt.error_11 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_10 ),
            .carryout(\pid_alt.error_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_3_20_4 .C_ON=1'b1;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_11_c_RNI5JAH_LC_3_20_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_cry_11_c_RNI5JAH_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23129),
            .in3(N__21482),
            .lcout(\pid_alt.error_12 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_11 ),
            .carryout(\pid_alt.error_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_3_20_5 .C_ON=1'b1;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_12_c_RNI7MBH_LC_3_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_12_c_RNI7MBH_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__23057),
            .in2(_gnd_net_),
            .in3(N__21434),
            .lcout(\pid_alt.error_13 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_12 ),
            .carryout(\pid_alt.error_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_3_20_6 .C_ON=1'b1;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_13_c_RNI9PCH_LC_3_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_cry_13_c_RNI9PCH_LC_3_20_6  (
            .in0(_gnd_net_),
            .in1(N__23045),
            .in2(_gnd_net_),
            .in3(N__22049),
            .lcout(\pid_alt.error_14 ),
            .ltout(),
            .carryin(\pid_alt.error_cry_13 ),
            .carryout(\pid_alt.error_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_3_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_14_c_RNIBSDH_LC_3_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \pid_alt.error_cry_14_c_RNIBSDH_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(N__22046),
            .in2(_gnd_net_),
            .in3(N__22040),
            .lcout(\pid_alt.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_21_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22007),
            .lcout(drone_altitude_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_11_LC_3_22_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_11_LC_3_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_11_LC_3_22_1 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_alt.error_i_acumm_11_LC_3_22_1  (
            .in0(N__23747),
            .in1(N__31988),
            .in2(N__21995),
            .in3(N__22660),
            .lcout(\pid_alt.error_i_acummZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51377),
            .ce(),
            .sr(N__33227));
    defparam \pid_alt.error_i_acumm_7_LC_3_22_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_7_LC_3_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_7_LC_3_22_2 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \pid_alt.error_i_acumm_7_LC_3_22_2  (
            .in0(N__31987),
            .in1(N__21970),
            .in2(N__22664),
            .in3(N__24043),
            .lcout(\pid_alt.error_i_acummZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51377),
            .ce(),
            .sr(N__33227));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_23_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_23_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_23_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__39652),
            .in2(_gnd_net_),
            .in3(N__50803),
            .lcout(alt_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51362),
            .ce(N__25948),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_23_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_23_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_23_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_23_7  (
            .in0(N__50804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40010),
            .lcout(alt_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51362),
            .ce(N__25948),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_6_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIRSI31_11_LC_4_6_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIRSI31_11_LC_4_6_7  (
            .in0(N__23534),
            .in1(N__27612),
            .in2(_gnd_net_),
            .in3(N__49772),
            .lcout(\Commands_frame_decoder.state_RNIRSI31Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_4_7_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_1_LC_4_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_1_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__39761),
            .in2(_gnd_net_),
            .in3(N__40001),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_4_7_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_1_LC_4_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_1_LC_4_7_1  (
            .in0(N__23545),
            .in1(N__39483),
            .in2(N__22136),
            .in3(N__40261),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_1_LC_4_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_1_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_1_LC_4_8_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_1_LC_4_8_1  (
            .in0(N__23655),
            .in1(N__26901),
            .in2(N__22133),
            .in3(N__27440),
            .lcout(\Commands_frame_decoder.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51524),
            .ce(),
            .sr(N__49504));
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_4_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNI6QPK_14_LC_4_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Commands_frame_decoder.state_RNI6QPK_14_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__27265),
            .in2(_gnd_net_),
            .in3(N__23650),
            .lcout(\Commands_frame_decoder.N_382_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_4_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_4_10_1 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH4data_ess_7_LC_4_10_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Commands_frame_decoder.source_CH4data_ess_7_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__39983),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51514),
            .ce(N__25318),
            .sr(N__49509));
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_5_LC_4_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_5_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40246),
            .lcout(frame_decoder_CH4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51514),
            .ce(N__25318),
            .sr(N__49509));
    defparam \pid_alt.state_1_LC_4_11_6 .C_ON=1'b0;
    defparam \pid_alt.state_1_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_1_LC_4_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.state_1_LC_4_11_6  (
            .in0(N__31167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51507),
            .ce(),
            .sr(N__49512));
    defparam \Commands_frame_decoder.state_5_LC_4_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_5_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_5_LC_4_11_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_5_LC_4_11_7  (
            .in0(N__23612),
            .in1(N__25451),
            .in2(_gnd_net_),
            .in3(N__26903),
            .lcout(\Commands_frame_decoder.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51507),
            .ce(),
            .sr(N__49512));
    defparam \pid_alt.error_d_reg_prev_esr_RNIFBF74_12_LC_4_12_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFBF74_12_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIFBF74_12_LC_4_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIFBF74_12_LC_4_12_0  (
            .in0(N__22228),
            .in1(N__22124),
            .in2(N__22708),
            .in3(N__22114),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_12_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_12_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_12_1  (
            .in0(N__22219),
            .in1(N__23989),
            .in2(_gnd_net_),
            .in3(N__23592),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_12_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_12_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_12_2  (
            .in0(N__22229),
            .in1(_gnd_net_),
            .in2(N__22118),
            .in3(N__22115),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_12_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_12_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_12_3  (
            .in0(N__22300),
            .in1(N__22277),
            .in2(_gnd_net_),
            .in3(N__22257),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJ0N32_11_LC_4_12_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJ0N32_11_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJ0N32_11_LC_4_12_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJ0N32_11_LC_4_12_5  (
            .in0(N__22199),
            .in1(N__23774),
            .in2(_gnd_net_),
            .in3(N__24220),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_12_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_12_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_12_6  (
            .in0(N__23593),
            .in1(_gnd_net_),
            .in2(N__23993),
            .in3(N__22220),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIKFGA4_11_LC_4_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKFGA4_11_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIKFGA4_11_LC_4_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIKFGA4_11_LC_4_12_7  (
            .in0(N__23845),
            .in1(N__23773),
            .in2(N__22193),
            .in3(N__24219),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_13_1 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_13_1  (
            .in0(N__22426),
            .in1(_gnd_net_),
            .in2(N__22406),
            .in3(N__22157),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_13_2 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__22171),
            .in2(N__22178),
            .in3(N__24127),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_13_3 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_13_3  (
            .in0(N__28624),
            .in1(_gnd_net_),
            .in2(N__28612),
            .in3(N__28572),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_13_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_13_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_13_4  (
            .in0(N__22156),
            .in1(N__22402),
            .in2(_gnd_net_),
            .in3(N__22425),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_13_5  (
            .in0(N__22393),
            .in1(N__23020),
            .in2(N__22430),
            .in3(N__24150),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_14_LC_4_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_14_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22427),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51486),
            .ce(N__25558),
            .sr(N__49519));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_13_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_13_7  (
            .in0(N__22394),
            .in1(N__22379),
            .in2(_gnd_net_),
            .in3(N__24151),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_5_LC_4_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_5_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_5_LC_4_14_0 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \pid_alt.error_i_acumm_esr_5_LC_4_14_0  (
            .in0(N__22316),
            .in1(N__22330),
            .in2(N__22343),
            .in3(N__22628),
            .lcout(\pid_alt.error_i_acummZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_4_14_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_4_14_1 .LUT_INIT=16'b0000110100000101;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_4_14_1  (
            .in0(N__33336),
            .in1(N__33314),
            .in2(N__33393),
            .in3(N__24099),
            .lcout(\pid_alt.N_295 ),
            .ltout(\pid_alt.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_1_LC_4_14_2 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_1_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__22676),
            .in2(N__22364),
            .in3(N__24056),
            .lcout(\pid_alt.error_i_acummZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_2_LC_4_14_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_2_LC_4_14_3  (
            .in0(N__22630),
            .in1(_gnd_net_),
            .in2(N__22682),
            .in3(N__24011),
            .lcout(\pid_alt.error_i_acummZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_3_LC_4_14_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_alt.error_i_acumm_esr_3_LC_4_14_4  (
            .in0(N__24071),
            .in1(N__22631),
            .in2(_gnd_net_),
            .in3(N__22680),
            .lcout(\pid_alt.error_i_acummZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIP4VR2_4_LC_4_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIP4VR2_4_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIP4VR2_4_LC_4_14_5 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIP4VR2_4_LC_4_14_5  (
            .in0(N__22603),
            .in1(N__22339),
            .in2(N__22331),
            .in3(N__22315),
            .lcout(\pid_alt.N_294 ),
            .ltout(\pid_alt.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_0_LC_4_14_6 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_0_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__22629),
            .in2(N__22685),
            .in3(N__24977),
            .lcout(\pid_alt.error_i_acummZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_4_LC_4_14_7 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \pid_alt.error_i_acumm_esr_4_LC_4_14_7  (
            .in0(N__22681),
            .in1(_gnd_net_),
            .in2(N__22647),
            .in3(N__22604),
            .lcout(\pid_alt.error_i_acummZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51474),
            .ce(N__33256),
            .sr(N__33197));
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_15_0 .C_ON=1'b1;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__23185),
            .in2(N__23189),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_0_LC_4_15_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_0_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_0_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__22567),
            .in2(N__22556),
            .in3(N__22541),
            .lcout(\pid_alt.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_1_LC_4_15_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_1_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_1_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__22538),
            .in2(N__24199),
            .in3(N__22526),
            .lcout(\pid_alt.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_0 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_2_LC_4_15_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_2_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_2_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__22523),
            .in2(N__24177),
            .in3(N__22511),
            .lcout(\pid_alt.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_1 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_3_LC_4_15_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_3_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_3_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__22508),
            .in2(N__24246),
            .in3(N__22496),
            .lcout(\pid_alt.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_2 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_4_LC_4_15_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_4_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_4_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__22489),
            .in2(N__22472),
            .in3(N__22460),
            .lcout(\pid_alt.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_3 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_5_LC_4_15_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_5_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_5_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__22457),
            .in2(N__22448),
            .in3(N__22829),
            .lcout(\pid_alt.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_4 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_6_LC_4_15_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_6_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_6_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__22826),
            .in2(N__22813),
            .in3(N__22784),
            .lcout(\pid_alt.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_5 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_6 ),
            .clk(N__51462),
            .ce(N__25562),
            .sr(N__49531));
    defparam \pid_alt.pid_prereg_esr_7_LC_4_16_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_7_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_7_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__24530),
            .in2(N__24575),
            .in3(N__22781),
            .lcout(\pid_alt.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_8_LC_4_16_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_8_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_8_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__24395),
            .in2(N__24670),
            .in3(N__22778),
            .lcout(\pid_alt.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_7 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_9_LC_4_16_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_9_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_9_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__22775),
            .in2(N__24358),
            .in3(N__22766),
            .lcout(\pid_alt.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_8 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_10_LC_4_16_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_10_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_10_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__22763),
            .in2(N__22757),
            .in3(N__22739),
            .lcout(\pid_alt.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_9 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_11_LC_4_16_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_11_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_11_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__23954),
            .in2(N__23977),
            .in3(N__22736),
            .lcout(\pid_alt.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_10 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_12_LC_4_16_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_12_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_12_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__22733),
            .in2(N__23852),
            .in3(N__22724),
            .lcout(\pid_alt.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_11 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_13_LC_4_16_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_13_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_13_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__22721),
            .in2(N__22712),
            .in3(N__22688),
            .lcout(\pid_alt.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_12 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_14_LC_4_16_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_14_LC_4_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_14_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(N__23021),
            .in2(N__23006),
            .in3(N__22994),
            .lcout(\pid_alt.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_13 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_14 ),
            .clk(N__51445),
            .ce(N__25566),
            .sr(N__49539));
    defparam \pid_alt.pid_prereg_esr_15_LC_4_17_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_15_LC_4_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_15_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__22991),
            .in2(N__22981),
            .in3(N__22955),
            .lcout(\pid_alt.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_16_LC_4_17_1 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_16_LC_4_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_16_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__22952),
            .in2(N__22946),
            .in3(N__22925),
            .lcout(\pid_alt.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_15 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_17_LC_4_17_2 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_17_LC_4_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_17_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__22922),
            .in2(N__22915),
            .in3(N__22898),
            .lcout(\pid_alt.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_16 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_18_LC_4_17_3 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_18_LC_4_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_18_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__22895),
            .in2(N__22886),
            .in3(N__22871),
            .lcout(\pid_alt.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_17 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_19_LC_4_17_4 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_19_LC_4_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_19_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__22868),
            .in2(N__22859),
            .in3(N__22838),
            .lcout(\pid_alt.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_18 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_20_LC_4_17_5 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_20_LC_4_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_20_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__24926),
            .in2(N__24949),
            .in3(N__22835),
            .lcout(\pid_alt.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_19 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_21_LC_4_17_6 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_21_LC_4_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_21_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(N__24695),
            .in2(N__24815),
            .in3(N__22832),
            .lcout(\pid_alt.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_20 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_22_LC_4_17_7 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_17_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_22_LC_4_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_22_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(N__23120),
            .in2(N__23105),
            .in3(N__23108),
            .lcout(\pid_alt.pid_preregZ0Z_22 ),
            .ltout(),
            .carryin(\pid_alt.un1_pid_prereg_0_cry_21 ),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_22 ),
            .clk(N__51431),
            .ce(N__25567),
            .sr(N__49546));
    defparam \pid_alt.pid_prereg_esr_23_LC_4_18_0 .C_ON=1'b1;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_23_LC_4_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.pid_prereg_esr_23_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__23104),
            .in2(N__23078),
            .in3(N__23063),
            .lcout(\pid_alt.pid_preregZ0Z_23 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\pid_alt.un1_pid_prereg_0_cry_23 ),
            .clk(N__51418),
            .ce(N__25571),
            .sr(N__49552));
    defparam \pid_alt.pid_prereg_esr_24_LC_4_18_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.pid_prereg_esr_24_LC_4_18_1 .LUT_INIT=16'b1000000101111110;
    LogicCell40 \pid_alt.pid_prereg_esr_24_LC_4_18_1  (
            .in0(N__24754),
            .in1(N__24727),
            .in2(N__24800),
            .in3(N__23060),
            .lcout(\pid_alt.pid_preregZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51418),
            .ce(N__25571),
            .sr(N__49552));
    defparam \pid_alt.error_axb_13_LC_4_19_0 .C_ON=1'b0;
    defparam \pid_alt.error_axb_13_LC_4_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_13_LC_4_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_13_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23051),
            .lcout(\pid_alt.error_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_4_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_4_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_13_LC_4_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_13_LC_4_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36879),
            .lcout(drone_altitude_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51403),
            .ce(N__25819),
            .sr(N__49562));
    defparam \pid_alt.error_axb_14_LC_4_19_2 .C_ON=1'b0;
    defparam \pid_alt.error_axb_14_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_14_LC_4_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_14_LC_4_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23039),
            .lcout(\pid_alt.error_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48435),
            .lcout(drone_altitude_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51403),
            .ce(N__25819),
            .sr(N__49562));
    defparam \pid_alt.error_axb_2_LC_4_19_4 .C_ON=1'b0;
    defparam \pid_alt.error_axb_2_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_2_LC_4_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_2_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24683),
            .lcout(\pid_alt.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_3_LC_4_19_5 .C_ON=1'b0;
    defparam \pid_alt.error_axb_3_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_3_LC_4_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_3_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24677),
            .lcout(\pid_alt.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_4_19_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_4_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_4_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23681),
            .lcout(\pid_alt.error_d_reg_prev_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_4_20_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_4_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23162),
            .lcout(drone_H_disp_side_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_4_20_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_4_20_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_4_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_4_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42606),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51388),
            .ce(N__29587),
            .sr(N__49569));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_4_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_4_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23156),
            .lcout(drone_H_disp_side_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_4_20_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_4_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_4_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36807),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51388),
            .ce(N__29587),
            .sr(N__49569));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_4_20_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_4_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23150),
            .lcout(drone_H_disp_side_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_4_20_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_4_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_4_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37128),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51388),
            .ce(N__29587),
            .sr(N__49569));
    defparam \pid_alt.error_axb_1_LC_4_20_6 .C_ON=1'b0;
    defparam \pid_alt.error_axb_1_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_1_LC_4_20_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pid_alt.error_axb_1_LC_4_20_6  (
            .in0(_gnd_net_),
            .in1(N__24689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_axb_12_LC_4_20_7 .C_ON=1'b0;
    defparam \pid_alt.error_axb_12_LC_4_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_axb_12_LC_4_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_axb_12_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(\pid_alt.error_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_inv_LC_4_21_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_inv_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_inv_LC_4_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_cry_0_c_inv_LC_4_21_0  (
            .in0(_gnd_net_),
            .in1(N__23321),
            .in2(_gnd_net_),
            .in3(N__27154),
            .lcout(\pid_side.error_axb_0 ),
            .ltout(),
            .carryin(bfn_4_21_0_),
            .carryout(\pid_side.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_4_21_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_4_21_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_c_RNI43F5_LC_4_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_0_c_RNI43F5_LC_4_21_1  (
            .in0(_gnd_net_),
            .in1(N__28466),
            .in2(_gnd_net_),
            .in3(N__23300),
            .lcout(\pid_side.error_1 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0 ),
            .carryout(\pid_side.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_4_21_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_c_RNI66G5_LC_4_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_1_c_RNI66G5_LC_4_21_2  (
            .in0(_gnd_net_),
            .in1(N__25991),
            .in2(_gnd_net_),
            .in3(N__23285),
            .lcout(\pid_side.error_2 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1 ),
            .carryout(\pid_side.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_4_21_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_c_RNI89H5_LC_4_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_2_c_RNI89H5_LC_4_21_3  (
            .in0(_gnd_net_),
            .in1(N__25982),
            .in2(_gnd_net_),
            .in3(N__23267),
            .lcout(\pid_side.error_3 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2 ),
            .carryout(\pid_side.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_4_21_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_c_RNI1SDJ_LC_4_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_c_RNI1SDJ_LC_4_21_4  (
            .in0(_gnd_net_),
            .in1(N__25223),
            .in2(N__25766),
            .in3(N__23252),
            .lcout(\pid_side.error_4 ),
            .ltout(),
            .carryin(\pid_side.error_cry_3 ),
            .carryout(\pid_side.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_4_21_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_4_21_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_0_0_c_RNIF3ET_LC_4_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_0_0_c_RNIF3ET_LC_4_21_5  (
            .in0(_gnd_net_),
            .in1(N__25214),
            .in2(N__25742),
            .in3(N__23237),
            .lcout(\pid_side.error_5 ),
            .ltout(),
            .carryin(\pid_side.error_cry_0_0 ),
            .carryout(\pid_side.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_4_21_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_4_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_1_0_c_RNII9K11_LC_4_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_1_0_c_RNII9K11_LC_4_21_6  (
            .in0(_gnd_net_),
            .in1(N__25229),
            .in2(N__25208),
            .in3(N__23219),
            .lcout(\pid_side.error_6 ),
            .ltout(),
            .carryin(\pid_side.error_cry_1_0 ),
            .carryout(\pid_side.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_4_21_7 .C_ON=1'b1;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_2_0_c_RNILFQL_LC_4_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_2_0_c_RNILFQL_LC_4_21_7  (
            .in0(_gnd_net_),
            .in1(N__25199),
            .in2(N__25754),
            .in3(N__23201),
            .lcout(\pid_side.error_7 ),
            .ltout(),
            .carryin(\pid_side.error_cry_2_0 ),
            .carryout(\pid_side.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_4_22_0 .C_ON=1'b1;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_4_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_3_0_c_RNIOL0Q_LC_4_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_3_0_c_RNIOL0Q_LC_4_22_0  (
            .in0(_gnd_net_),
            .in1(N__23198),
            .in2(N__25193),
            .in3(N__23480),
            .lcout(\pid_side.error_8 ),
            .ltout(),
            .carryin(bfn_4_22_0_),
            .carryout(\pid_side.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_4_22_1 .C_ON=1'b1;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_4_c_RNIC8FJ_LC_4_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_4_c_RNIC8FJ_LC_4_22_1  (
            .in0(_gnd_net_),
            .in1(N__23477),
            .in2(N__25184),
            .in3(N__23453),
            .lcout(\pid_side.error_9 ),
            .ltout(),
            .carryin(\pid_side.error_cry_4 ),
            .carryout(\pid_side.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_4_22_2 .C_ON=1'b1;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_4_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_5_c_RNIM4IS_LC_4_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_5_c_RNIM4IS_LC_4_22_2  (
            .in0(_gnd_net_),
            .in1(N__25175),
            .in2(N__23450),
            .in3(N__23423),
            .lcout(\pid_side.error_10 ),
            .ltout(),
            .carryin(\pid_side.error_cry_5 ),
            .carryout(\pid_side.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_4_22_3 .C_ON=1'b1;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_6_c_RNIQBMT_LC_4_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_side.error_cry_6_c_RNIQBMT_LC_4_22_3  (
            .in0(_gnd_net_),
            .in1(N__28493),
            .in2(_gnd_net_),
            .in3(N__23405),
            .lcout(\pid_side.error_11 ),
            .ltout(),
            .carryin(\pid_side.error_cry_6 ),
            .carryout(\pid_side.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_4_22_4 .C_ON=1'b1;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_4_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_7_c_RNIPRDP1_LC_4_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_7_c_RNIPRDP1_LC_4_22_4  (
            .in0(_gnd_net_),
            .in1(N__28520),
            .in2(N__29549),
            .in3(N__23387),
            .lcout(\pid_side.error_12 ),
            .ltout(),
            .carryin(\pid_side.error_cry_7 ),
            .carryout(\pid_side.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_4_22_5 .C_ON=1'b1;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_4_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_8_c_RNIUUKS_LC_4_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_8_c_RNIUUKS_LC_4_22_5  (
            .in0(_gnd_net_),
            .in1(N__29636),
            .in2(N__29522),
            .in3(N__23369),
            .lcout(\pid_side.error_13 ),
            .ltout(),
            .carryin(\pid_side.error_cry_8 ),
            .carryout(\pid_side.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_4_22_6 .C_ON=1'b1;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_9_c_RNI13MS_LC_4_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_side.error_cry_9_c_RNI13MS_LC_4_22_6  (
            .in0(_gnd_net_),
            .in1(N__24956),
            .in2(N__29612),
            .in3(N__23351),
            .lcout(\pid_side.error_14 ),
            .ltout(),
            .carryin(\pid_side.error_cry_9 ),
            .carryout(\pid_side.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_4_22_7 .C_ON=1'b0;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_4_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_cry_10_c_RNIBCT11_LC_4_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_side.error_cry_10_c_RNIBCT11_LC_4_22_7  (
            .in0(N__25169),
            .in1(N__29611),
            .in2(_gnd_net_),
            .in3(N__23348),
            .lcout(\pid_side.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_4_23_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_4_23_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_kp_e_0_0_LC_4_23_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_e_0_0_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__39768),
            .in2(_gnd_net_),
            .in3(N__50802),
            .lcout(alt_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51352),
            .ce(N__25947),
            .sr(_gnd_net_));
    defparam \pid_alt.state_0_LC_5_6_7 .C_ON=1'b0;
    defparam \pid_alt.state_0_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.state_0_LC_5_6_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_alt.state_0_LC_5_6_7  (
            .in0(N__31147),
            .in1(N__32842),
            .in2(_gnd_net_),
            .in3(N__32022),
            .lcout(\pid_alt.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51529),
            .ce(),
            .sr(N__49498));
    defparam \Commands_frame_decoder.state_12_LC_5_7_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_12_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_12_LC_5_7_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_12_LC_5_7_3  (
            .in0(N__23533),
            .in1(N__27609),
            .in2(N__25306),
            .in3(N__26913),
            .lcout(\Commands_frame_decoder.stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51525),
            .ce(),
            .sr(N__49500));
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_0_LC_5_8_4 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_0_LC_5_8_4  (
            .in0(N__23560),
            .in1(N__27438),
            .in2(N__23669),
            .in3(N__23570),
            .lcout(),
            .ltout(\Commands_frame_decoder.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_8_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_0_LC_5_8_5 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_0_LC_5_8_5  (
            .in0(N__23546),
            .in1(N__23561),
            .in2(N__23552),
            .in3(N__25352),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_0_LC_5_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_0_LC_5_8_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.state_0_LC_5_8_6 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Commands_frame_decoder.state_0_LC_5_8_6  (
            .in0(N__26880),
            .in1(N__23656),
            .in2(N__23549),
            .in3(N__25340),
            .lcout(\Commands_frame_decoder.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51520),
            .ce(),
            .sr(N__49502));
    defparam \Commands_frame_decoder.state_2_LC_5_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_2_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_2_LC_5_8_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_2_LC_5_8_7  (
            .in0(N__27439),
            .in1(N__23621),
            .in2(N__25429),
            .in3(N__26879),
            .lcout(\Commands_frame_decoder.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51520),
            .ce(),
            .sr(N__49502));
    defparam \Commands_frame_decoder.preinit_LC_5_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_LC_5_9_2 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.preinit_LC_5_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.preinit_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__25251),
            .in2(_gnd_net_),
            .in3(N__27607),
            .lcout(\Commands_frame_decoder.preinitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51515),
            .ce(),
            .sr(N__49505));
    defparam \Commands_frame_decoder.state_11_LC_5_9_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_11_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_11_LC_5_9_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_11_LC_5_9_7  (
            .in0(N__27606),
            .in1(N__23529),
            .in2(N__26825),
            .in3(N__26902),
            .lcout(\Commands_frame_decoder.stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51515),
            .ce(),
            .sr(N__49505));
    defparam \scaler_4.N_1684_i_l_ofx_LC_5_10_2 .C_ON=1'b0;
    defparam \scaler_4.N_1684_i_l_ofx_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.N_1684_i_l_ofx_LC_5_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.N_1684_i_l_ofx_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__25394),
            .in2(_gnd_net_),
            .in3(N__23510),
            .lcout(\scaler_4.N_1684_i_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_3_0_LC_5_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_3_0_LC_5_10_3  (
            .in0(N__39697),
            .in1(N__39974),
            .in2(N__39467),
            .in3(N__40238),
            .lcout(\Commands_frame_decoder.state_ns_i_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_1_2_LC_5_10_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Commands_frame_decoder.state_RNO_1_2_LC_5_10_4  (
            .in0(N__39975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39698),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNO_0_2_LC_5_10_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Commands_frame_decoder.state_RNO_0_2_LC_5_10_5  (
            .in0(N__39439),
            .in1(N__23657),
            .in2(N__23624),
            .in3(N__40239),
            .lcout(\Commands_frame_decoder.state_ns_0_a3_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_2_LC_5_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_2_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_2_LC_5_10_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \uart_pc.data_2_LC_5_10_6  (
            .in0(N__28769),
            .in1(N__27421),
            .in2(N__39474),
            .in3(N__28874),
            .lcout(uart_pc_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51508),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_5_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIHL1J_5_LC_5_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIHL1J_5_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__23611),
            .in2(_gnd_net_),
            .in3(N__27568),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_5_11_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIE28S_5_LC_5_11_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Commands_frame_decoder.state_RNIE28S_5_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23600),
            .in3(N__49750),
            .lcout(\Commands_frame_decoder.source_CH4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_0_LC_5_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_0_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_0_LC_5_11_5 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_0_LC_5_11_5  (
            .in0(N__28775),
            .in1(N__27420),
            .in2(N__27344),
            .in3(N__39706),
            .lcout(uart_pc_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51497),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_5_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIQRI31_10_LC_5_11_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIQRI31_10_LC_5_11_6  (
            .in0(N__27567),
            .in1(N__26818),
            .in2(_gnd_net_),
            .in3(N__49749),
            .lcout(\Commands_frame_decoder.state_RNIQRI31Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_12_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_15_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_15_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28576),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51487),
            .ce(N__25554),
            .sr(N__49513));
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_12_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_12_LC_5_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_12_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23597),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51487),
            .ce(N__25554),
            .sr(N__49513));
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_5_13_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_5_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_5_13_0  (
            .in0(N__23830),
            .in1(N__23861),
            .in2(N__23981),
            .in3(N__23763),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_13_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_13_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_13_1  (
            .in0(N__23942),
            .in1(N__23915),
            .in2(_gnd_net_),
            .in3(N__23891),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_5_13_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_5_13_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_5_13_2  (
            .in0(N__23831),
            .in1(_gnd_net_),
            .in2(N__23855),
            .in3(N__23764),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_5_13_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_5_13_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_5_13_3  (
            .in0(N__23788),
            .in1(N__23797),
            .in2(_gnd_net_),
            .in3(N__23820),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_13_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_11_LC_5_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_11_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23822),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51475),
            .ce(N__25555),
            .sr(N__49516));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_5_13_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_5_13_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_5_13_6  (
            .in0(N__23821),
            .in1(_gnd_net_),
            .in2(N__23801),
            .in3(N__23789),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_5_13_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_11_LC_5_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_11_LC_5_13_7  (
            .in0(N__23765),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51475),
            .ce(N__25555),
            .sr(N__49516));
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_5_14_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_0_LC_5_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_0_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23717),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_5_14_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_3_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_3_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24247),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_5_14_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_12_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_12_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24224),
            .lcout(\pid_alt.error_i_acumm7lto12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_5_14_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_1_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_1_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24200),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_5_14_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_2_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_2_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24178),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_5_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_14_LC_5_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_14_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24155),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_5_14_7 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_15_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_15_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24131),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51463),
            .ce(N__25559),
            .sr(N__49520));
    defparam \pid_alt.error_i_acumm_esr_12_LC_5_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_12_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_12_LC_5_15_0 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \pid_alt.error_i_acumm_esr_12_LC_5_15_0  (
            .in0(N__33319),
            .in1(N__33395),
            .in2(N__33346),
            .in3(N__24100),
            .lcout(\pid_alt.error_i_acummZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51446),
            .ce(N__33255),
            .sr(N__33196));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRFAQ1_0_LC_5_15_1 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRFAQ1_0_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRFAQ1_0_LC_5_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRFAQ1_0_LC_5_15_1  (
            .in0(N__24067),
            .in1(N__24055),
            .in2(N__24044),
            .in3(N__24973),
            .lcout(),
            .ltout(\pid_alt.un1_reset_1_i_a5_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE78O2_2_LC_5_15_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE78O2_2_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIE78O2_2_LC_5_15_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIE78O2_2_LC_5_15_2  (
            .in0(N__33318),
            .in1(N__24007),
            .in2(N__23996),
            .in3(N__31968),
            .lcout(\pid_alt.un1_reset_1_i_a5_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_5_15_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_5_15_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_5_15_3  (
            .in0(N__24446),
            .in1(N__25730),
            .in2(N__25616),
            .in3(N__24440),
            .lcout(\pid_alt.N_557 ),
            .ltout(\pid_alt.N_557_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIVV9C5_10_LC_5_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIVV9C5_10_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIVV9C5_10_LC_5_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIVV9C5_10_LC_5_15_4  (
            .in0(N__24434),
            .in1(N__24422),
            .in2(N__24410),
            .in3(N__24407),
            .lcout(),
            .ltout(\pid_alt.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HS46_21_LC_5_15_5 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HS46_21_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNI8HS46_21_LC_5_15_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNI8HS46_21_LC_5_15_5  (
            .in0(N__31969),
            .in1(N__33394),
            .in2(N__24401),
            .in3(N__49042),
            .lcout(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21 ),
            .ltout(\pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIT64J6_1_LC_5_15_6 .C_ON=1'b0;
    defparam \pid_alt.state_RNIT64J6_1_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIT64J6_1_LC_5_15_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_alt.state_RNIT64J6_1_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24398),
            .in3(N__31970),
            .lcout(\pid_alt.N_72_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_0  (
            .in0(N__24262),
            .in1(N__24389),
            .in2(N__24671),
            .in3(N__24379),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_1 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_1  (
            .in0(N__24616),
            .in1(N__24625),
            .in2(_gnd_net_),
            .in3(N__24651),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2  (
            .in0(N__24263),
            .in1(_gnd_net_),
            .in2(N__24383),
            .in3(N__24380),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_3 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_3  (
            .in0(N__24341),
            .in1(N__24317),
            .in2(_gnd_net_),
            .in3(N__24296),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_7_LC_5_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_7_LC_5_16_4  (
            .in0(N__24653),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51432),
            .ce(N__25563),
            .sr(N__49532));
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_16_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_16_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_16_5  (
            .in0(N__24590),
            .in1(_gnd_net_),
            .in2(N__24599),
            .in3(N__24551),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_6 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_6  (
            .in0(N__24652),
            .in1(_gnd_net_),
            .in2(N__24629),
            .in3(N__24617),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_16_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_16_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_16_7  (
            .in0(N__24589),
            .in1(N__24574),
            .in2(N__24554),
            .in3(N__24550),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_17_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_17_6  (
            .in0(N__24524),
            .in1(N__24518),
            .in2(N__24512),
            .in3(N__24503),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_17_7 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_17_7  (
            .in0(N__24497),
            .in1(N__24491),
            .in2(N__24485),
            .in3(N__24476),
            .lcout(\pid_alt.source_pid_1_sqmuxa_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_5_18_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_5_18_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_5_18_0  (
            .in0(N__24862),
            .in1(N__24871),
            .in2(_gnd_net_),
            .in3(N__24843),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_5_18_1 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_5_18_1 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_5_18_1  (
            .in0(N__24919),
            .in1(N__24470),
            .in2(_gnd_net_),
            .in3(N__24886),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_5_18_2 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_5_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_5_18_2  (
            .in0(N__24950),
            .in1(N__24785),
            .in2(N__24929),
            .in3(N__25635),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_5_18_3 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_5_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_19_LC_5_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_19_LC_5_18_3  (
            .in0(N__24920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51404),
            .ce(N__25568),
            .sr(N__49547));
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_5_18_4 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_5_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_d_reg_prev_esr_20_LC_5_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_20_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24844),
            .lcout(\pid_alt.error_d_reg_prevZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51404),
            .ce(N__25568),
            .sr(N__49547));
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_5_18_5 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_5_18_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_5_18_5  (
            .in0(N__24872),
            .in1(N__24863),
            .in2(_gnd_net_),
            .in3(N__24845),
            .lcout(\pid_alt.un1_pid_prereg_236_1 ),
            .ltout(\pid_alt.un1_pid_prereg_236_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_5_18_6 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_5_18_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_5_18_6  (
            .in0(_gnd_net_),
            .in1(N__24824),
            .in2(N__24818),
            .in3(N__25636),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19 ),
            .ltout(\pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_5_18_7 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_5_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_5_18_7  (
            .in0(N__24786),
            .in1(N__24750),
            .in2(N__24734),
            .in3(N__24726),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_19_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36796),
            .lcout(drone_altitude_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_5_19_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_5_19_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_2_LC_5_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_2_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37118),
            .lcout(drone_altitude_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_5_19_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_5_19_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_3_LC_5_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_3_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37044),
            .lcout(drone_altitude_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_19_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36969),
            .lcout(\dron_frame_decoder_1.drone_altitude_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36878),
            .lcout(\dron_frame_decoder_1.drone_altitude_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_19_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48434),
            .lcout(\dron_frame_decoder_1.drone_altitude_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51389),
            .ce(N__33470),
            .sr(N__49553));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_5_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_5_20_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_0_LC_5_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_0_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(N__39755),
            .in2(_gnd_net_),
            .in3(N__50809),
            .lcout(xy_kp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51378),
            .ce(N__39026),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_5_20_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_2_LC_5_20_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_2_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(N__39525),
            .in2(_gnd_net_),
            .in3(N__50810),
            .lcout(xy_kp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51378),
            .ce(N__39026),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_5_20_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_5_20_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_5_LC_5_20_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_5_LC_5_20_5  (
            .in0(N__50811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40093),
            .lcout(xy_kp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51378),
            .ce(N__39026),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_20_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25040),
            .lcout(drone_altitude_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_5_21_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_0_LC_5_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_0_LC_5_21_0  (
            .in0(_gnd_net_),
            .in1(N__25022),
            .in2(_gnd_net_),
            .in3(N__24998),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51363),
            .ce(N__25574),
            .sr(N__49570));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_5_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_5_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_5_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29632),
            .lcout(drone_H_disp_side_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_5_21_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_5_21_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_5_21_6  (
            .in0(_gnd_net_),
            .in1(N__27113),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_5_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_5_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_0_LC_5_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_0_LC_5_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39759),
            .lcout(side_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_5_22_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_5_22_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_1_LC_5_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_1_LC_5_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39653),
            .lcout(side_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_5_22_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_5_22_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_2_LC_5_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_2_LC_5_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39526),
            .lcout(side_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_5_22_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_5_22_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_3_LC_5_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_3_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39366),
            .lcout(side_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_5_22_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_5_22_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_4_LC_5_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_4_LC_5_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40402),
            .lcout(side_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_5_22_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_5_22_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_5_LC_5_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_5_LC_5_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40274),
            .lcout(side_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_5_22_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_5_22_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH2data_esr_6_LC_5_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_esr_6_LC_5_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40121),
            .lcout(side_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51353),
            .ce(N__27047),
            .sr(N__49580));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_5_23_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_5_23_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_5_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_5_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36627),
            .lcout(drone_H_disp_side_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51343),
            .ce(N__29591),
            .sr(N__49589));
    defparam \Commands_frame_decoder.source_data_valid_LC_7_6_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_data_valid_LC_7_6_4 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \Commands_frame_decoder.source_data_valid_LC_7_6_4  (
            .in0(N__26090),
            .in1(N__25262),
            .in2(N__27186),
            .in3(N__27614),
            .lcout(debug_CH3_20A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51521),
            .ce(),
            .sr(N__49499));
    defparam \Commands_frame_decoder.state_13_LC_7_7_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_13_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_13_LC_7_7_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_13_LC_7_7_3  (
            .in0(N__27597),
            .in1(N__25286),
            .in2(N__25307),
            .in3(N__26851),
            .lcout(\Commands_frame_decoder.stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51516),
            .ce(),
            .sr(N__49501));
    defparam \Commands_frame_decoder.state_14_LC_7_7_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_14_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_14_LC_7_7_4 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_14_LC_7_7_4  (
            .in0(N__25285),
            .in1(N__27598),
            .in2(_gnd_net_),
            .in3(N__25336),
            .lcout(\Commands_frame_decoder.stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51516),
            .ce(),
            .sr(N__49501));
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_8_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_8_0 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_8_0  (
            .in0(N__26178),
            .in1(N__26196),
            .in2(N__26162),
            .in3(N__26212),
            .lcout(\Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_7_8_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNII19A1_4_LC_7_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Commands_frame_decoder.WDT_RNII19A1_4_LC_7_8_1  (
            .in0(N__26245),
            .in1(N__26020),
            .in2(N__26231),
            .in3(N__26035),
            .lcout(\Commands_frame_decoder.WDT_RNII19A1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_7_8_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNID7P31_6_LC_7_8_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Commands_frame_decoder.WDT_RNID7P31_6_LC_7_8_2  (
            .in0(N__26179),
            .in1(N__26005),
            .in2(_gnd_net_),
            .in3(N__26197),
            .lcout(),
            .ltout(\Commands_frame_decoder.WDT8lto13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_7_8_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_7_8_3 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_7_8_3  (
            .in0(N__26260),
            .in1(N__25277),
            .in2(N__25271),
            .in3(N__25268),
            .lcout(\Commands_frame_decoder.WDT8lt14_0 ),
            .ltout(\Commands_frame_decoder.WDT8lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_7_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.preinit_RNIF92K5_LC_7_8_4 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \Commands_frame_decoder.preinit_RNIF92K5_LC_7_8_4  (
            .in0(N__26141),
            .in1(N__25261),
            .in2(N__25232),
            .in3(N__26115),
            .lcout(\Commands_frame_decoder.state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_7_8_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_7_8_5 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_7_8_5  (
            .in0(N__25361),
            .in1(N__26143),
            .in2(N__27608),
            .in3(N__26116),
            .lcout(\Commands_frame_decoder.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_7_8_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_7_8_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_7_8_6  (
            .in0(N__26142),
            .in1(N__27577),
            .in2(N__26120),
            .in3(N__25360),
            .lcout(\Commands_frame_decoder.N_377_0 ),
            .ltout(\Commands_frame_decoder.N_377_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_8_7 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_8_7  (
            .in0(N__27254),
            .in1(N__27230),
            .in2(N__25343),
            .in3(N__27578),
            .lcout(\Commands_frame_decoder.N_384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_9_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_0_LC_7_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_0_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39754),
            .lcout(frame_decoder_CH4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_9_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_1_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_1_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39577),
            .lcout(frame_decoder_CH4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_9_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_2_LC_7_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_2_LC_7_9_2  (
            .in0(N__39487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(frame_decoder_CH4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_9_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_3_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_3_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39344),
            .lcout(frame_decoder_CH4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_9_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_4_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_4_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40359),
            .lcout(frame_decoder_CH4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_9_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH4data_esr_6_LC_7_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH4data_esr_6_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40106),
            .lcout(frame_decoder_CH4data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51498),
            .ce(N__25325),
            .sr(N__49506));
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_10_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_0_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_0_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39753),
            .lcout(frame_decoder_OFF4data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_10_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_1_LC_7_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_1_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39594),
            .lcout(frame_decoder_OFF4data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_10_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_2_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_2_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39466),
            .lcout(frame_decoder_OFF4data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39343),
            .lcout(frame_decoder_OFF4data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_10_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_4_LC_7_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_4_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40378),
            .lcout(frame_decoder_OFF4data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_offset4data_esr_5_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_esr_5_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40254),
            .lcout(frame_decoder_OFF4data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_10_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_10_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_offset4data_ess_7_LC_7_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_offset4data_ess_7_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39982),
            .lcout(frame_decoder_OFF4data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51488),
            .ce(N__26956),
            .sr(N__49508));
    defparam \Commands_frame_decoder.state_6_LC_7_11_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_6_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_6_LC_7_11_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \Commands_frame_decoder.state_6_LC_7_11_1  (
            .in0(N__25379),
            .in1(N__26702),
            .in2(_gnd_net_),
            .in3(N__26894),
            .lcout(\Commands_frame_decoder.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51476),
            .ce(),
            .sr(N__49510));
    defparam \uart_pc.data_rdy_LC_7_11_5 .C_ON=1'b0;
    defparam \uart_pc.data_rdy_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_rdy_LC_7_11_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.data_rdy_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__40704),
            .in2(_gnd_net_),
            .in3(N__28799),
            .lcout(uart_pc_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51476),
            .ce(),
            .sr(N__49510));
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_11_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIGK1J_4_LC_7_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIGK1J_4_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__25369),
            .in2(_gnd_net_),
            .in3(N__27491),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_4_LC_7_11_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Commands_frame_decoder.state_4_LC_7_11_7  (
            .in0(N__25370),
            .in1(N__25786),
            .in2(_gnd_net_),
            .in3(N__26893),
            .lcout(\Commands_frame_decoder.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51476),
            .ce(),
            .sr(N__49510));
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_7_12_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_7_12_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_7_12_0  (
            .in0(N__26676),
            .in1(N__26493),
            .in2(_gnd_net_),
            .in3(N__26569),
            .lcout(\dron_frame_decoder_1.WDT10lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_7_12_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_7_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_7_12_2  (
            .in0(N__26524),
            .in1(N__26584),
            .in2(N__26603),
            .in3(N__26539),
            .lcout(),
            .ltout(\dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_7_12_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_7_12_3 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_7_12_3  (
            .in0(N__26554),
            .in1(N__25457),
            .in2(N__25469),
            .in3(N__25466),
            .lcout(\dron_frame_decoder_1.WDT10lt14_0 ),
            .ltout(\dron_frame_decoder_1.WDT10lt14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_7_12_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_7_12_4 .LUT_INIT=16'b0000001111111111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__27780),
            .in2(N__25460),
            .in3(N__27801),
            .lcout(\dron_frame_decoder_1.WDT10_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_7_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_7_12_7 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_7_12_7  (
            .in0(N__26494),
            .in1(N__26509),
            .in2(N__26660),
            .in3(N__26677),
            .lcout(\dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNID18S_4_LC_7_13_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNID18S_4_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__25450),
            .in2(_gnd_net_),
            .in3(N__49748),
            .lcout(\Commands_frame_decoder.source_CH3data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_6_LC_7_13_2 .C_ON=1'b0;
    defparam \uart_pc.data_6_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_6_LC_7_13_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_6_LC_7_13_2  (
            .in0(N__28774),
            .in1(N__27422),
            .in2(N__40562),
            .in3(N__39930),
            .lcout(uart_pc_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51447),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__25405),
            .in2(_gnd_net_),
            .in3(N__27536),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_14_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIEI1J_2_LC_7_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNIEI1J_2_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(_gnd_net_),
            .in3(N__27537),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0 ),
            .ltout(\Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_3_LC_7_14_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_3_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_3_LC_7_14_3 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_3_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__25406),
            .in2(N__25409),
            .in3(N__26914),
            .lcout(\Commands_frame_decoder.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51433),
            .ce(),
            .sr(N__49521));
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_7_15_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_7_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_7_15_0  (
            .in0(N__25670),
            .in1(N__25646),
            .in2(N__25700),
            .in3(N__25583),
            .lcout(\pid_alt.m7_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_7_15_4 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_19_LC_7_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_19_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25721),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51419),
            .ce(N__25556),
            .sr(N__49524));
    defparam \pid_alt.pid_prereg_esr_RNI046H1_1_LC_7_15_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI046H1_1_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI046H1_1_LC_7_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI046H1_1_LC_7_15_5  (
            .in0(N__30590),
            .in1(N__31483),
            .in2(N__30648),
            .in3(N__31516),
            .lcout(),
            .ltout(\pid_alt.un1_reset_i_a5_1_10_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIJF5N2_10_LC_7_15_6 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIJF5N2_10_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIJF5N2_10_LC_7_15_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIJF5N2_10_LC_7_15_6  (
            .in0(N__30547),
            .in1(N__30298),
            .in2(N__25691),
            .in3(N__29140),
            .lcout(\pid_alt.un1_reset_i_a5_1_10_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_7_16_0 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_18_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_18_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25688),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51405),
            .ce(N__25560),
            .sr(N__49533));
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_7_16_2 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_17_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_17_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25664),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51405),
            .ce(N__25560),
            .sr(N__49533));
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_7_16_3 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_20_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_20_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25640),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51405),
            .ce(N__25560),
            .sr(N__49533));
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_7_16_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_prereg_esr_16_LC_7_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.error_i_acumm_prereg_esr_16_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25601),
            .lcout(\pid_alt.error_i_acumm_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51405),
            .ce(N__25560),
            .sr(N__49533));
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_17_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIBV7S_2_LC_7_17_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIBV7S_2_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__25486),
            .in2(_gnd_net_),
            .in3(N__49767),
            .lcout(\Commands_frame_decoder.un1_sink_data_valid_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_7_17_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_7_17_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_7_17_5  (
            .in0(N__25865),
            .in1(N__25853),
            .in2(N__25844),
            .in3(N__25832),
            .lcout(\pid_alt.N_551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIFCSD1_0_LC_7_18_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIFCSD1_0_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIFCSD1_0_LC_7_18_4 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \pid_alt.state_RNIFCSD1_0_LC_7_18_4  (
            .in0(N__32841),
            .in1(N__31986),
            .in2(N__31178),
            .in3(N__49747),
            .lcout(\pid_alt.state_RNIFCSD1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_18_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_18_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__26780),
            .in2(_gnd_net_),
            .in3(N__49033),
            .lcout(\dron_frame_decoder_1.N_755_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_7_19_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_7_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_7_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36616),
            .lcout(\dron_frame_decoder_1.drone_altitude_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51364),
            .ce(N__33462),
            .sr(N__49554));
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_20_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIC08S_3_LC_7_20_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.state_RNIC08S_3_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__25787),
            .in2(_gnd_net_),
            .in3(N__49768),
            .lcout(\Commands_frame_decoder.source_CH2data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_7_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI36DT_4_LC_7_21_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI36DT_4_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__28097),
            .in2(_gnd_net_),
            .in3(N__49773),
            .lcout(\dron_frame_decoder_1.N_747_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_7_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_7_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27125),
            .lcout(drone_H_disp_side_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_7_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_7_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27104),
            .lcout(drone_H_disp_side_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_7_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_7_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27119),
            .lcout(drone_H_disp_side_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_2_LC_7_21_6 .C_ON=1'b0;
    defparam \pid_side.error_axb_2_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_2_LC_7_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_2_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27137),
            .lcout(\pid_side.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_3_LC_7_21_7 .C_ON=1'b0;
    defparam \pid_side.error_axb_3_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_3_LC_7_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_side.error_axb_3_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27131),
            .lcout(\pid_side.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_22_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_22_6 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_alt_kp_4_LC_7_22_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_alt_kp_4_LC_7_22_6  (
            .in0(N__25966),
            .in1(N__27611),
            .in2(N__26719),
            .in3(N__40401),
            .lcout(alt_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51336),
            .ce(),
            .sr(N__49581));
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIF38S_6_LC_7_23_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIF38S_6_LC_7_23_5  (
            .in0(N__26712),
            .in1(N__27610),
            .in2(_gnd_net_),
            .in3(N__49771),
            .lcout(\Commands_frame_decoder.state_RNIF38SZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_7 .C_ON=1'b0;
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNICP2N1_0_LC_7_29_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNICP2N1_0_LC_7_29_7  (
            .in0(_gnd_net_),
            .in1(N__25922),
            .in2(_gnd_net_),
            .in3(N__50795),
            .lcout(\pid_alt.N_850_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_1 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_1__0__0_LC_8_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_1__0__0_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25892),
            .lcout(\uart_drone_sync.aux_1__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51536),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_7 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_0__0__0_LC_8_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_0__0__0_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25898),
            .lcout(\uart_drone_sync.aux_0__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51536),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_1 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_2__0__0_LC_8_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_2__0__0_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25886),
            .lcout(\uart_drone_sync.aux_2__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51533),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_6_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.source_data_1_esr_ctle_14_LC_8_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \scaler_4.source_data_1_esr_ctle_14_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__27176),
            .in2(_gnd_net_),
            .in3(N__49752),
            .lcout(\scaler_4.debug_CH3_20A_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_8_6_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.source_data_valid_RNO_0_LC_8_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.source_data_valid_RNO_0_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__27219),
            .in2(_gnd_net_),
            .in3(N__27255),
            .lcout(\Commands_frame_decoder.count_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.WDT_0_LC_8_7_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_0_LC_8_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_0_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__26069),
            .in2(N__26084),
            .in3(N__26083),
            .lcout(\Commands_frame_decoder.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_1_LC_8_7_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_1_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_1_LC_8_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_1_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__26063),
            .in2(_gnd_net_),
            .in3(N__26057),
            .lcout(\Commands_frame_decoder.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_0 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_2_LC_8_7_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_2_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_2_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_2_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__26054),
            .in2(_gnd_net_),
            .in3(N__26048),
            .lcout(\Commands_frame_decoder.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_1 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_3_LC_8_7_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_3_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_3_LC_8_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_3_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__26045),
            .in2(_gnd_net_),
            .in3(N__26039),
            .lcout(\Commands_frame_decoder.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_2 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_4_LC_8_7_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_4_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_4_LC_8_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_4_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__26036),
            .in2(_gnd_net_),
            .in3(N__26024),
            .lcout(\Commands_frame_decoder.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_3 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_5_LC_8_7_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_5_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_5_LC_8_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_5_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__26021),
            .in2(_gnd_net_),
            .in3(N__26009),
            .lcout(\Commands_frame_decoder.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_4 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_6_LC_8_7_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_6_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_6_LC_8_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_6_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__26006),
            .in2(_gnd_net_),
            .in3(N__25994),
            .lcout(\Commands_frame_decoder.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_5 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_7_LC_8_7_7 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_7_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_7_LC_8_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_7_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__26261),
            .in2(_gnd_net_),
            .in3(N__26249),
            .lcout(\Commands_frame_decoder.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_6 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_7 ),
            .clk(N__51509),
            .ce(),
            .sr(N__26462));
    defparam \Commands_frame_decoder.WDT_8_LC_8_8_0 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_8_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_8_LC_8_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_8_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__26246),
            .in2(_gnd_net_),
            .in3(N__26234),
            .lcout(\Commands_frame_decoder.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_9_LC_8_8_1 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_9_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_9_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_9_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__26230),
            .in2(_gnd_net_),
            .in3(N__26216),
            .lcout(\Commands_frame_decoder.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_8 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_10_LC_8_8_2 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_10_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_10_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_10_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__26213),
            .in2(_gnd_net_),
            .in3(N__26201),
            .lcout(\Commands_frame_decoder.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_9 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_11_LC_8_8_3 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_11_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_11_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_11_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__26198),
            .in2(_gnd_net_),
            .in3(N__26183),
            .lcout(\Commands_frame_decoder.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_10 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_12_LC_8_8_4 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_12_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_12_LC_8_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_12_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__26180),
            .in2(_gnd_net_),
            .in3(N__26165),
            .lcout(\Commands_frame_decoder.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_11 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_13_LC_8_8_5 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_13_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_13_LC_8_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_13_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__26161),
            .in2(_gnd_net_),
            .in3(N__26147),
            .lcout(\Commands_frame_decoder.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_12 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_14_LC_8_8_6 .C_ON=1'b1;
    defparam \Commands_frame_decoder.WDT_14_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_14_LC_8_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Commands_frame_decoder.WDT_14_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__26144),
            .in2(_gnd_net_),
            .in3(N__26126),
            .lcout(\Commands_frame_decoder.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\Commands_frame_decoder.un1_WDT_cry_13 ),
            .carryout(\Commands_frame_decoder.un1_WDT_cry_14 ),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \Commands_frame_decoder.WDT_15_LC_8_8_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.WDT_15_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.WDT_15_LC_8_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Commands_frame_decoder.WDT_15_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__26114),
            .in2(_gnd_net_),
            .in3(N__26123),
            .lcout(\Commands_frame_decoder.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51499),
            .ce(),
            .sr(N__26458));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_9_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__28937),
            .in2(N__28974),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_9_1 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__26399),
            .in2(N__26393),
            .in3(N__26384),
            .lcout(\scaler_4.un2_source_data_0 ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_0 ),
            .carryout(\scaler_4.un3_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_9_2 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__26381),
            .in2(N__26375),
            .in3(N__26366),
            .lcout(\scaler_4.un3_source_data_0_cry_1_c_RNI74CL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_1 ),
            .carryout(\scaler_4.un3_source_data_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_9_3 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__26363),
            .in2(N__26357),
            .in3(N__26348),
            .lcout(\scaler_4.un3_source_data_0_cry_2_c_RNIA8DL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_2 ),
            .carryout(\scaler_4.un3_source_data_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_9_4 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__26345),
            .in2(N__26339),
            .in3(N__26330),
            .lcout(\scaler_4.un3_source_data_0_cry_3_c_RNIDCEL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_3 ),
            .carryout(\scaler_4.un3_source_data_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_9_5 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__26327),
            .in2(N__26315),
            .in3(N__26306),
            .lcout(\scaler_4.un3_source_data_0_cry_4_c_RNIGGFL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_4 ),
            .carryout(\scaler_4.un3_source_data_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_9_6 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__26303),
            .in2(N__26297),
            .in3(N__26279),
            .lcout(\scaler_4.un3_source_data_0_cry_5_c_RNIJKGL ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_5 ),
            .carryout(\scaler_4.un3_source_data_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_9_7 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__26276),
            .in2(_gnd_net_),
            .in3(N__26264),
            .lcout(\scaler_4.un3_source_data_0_cry_6_c_RNIOUNN ),
            .ltout(),
            .carryin(\scaler_4.un3_source_data_0_cry_6 ),
            .carryout(\scaler_4.un3_source_data_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_10_0 .C_ON=1'b1;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__26477),
            .in2(N__48128),
            .in3(N__26468),
            .lcout(\scaler_4.un3_source_data_0_cry_7_c_RNIP0PN ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\scaler_4.un3_source_data_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_10_1 .C_ON=1'b0;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26465),
            .lcout(\scaler_4.un3_source_data_0_cry_8_c_RNIS918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_10_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.un1_state57_i_LC_8_10_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Commands_frame_decoder.un1_state57_i_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__27535),
            .in2(_gnd_net_),
            .in3(N__49755),
            .lcout(\Commands_frame_decoder.un1_state57_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_1_LC_8_10_6 .C_ON=1'b0;
    defparam \uart_pc.data_1_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_LC_8_10_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_LC_8_10_6  (
            .in0(N__28756),
            .in1(N__27406),
            .in2(N__28856),
            .in3(N__39576),
            .lcout(uart_pc_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51477),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_10_7 .C_ON=1'b0;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_10_7  (
            .in0(N__29007),
            .in1(N__28968),
            .in2(_gnd_net_),
            .in3(N__28938),
            .lcout(\scaler_4.un2_source_data_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_0_LC_8_11_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_0_LC_8_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_0_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__26423),
            .in2(N__26438),
            .in3(N__26437),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_1_LC_8_11_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_1_LC_8_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__26417),
            .in2(_gnd_net_),
            .in3(N__26411),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_1 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_0 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_2_LC_8_11_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_2_LC_8_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_2_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__26408),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_2 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_1 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_3_LC_8_11_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_3_LC_8_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_3_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__26612),
            .in2(_gnd_net_),
            .in3(N__26606),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_3 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_2 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_4_LC_8_11_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_4_LC_8_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_4_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__26588),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_4 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_3 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_5_LC_8_11_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_5_LC_8_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_5_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__26585),
            .in2(_gnd_net_),
            .in3(N__26573),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_5 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_4 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_6_LC_8_11_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_6_LC_8_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_6_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__26570),
            .in2(_gnd_net_),
            .in3(N__26558),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_6 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_5 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_7_LC_8_11_7 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_7_LC_8_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_7_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__26555),
            .in2(_gnd_net_),
            .in3(N__26543),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_7 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_6 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_7 ),
            .clk(N__51464),
            .ce(),
            .sr(N__26633));
    defparam \dron_frame_decoder_1.WDT_8_LC_8_12_0 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_8_LC_8_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_8_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__26540),
            .in2(_gnd_net_),
            .in3(N__26528),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_9_LC_8_12_1 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_9_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_9_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__26525),
            .in2(_gnd_net_),
            .in3(N__26513),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_9 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_8 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_10_LC_8_12_2 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_10_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_10_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__26510),
            .in2(_gnd_net_),
            .in3(N__26498),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_10 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_9 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_11_LC_8_12_3 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_11_LC_8_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_11_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__26495),
            .in2(_gnd_net_),
            .in3(N__26480),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_11 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_10 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_12_LC_8_12_4 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_12_LC_8_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_12_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__26678),
            .in2(_gnd_net_),
            .in3(N__26663),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_12 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_11 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_13_LC_8_12_5 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_13_LC_8_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_13_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__26659),
            .in2(_gnd_net_),
            .in3(N__26645),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_13 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_12 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_14_LC_8_12_6 .C_ON=1'b1;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_14_LC_8_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \dron_frame_decoder_1.WDT_14_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__27784),
            .in2(_gnd_net_),
            .in3(N__26642),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_14 ),
            .ltout(),
            .carryin(\dron_frame_decoder_1.un1_WDT_cry_13 ),
            .carryout(\dron_frame_decoder_1.un1_WDT_cry_14 ),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \dron_frame_decoder_1.WDT_15_LC_8_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.WDT_15_LC_8_12_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \dron_frame_decoder_1.WDT_15_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__27803),
            .in2(_gnd_net_),
            .in3(N__26639),
            .lcout(\dron_frame_decoder_1.WDTZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51448),
            .ce(),
            .sr(N__26623));
    defparam \uart_pc.data_1_4_LC_8_13_0 .C_ON=1'b0;
    defparam \uart_pc.data_1_4_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_1_4_LC_8_13_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \uart_pc.data_1_4_LC_8_13_0  (
            .in0(N__28773),
            .in1(N__27419),
            .in2(N__29081),
            .in3(N__40194),
            .lcout(uart_pc_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51434),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_8_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_8_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__36919),
            .in2(_gnd_net_),
            .in3(N__37009),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_8_13_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_8_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_8_13_2  (
            .in0(N__48426),
            .in1(N__27749),
            .in2(N__26636),
            .in3(N__36759),
            .lcout(\dron_frame_decoder_1.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_13_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__29210),
            .in2(_gnd_net_),
            .in3(N__49759),
            .lcout(\dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_8_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI0TLI1_4_LC_8_14_0 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \dron_frame_decoder_1.state_RNI0TLI1_4_LC_8_14_0  (
            .in0(N__28052),
            .in1(N__26765),
            .in2(N__49796),
            .in3(N__28120),
            .lcout(\dron_frame_decoder_1.N_763_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_14_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_14_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_14_2  (
            .in0(N__28051),
            .in1(N__26764),
            .in2(N__28078),
            .in3(N__28119),
            .lcout(\dron_frame_decoder_1.state_RNI3T3K1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_rdy_LC_8_14_5 .C_ON=1'b0;
    defparam \uart_drone.data_rdy_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_rdy_LC_8_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.data_rdy_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__31054),
            .in2(_gnd_net_),
            .in3(N__29879),
            .lcout(uart_drone_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51420),
            .ce(),
            .sr(N__49525));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_0_1_LC_8_14_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_0_1_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_0_1_LC_8_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_2_0_1_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__29206),
            .in2(_gnd_net_),
            .in3(N__37112),
            .lcout(),
            .ltout(\dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_1_LC_8_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_0_i_a2_2_1_LC_8_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \dron_frame_decoder_1.state_ns_0_i_a2_2_1_LC_8_14_7  (
            .in0(N__36609),
            .in1(N__36848),
            .in2(N__26768),
            .in3(N__42570),
            .lcout(\dron_frame_decoder_1.N_435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_8_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI7Q6K_5_LC_8_15_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \dron_frame_decoder_1.state_RNI7Q6K_5_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__27998),
            .in2(_gnd_net_),
            .in3(N__29195),
            .lcout(\dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_15_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_2_0_LC_8_15_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \dron_frame_decoder_1.state_RNO_2_0_LC_8_15_5  (
            .in0(N__28050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27752),
            .lcout(\dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_8_15_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNITC181_2_LC_8_15_7 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \dron_frame_decoder_1.state_RNITC181_2_LC_8_15_7  (
            .in0(N__29239),
            .in1(N__29196),
            .in2(N__27839),
            .in3(N__49751),
            .lcout(\dron_frame_decoder_1.N_723_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_8_16_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_8_16_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_xy_kp_4_LC_8_16_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_4_LC_8_16_0  (
            .in0(N__26745),
            .in1(N__27603),
            .in2(N__26998),
            .in3(N__40369),
            .lcout(xy_kp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51390),
            .ce(),
            .sr(N__49540));
    defparam \Commands_frame_decoder.state_7_LC_8_16_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_7_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_7_LC_8_16_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_7_LC_8_16_1  (
            .in0(N__27601),
            .in1(N__26991),
            .in2(N__26720),
            .in3(N__26916),
            .lcout(\Commands_frame_decoder.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51390),
            .ce(),
            .sr(N__49540));
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_16_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNIG48S_7_LC_8_16_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \Commands_frame_decoder.state_RNIG48S_7_LC_8_16_2  (
            .in0(N__26990),
            .in1(N__27600),
            .in2(_gnd_net_),
            .in3(N__49756),
            .lcout(\Commands_frame_decoder.state_RNIG48SZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_8_LC_8_16_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_8_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_8_LC_8_16_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \Commands_frame_decoder.state_8_LC_8_16_3  (
            .in0(N__27602),
            .in1(N__26974),
            .in2(N__26999),
            .in3(N__26917),
            .lcout(\Commands_frame_decoder.stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51390),
            .ce(),
            .sr(N__49540));
    defparam \Commands_frame_decoder.state_9_LC_8_16_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_9_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_9_LC_8_16_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Commands_frame_decoder.state_9_LC_8_16_4  (
            .in0(N__26918),
            .in1(N__26936),
            .in2(N__26975),
            .in3(N__27604),
            .lcout(\Commands_frame_decoder.stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51390),
            .ce(),
            .sr(N__49540));
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_16_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNII68S_9_LC_8_16_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Commands_frame_decoder.state_RNII68S_9_LC_8_16_5  (
            .in0(N__49757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26927),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_16_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_RNILP1J_9_LC_8_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_RNILP1J_9_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__26935),
            .in2(_gnd_net_),
            .in3(N__27599),
            .lcout(\Commands_frame_decoder.source_offset4data_1_sqmuxa ),
            .ltout(\Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_10_LC_8_16_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_10_LC_8_16_7 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.state_10_LC_8_16_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \Commands_frame_decoder.state_10_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__26811),
            .in2(N__26921),
            .in3(N__26915),
            .lcout(\Commands_frame_decoder.stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51390),
            .ce(),
            .sr(N__49540));
    defparam \pid_side.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_8_17_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_side.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__49868),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_8_17_1 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_8_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__34708),
            .in2(_gnd_net_),
            .in3(N__26789),
            .lcout(\pid_side.un1_pid_prereg_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_1 ),
            .carryout(\pid_side.un1_pid_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_8_17_2 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_8_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__50107),
            .in2(_gnd_net_),
            .in3(N__26786),
            .lcout(\pid_side.un1_pid_prereg_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_2 ),
            .carryout(\pid_side.un1_pid_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_8_17_3 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_8_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__28381),
            .in2(_gnd_net_),
            .in3(N__26783),
            .lcout(\pid_side.un1_pid_prereg_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_3 ),
            .carryout(\pid_side.un1_pid_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_8_17_4 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_8_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__30865),
            .in2(N__48129),
            .in3(N__27026),
            .lcout(\pid_side.un1_pid_prereg_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_4 ),
            .carryout(\pid_side.un1_pid_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_8_17_5 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_8_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__28348),
            .in2(N__48131),
            .in3(N__27023),
            .lcout(\pid_side.un1_pid_prereg_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_5 ),
            .carryout(\pid_side.un1_pid_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_8_17_6 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_8_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__30361),
            .in2(N__48130),
            .in3(N__27020),
            .lcout(\pid_side.un1_pid_prereg_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_6 ),
            .carryout(\pid_side.un1_pid_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_8_17_7 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_8_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__28450),
            .in2(N__48132),
            .in3(N__27017),
            .lcout(\pid_side.un1_pid_prereg_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_7 ),
            .carryout(\pid_side.un1_pid_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_8_18_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_8_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__48136),
            .in2(N__27907),
            .in3(N__27014),
            .lcout(\pid_side.un1_pid_prereg_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_8_18_1 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_8_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__29405),
            .in2(N__48191),
            .in3(N__27011),
            .lcout(\pid_side.un1_pid_prereg_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_9 ),
            .carryout(\pid_side.un1_pid_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_8_18_2 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_8_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__28420),
            .in2(_gnd_net_),
            .in3(N__27008),
            .lcout(\pid_side.un1_pid_prereg_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_10 ),
            .carryout(\pid_side.un1_pid_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_8_18_3 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_8_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__28709),
            .in2(N__48190),
            .in3(N__27005),
            .lcout(\pid_side.un1_pid_prereg_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_11 ),
            .carryout(\pid_side.un1_pid_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_8_18_4 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_8_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__30832),
            .in2(_gnd_net_),
            .in3(N__27002),
            .lcout(\pid_side.un1_pid_prereg_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_12 ),
            .carryout(\pid_side.un1_pid_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_8_18_5 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_8_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__28234),
            .in2(_gnd_net_),
            .in3(N__27071),
            .lcout(\pid_side.un1_pid_prereg_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_13 ),
            .carryout(\pid_side.un1_pid_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_8_18_6 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_8_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__28267),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\pid_side.un1_pid_prereg_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_14 ),
            .carryout(\pid_side.un1_pid_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_8_18_7 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_8_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__30922),
            .in2(_gnd_net_),
            .in3(N__27065),
            .lcout(\pid_side.un1_pid_prereg_cry_15_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_15 ),
            .carryout(\pid_side.un1_pid_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_8_19_0 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_8_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__28189),
            .in2(_gnd_net_),
            .in3(N__27062),
            .lcout(\pid_side.un1_pid_prereg_cry_16_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\pid_side.un1_pid_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_8_19_1 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_8_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__28657),
            .in2(_gnd_net_),
            .in3(N__27059),
            .lcout(\pid_side.un1_pid_prereg_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_17 ),
            .carryout(\pid_side.un1_pid_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_8_19_2 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_8_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__28306),
            .in2(_gnd_net_),
            .in3(N__27056),
            .lcout(\pid_side.un1_pid_prereg_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_18 ),
            .carryout(\pid_side.un1_pid_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_8_19_3 .C_ON=1'b1;
    defparam \pid_side.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_8_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__28146),
            .in2(_gnd_net_),
            .in3(N__27053),
            .lcout(\pid_side.un1_pid_prereg_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\pid_side.un1_pid_prereg_cry_19 ),
            .carryout(\pid_side.un1_pid_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_21_LC_8_19_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_21_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_21_LC_8_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_side.pid_prereg_esr_21_LC_8_19_4  (
            .in0(N__28147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27050),
            .lcout(\pid_side.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51354),
            .ce(N__41891),
            .sr(N__49563));
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_20_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_20_0 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH2data_ess_7_LC_8_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH2data_ess_7_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40006),
            .lcout(side_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51344),
            .ce(N__27037),
            .sr(N__49571));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_8_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_8_21_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_8_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42605),
            .lcout(drone_H_disp_side_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_8_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_8_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_8_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36803),
            .lcout(drone_H_disp_side_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_8_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_8_21_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_8_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37114),
            .lcout(drone_H_disp_side_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_8_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_8_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_8_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37034),
            .lcout(drone_H_disp_side_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_8_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_8_21_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_8_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36959),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_8_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_8_21_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_8_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36877),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_8_21_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_8_21_6 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_8_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48436),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_8_21_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_8_21_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_8_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36628),
            .lcout(\dron_frame_decoder_1.drone_H_disp_side_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51337),
            .ce(N__27098),
            .sr(N__49582));
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_8_22_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_8_22_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_7_LC_8_22_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_7_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__40005),
            .in2(_gnd_net_),
            .in3(N__50801),
            .lcout(alt_ki_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51329),
            .ce(N__38848),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_0 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_1__0__0_LC_9_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_1__0__0_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27290),
            .lcout(\uart_pc_sync.aux_1__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51534),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_5 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_0__0__0_LC_9_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_0__0__0_LC_9_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27296),
            .lcout(\uart_pc_sync.aux_0__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51534),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_2__0__0_LC_9_2_7 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_2__0__0_LC_9_2_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_pc_sync.aux_2__0__0_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(N__27284),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_pc_sync.aux_2__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51530),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.aux_3__0__0_LC_9_3_1 .C_ON=1'b0;
    defparam \uart_pc_sync.aux_3__0__0_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.aux_3__0__0_LC_9_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.aux_3__0__0_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27278),
            .lcout(\uart_pc_sync.aux_3__0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51526),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc_sync.Q_0__0_LC_9_3_6 .C_ON=1'b0;
    defparam \uart_pc_sync.Q_0__0_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc_sync.Q_0__0_LC_9_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_pc_sync.Q_0__0_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27272),
            .lcout(debug_CH2_18A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51526),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.count_0_LC_9_6_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.count_0_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.count_0_LC_9_6_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \Commands_frame_decoder.count_0_LC_9_6_0  (
            .in0(N__27613),
            .in1(N__27266),
            .in2(N__27229),
            .in3(N__49795),
            .lcout(\Commands_frame_decoder.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51510),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_4_LC_9_7_6 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_4_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_4_LC_9_7_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \scaler_4.source_data_1_4_LC_9_7_6  (
            .in0(N__27193),
            .in1(N__28982),
            .in2(N__36730),
            .in3(N__28949),
            .lcout(scaler_4_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51500),
            .ce(),
            .sr(N__49507));
    defparam \uart_pc.data_5_LC_9_8_0 .C_ON=1'b0;
    defparam \uart_pc.data_5_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_5_LC_9_8_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uart_pc.data_5_LC_9_8_0  (
            .in0(N__27390),
            .in1(N__28730),
            .in2(N__39821),
            .in3(N__40041),
            .lcout(uart_pc_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51489),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_3_LC_9_8_1 .C_ON=1'b0;
    defparam \uart_pc.data_3_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_3_LC_9_8_1 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \uart_pc.data_3_LC_9_8_1  (
            .in0(N__39284),
            .in1(N__28829),
            .in2(N__28741),
            .in3(N__27389),
            .lcout(uart_pc_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51489),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_8_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__40299),
            .in2(_gnd_net_),
            .in3(N__39581),
            .lcout(),
            .ltout(\Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_8_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_8_4  (
            .in0(N__27605),
            .in1(N__40040),
            .in2(N__27443),
            .in3(N__39283),
            .lcout(\Commands_frame_decoder.N_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_9_8_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNILR1B2_2_LC_9_8_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_pc.timer_Count_RNILR1B2_2_LC_9_8_6  (
            .in0(N__40643),
            .in1(N__28791),
            .in2(_gnd_net_),
            .in3(N__48993),
            .lcout(\uart_pc.timer_Count_RNILR1B2Z0Z_2 ),
            .ltout(\uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_4_LC_9_8_7 .C_ON=1'b0;
    defparam \uart_pc.data_4_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_4_LC_9_8_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \uart_pc.data_4_LC_9_8_7  (
            .in0(N__28792),
            .in1(N__27358),
            .in2(N__27362),
            .in3(N__40300),
            .lcout(uart_pc_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51489),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_4_LC_9_9_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_4_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_4_LC_9_9_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_4_LC_9_9_0  (
            .in0(N__29057),
            .in1(N__40650),
            .in2(N__27359),
            .in3(N__40758),
            .lcout(\uart_pc.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51478),
            .ce(),
            .sr(N__40524));
    defparam \uart_pc.data_Aux_0_LC_9_9_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_0_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_0_LC_9_9_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_pc.data_Aux_0_LC_9_9_4  (
            .in0(N__30068),
            .in1(N__27334),
            .in2(N__40676),
            .in3(N__40757),
            .lcout(\uart_pc.data_AuxZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51478),
            .ce(),
            .sr(N__40524));
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_10_0 .C_ON=1'b1;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \scaler_4.un2_source_data_0_cry_1_c_LC_9_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \scaler_4.un2_source_data_0_cry_1_c_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__29000),
            .in2(N__27323),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_6_LC_9_10_1 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_6_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_6_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_6_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__27307),
            .in2(N__29008),
            .in3(N__27314),
            .lcout(scaler_4_data_6),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_1 ),
            .carryout(\scaler_4.un2_source_data_0_cry_2 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_7_LC_9_10_2 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_7_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_7_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_7_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__27715),
            .in2(N__27311),
            .in3(N__27299),
            .lcout(scaler_4_data_7),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_2 ),
            .carryout(\scaler_4.un2_source_data_0_cry_3 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_8_LC_9_10_3 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_8_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_8_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_8_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__27700),
            .in2(N__27719),
            .in3(N__27707),
            .lcout(scaler_4_data_8),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_3 ),
            .carryout(\scaler_4.un2_source_data_0_cry_4 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_9_LC_9_10_4 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_9_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_9_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_9_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__27685),
            .in2(N__27704),
            .in3(N__27692),
            .lcout(scaler_4_data_9),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_4 ),
            .carryout(\scaler_4.un2_source_data_0_cry_5 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_10_LC_9_10_5 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_10_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_10_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_10_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__27670),
            .in2(N__27689),
            .in3(N__27677),
            .lcout(scaler_4_data_10),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_5 ),
            .carryout(\scaler_4.un2_source_data_0_cry_6 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_11_LC_9_10_6 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_11_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_11_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_11_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__27655),
            .in2(N__27674),
            .in3(N__27662),
            .lcout(scaler_4_data_11),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_6 ),
            .carryout(\scaler_4.un2_source_data_0_cry_7 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_12_LC_9_10_7 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_12_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_12_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_12_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__27643),
            .in2(N__27659),
            .in3(N__27647),
            .lcout(scaler_4_data_12),
            .ltout(),
            .carryin(\scaler_4.un2_source_data_0_cry_7 ),
            .carryout(\scaler_4.un2_source_data_0_cry_8 ),
            .clk(N__51465),
            .ce(N__28916),
            .sr(N__49514));
    defparam \scaler_4.source_data_1_esr_13_LC_9_11_0 .C_ON=1'b1;
    defparam \scaler_4.source_data_1_esr_13_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_13_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \scaler_4.source_data_1_esr_13_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__27644),
            .in2(N__27632),
            .in3(N__27623),
            .lcout(scaler_4_data_13),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\scaler_4.un2_source_data_0_cry_9 ),
            .clk(N__51449),
            .ce(N__28911),
            .sr(N__49517));
    defparam \scaler_4.source_data_1_esr_14_LC_9_11_1 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_14_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_14_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \scaler_4.source_data_1_esr_14_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27620),
            .lcout(scaler_4_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51449),
            .ce(N__28911),
            .sr(N__49517));
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_12_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIES9Q1_2_LC_9_12_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uart_drone.timer_Count_RNIES9Q1_2_LC_9_12_3  (
            .in0(N__31042),
            .in1(N__29874),
            .in2(_gnd_net_),
            .in3(N__49022),
            .lcout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2 ),
            .ltout(\uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_12_4 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIRC5U2_2_LC_9_12_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_drone.timer_Count_RNIRC5U2_2_LC_9_12_4  (
            .in0(N__29875),
            .in1(_gnd_net_),
            .in2(N__27617),
            .in3(_gnd_net_),
            .lcout(\uart_drone.data_rdyc_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_ns_i_i_0_a2_2_4_0_LC_9_12_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_ns_i_i_0_a2_2_4_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_ns_i_i_0_a2_2_4_0_LC_9_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \dron_frame_decoder_1.state_ns_i_i_0_a2_2_4_0_LC_9_12_5  (
            .in0(N__36749),
            .in1(N__36908),
            .in2(N__48408),
            .in3(N__36996),
            .lcout(\dron_frame_decoder_1.N_412_4 ),
            .ltout(\dron_frame_decoder_1.N_412_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_12_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_3_LC_9_12_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_3_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27806),
            .in3(N__27942),
            .lcout(\dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_12_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_12_7 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_12_7  (
            .in0(N__27802),
            .in1(N__29220),
            .in2(N__27785),
            .in3(N__27764),
            .lcout(\dron_frame_decoder_1.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_0  (
            .in0(N__28053),
            .in1(N__27750),
            .in2(N__27947),
            .in3(N__29211),
            .lcout(),
            .ltout(\dron_frame_decoder_1.N_177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_0_LC_9_13_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_0_LC_9_13_1 .SEQ_MODE=4'b1001;
    defparam \dron_frame_decoder_1.state_0_LC_9_13_1 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \dron_frame_decoder_1.state_0_LC_9_13_1  (
            .in0(N__28007),
            .in1(N__27751),
            .in2(N__27755),
            .in3(N__27855),
            .lcout(\dron_frame_decoder_1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51421),
            .ce(),
            .sr(N__49526));
    defparam \dron_frame_decoder_1.state_3_LC_9_13_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_3_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_3_LC_9_13_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \dron_frame_decoder_1.state_3_LC_9_13_3  (
            .in0(N__27725),
            .in1(N__27964),
            .in2(N__27834),
            .in3(N__27854),
            .lcout(\dron_frame_decoder_1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51421),
            .ce(),
            .sr(N__49526));
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_13_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_data_valid_LC_9_13_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \dron_frame_decoder_1.source_data_valid_LC_9_13_4  (
            .in0(N__28054),
            .in1(N__32802),
            .in2(_gnd_net_),
            .in3(N__29212),
            .lcout(debug_CH1_0A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51421),
            .ce(),
            .sr(N__49526));
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_9_14_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI1H181_5_LC_9_14_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \dron_frame_decoder_1.state_RNI1H181_5_LC_9_14_0  (
            .in0(N__29204),
            .in1(N__27999),
            .in2(N__28121),
            .in3(N__49754),
            .lcout(\dron_frame_decoder_1.N_739_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_4_LC_9_14_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_4_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_4_LC_9_14_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_4_LC_9_14_1  (
            .in0(N__28000),
            .in1(N__28118),
            .in2(N__29222),
            .in3(N__27870),
            .lcout(\dron_frame_decoder_1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51406),
            .ce(),
            .sr(N__49534));
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_14_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_14_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__28114),
            .in2(_gnd_net_),
            .in3(N__29203),
            .lcout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4 ),
            .ltout(\dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_7_LC_9_14_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_7_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_7_LC_9_14_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \dron_frame_decoder_1.state_7_LC_9_14_4  (
            .in0(N__27872),
            .in1(_gnd_net_),
            .in2(N__28082),
            .in3(N__28077),
            .lcout(\dron_frame_decoder_1.stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51406),
            .ce(),
            .sr(N__49534));
    defparam \dron_frame_decoder_1.state_6_LC_9_14_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_6_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_6_LC_9_14_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \dron_frame_decoder_1.state_6_LC_9_14_5  (
            .in0(N__28058),
            .in1(N__29205),
            .in2(N__28079),
            .in3(N__27871),
            .lcout(\dron_frame_decoder_1.stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51406),
            .ce(),
            .sr(N__49534));
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_14_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNO_0_0_LC_9_14_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNO_0_0_LC_9_14_7  (
            .in0(N__28025),
            .in1(N__27976),
            .in2(N__28016),
            .in3(N__27963),
            .lcout(\dron_frame_decoder_1.N_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_5_LC_9_15_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_5_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_5_LC_9_15_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \dron_frame_decoder_1.state_5_LC_9_15_0  (
            .in0(N__29314),
            .in1(N__28001),
            .in2(_gnd_net_),
            .in3(N__27875),
            .lcout(\dron_frame_decoder_1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51391),
            .ce(),
            .sr(N__49541));
    defparam \dron_frame_decoder_1.state_1_LC_9_15_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_1_LC_9_15_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_1_LC_9_15_1  (
            .in0(N__27873),
            .in1(N__27980),
            .in2(N__27946),
            .in3(N__27965),
            .lcout(\dron_frame_decoder_1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51391),
            .ce(),
            .sr(N__49541));
    defparam \pid_side.pid_prereg_9_LC_9_15_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_9_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_9_LC_9_15_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_side.pid_prereg_9_LC_9_15_3  (
            .in0(N__27920),
            .in1(N__27908),
            .in2(N__50047),
            .in3(N__34559),
            .lcout(\pid_side.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51391),
            .ce(),
            .sr(N__49541));
    defparam \dron_frame_decoder_1.state_2_LC_9_15_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_2_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.state_2_LC_9_15_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \dron_frame_decoder_1.state_2_LC_9_15_5  (
            .in0(N__27874),
            .in1(N__27835),
            .in2(N__29243),
            .in3(N__29213),
            .lcout(\dron_frame_decoder_1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51391),
            .ce(),
            .sr(N__49541));
    defparam \pid_side.pid_prereg_8_LC_9_17_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_8_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_8_LC_9_17_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_side.pid_prereg_8_LC_9_17_0  (
            .in0(N__28457),
            .in1(N__28451),
            .in2(N__50022),
            .in3(N__34593),
            .lcout(\pid_side.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51365),
            .ce(),
            .sr(N__49555));
    defparam \pid_side.pid_prereg_11_LC_9_17_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_11_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_11_LC_9_17_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_11_LC_9_17_1  (
            .in0(N__28424),
            .in1(N__28394),
            .in2(N__50020),
            .in3(N__34431),
            .lcout(\pid_side.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51365),
            .ce(),
            .sr(N__49555));
    defparam \pid_side.pid_prereg_4_LC_9_17_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_4_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_4_LC_9_17_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_4_LC_9_17_5  (
            .in0(N__28388),
            .in1(N__28382),
            .in2(N__50021),
            .in3(N__38230),
            .lcout(\pid_side.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51365),
            .ce(),
            .sr(N__49555));
    defparam \pid_side.pid_prereg_6_LC_9_17_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_6_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_6_LC_9_17_6 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pid_side.pid_prereg_6_LC_9_17_6  (
            .in0(N__49985),
            .in1(N__28352),
            .in2(N__34204),
            .in3(N__28322),
            .lcout(\pid_side.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51365),
            .ce(),
            .sr(N__49555));
    defparam \pid_side.pid_prereg_19_LC_9_18_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_19_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_19_LC_9_18_0 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \pid_side.pid_prereg_19_LC_9_18_0  (
            .in0(N__28316),
            .in1(N__50027),
            .in2(N__28310),
            .in3(N__29344),
            .lcout(\pid_side.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51355),
            .ce(),
            .sr(N__49564));
    defparam \pid_side.pid_prereg_15_LC_9_18_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_15_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_15_LC_9_18_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_15_LC_9_18_1  (
            .in0(N__28274),
            .in1(N__28244),
            .in2(N__50044),
            .in3(N__34804),
            .lcout(\pid_side.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51355),
            .ce(),
            .sr(N__49564));
    defparam \pid_side.pid_prereg_14_LC_9_18_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_14_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_14_LC_9_18_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pid_side.pid_prereg_14_LC_9_18_2  (
            .in0(N__28238),
            .in1(N__28205),
            .in2(N__34790),
            .in3(N__50023),
            .lcout(\pid_side.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51355),
            .ce(),
            .sr(N__49564));
    defparam \pid_side.pid_prereg_17_LC_9_19_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_17_LC_9_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_17_LC_9_19_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_17_LC_9_19_0  (
            .in0(N__28199),
            .in1(N__28193),
            .in2(N__50046),
            .in3(N__29357),
            .lcout(\pid_side.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51345),
            .ce(),
            .sr(N__49572));
    defparam \pid_side.pid_prereg_20_LC_9_19_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_20_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_20_LC_9_19_1 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \pid_side.pid_prereg_20_LC_9_19_1  (
            .in0(N__50035),
            .in1(N__28154),
            .in2(N__29330),
            .in3(N__28148),
            .lcout(\pid_side.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51345),
            .ce(),
            .sr(N__49572));
    defparam \pid_side.pid_prereg_12_LC_9_19_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_12_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_12_LC_9_19_4 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_side.pid_prereg_12_LC_9_19_4  (
            .in0(N__28708),
            .in1(N__28676),
            .in2(N__50045),
            .in3(N__37841),
            .lcout(\pid_side.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51345),
            .ce(),
            .sr(N__49572));
    defparam \pid_side.pid_prereg_18_LC_9_19_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_18_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_18_LC_9_19_6 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_side.pid_prereg_18_LC_9_19_6  (
            .in0(N__50034),
            .in1(N__28670),
            .in2(N__28664),
            .in3(N__29369),
            .lcout(\pid_side.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51345),
            .ce(),
            .sr(N__49572));
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_9_20_0 .C_ON=1'b0;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_9_20_0 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_9_20_0  (
            .in0(N__28631),
            .in1(N__28613),
            .in2(_gnd_net_),
            .in3(N__28583),
            .lcout(\pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_8_l_ofx_LC_9_20_5 .C_ON=1'b0;
    defparam \pid_side.error_axb_8_l_ofx_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_8_l_ofx_LC_9_20_5 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \pid_side.error_axb_8_l_ofx_LC_9_20_5  (
            .in0(N__29300),
            .in1(_gnd_net_),
            .in2(N__28505),
            .in3(N__29542),
            .lcout(\pid_side.error_axb_8_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_axb_7_LC_9_20_6 .C_ON=1'b0;
    defparam \pid_side.error_axb_7_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_7_LC_9_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pid_side.error_axb_7_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__28501),
            .in2(_gnd_net_),
            .in3(N__29299),
            .lcout(\pid_side.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_2_LC_9_21_0 .C_ON=1'b0;
    defparam \pid_front.error_axb_2_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_2_LC_9_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_2_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28478),
            .lcout(\pid_front.error_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_9_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_9_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37113),
            .lcout(drone_H_disp_front_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51330),
            .ce(N__42509),
            .sr(N__49590));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_9_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_9_21_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__37022),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51330),
            .ce(N__42509),
            .sr(N__49590));
    defparam \pid_side.error_axb_1_LC_9_21_4 .C_ON=1'b0;
    defparam \pid_side.error_axb_1_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.error_axb_1_LC_9_21_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pid_side.error_axb_1_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__28472),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_RNO_LC_10_5_2 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.source_data_valid_esr_RNO_LC_10_5_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \pid_alt.source_data_valid_esr_RNO_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__31177),
            .in2(_gnd_net_),
            .in3(N__49776),
            .lcout(\pid_alt.state_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_data_valid_esr_LC_10_6_0 .C_ON=1'b0;
    defparam \pid_alt.source_data_valid_esr_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_data_valid_esr_LC_10_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_alt.source_data_valid_esr_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32018),
            .lcout(pid_altitude_dv),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51490),
            .ce(N__28811),
            .sr(N__49503));
    defparam \uart_pc.state_RNO_0_0_LC_10_7_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_0_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_0_LC_10_7_1 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_pc.state_RNO_0_0_LC_10_7_1  (
            .in0(N__32146),
            .in1(N__40705),
            .in2(_gnd_net_),
            .in3(N__49777),
            .lcout(),
            .ltout(\uart_pc.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_0_LC_10_7_2 .C_ON=1'b0;
    defparam \uart_pc.state_0_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_0_LC_10_7_2 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \uart_pc.state_0_LC_10_7_2  (
            .in0(N__29795),
            .in1(N__31100),
            .in2(N__28805),
            .in3(N__31265),
            .lcout(\uart_pc.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51479),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIMQ8T1_4_LC_10_8_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIMQ8T1_4_LC_10_8_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart_pc.state_RNIMQ8T1_4_LC_10_8_0  (
            .in0(N__48988),
            .in1(N__31261),
            .in2(N__31110),
            .in3(N__29789),
            .lcout(\uart_pc.N_143 ),
            .ltout(\uart_pc.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_3_LC_10_8_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_3_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_3_LC_10_8_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_pc.timer_Count_3_LC_10_8_1  (
            .in0(N__29696),
            .in1(N__29750),
            .in2(N__28802),
            .in3(N__48989),
            .lcout(\uart_pc.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51466),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_1_LC_10_8_2 .C_ON=1'b0;
    defparam \uart_drone.state_1_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_1_LC_10_8_2 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \uart_drone.state_1_LC_10_8_2  (
            .in0(N__29028),
            .in1(N__31010),
            .in2(N__30953),
            .in3(N__49780),
            .lcout(\uart_drone.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51466),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_10_8_4 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIPD2K1_2_LC_10_8_4 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \uart_pc.timer_Count_RNIPD2K1_2_LC_10_8_4  (
            .in0(N__31334),
            .in1(N__31306),
            .in2(N__31109),
            .in3(N__29788),
            .lcout(\uart_pc.data_rdyc_1 ),
            .ltout(\uart_pc.data_rdyc_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_10_8_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIMQ8T1_2_LC_10_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_pc.timer_Count_RNIMQ8T1_2_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28778),
            .in3(N__48987),
            .lcout(\uart_pc.timer_Count_RNIMQ8T1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_2_LC_10_8_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_2_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_2_LC_10_8_6 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \uart_drone.state_RNO_0_2_LC_10_8_6  (
            .in0(N__32958),
            .in1(N__31009),
            .in2(N__29030),
            .in3(N__49779),
            .lcout(),
            .ltout(\uart_drone.state_srsts_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_2_LC_10_8_7 .C_ON=1'b0;
    defparam \uart_drone.state_2_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_2_LC_10_8_7 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_drone.state_2_LC_10_8_7  (
            .in0(N__29029),
            .in1(N__33100),
            .in2(N__29012),
            .in3(N__33023),
            .lcout(\uart_drone.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51466),
            .ce(),
            .sr(_gnd_net_));
    defparam \scaler_4.source_data_1_esr_5_LC_10_9_0 .C_ON=1'b0;
    defparam \scaler_4.source_data_1_esr_5_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \scaler_4.source_data_1_esr_5_LC_10_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \scaler_4.source_data_1_esr_5_LC_10_9_0  (
            .in0(N__29009),
            .in1(N__28981),
            .in2(_gnd_net_),
            .in3(N__28948),
            .lcout(scaler_4_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51451),
            .ce(N__28912),
            .sr(N__49511));
    defparam \uart_pc.data_Aux_RNO_0_3_LC_10_9_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_3_LC_10_9_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_3_LC_10_9_2  (
            .in0(N__29998),
            .in1(N__30052),
            .in2(_gnd_net_),
            .in3(N__29952),
            .lcout(\uart_pc.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_9_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_6_LC_10_9_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_6_LC_10_9_5  (
            .in0(N__29953),
            .in1(_gnd_net_),
            .in2(N__30056),
            .in3(N__29999),
            .lcout(\uart_pc.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIEAGS_4_LC_10_9_6 .C_ON=1'b0;
    defparam \uart_pc.state_RNIEAGS_4_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIEAGS_4_LC_10_9_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_pc.state_RNIEAGS_4_LC_10_9_6  (
            .in0(N__29791),
            .in1(N__30140),
            .in2(_gnd_net_),
            .in3(N__49758),
            .lcout(\uart_pc.state_RNIEAGSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_2_LC_10_10_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_2_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_2_LC_10_10_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \uart_pc.data_Aux_2_LC_10_10_2  (
            .in0(N__40749),
            .in1(N__29039),
            .in2(N__28873),
            .in3(N__40694),
            .lcout(\uart_pc.data_AuxZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51436),
            .ce(),
            .sr(N__40528));
    defparam \uart_pc.data_Aux_1_LC_10_10_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_1_LC_10_10_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_1_LC_10_10_3 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_1_LC_10_10_3  (
            .in0(N__29900),
            .in1(N__40691),
            .in2(N__28852),
            .in3(N__40748),
            .lcout(\uart_pc.data_AuxZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51436),
            .ce(),
            .sr(N__40528));
    defparam \uart_pc.data_Aux_3_LC_10_10_5 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_3_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_3_LC_10_10_5 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_3_LC_10_10_5  (
            .in0(N__28835),
            .in1(N__40692),
            .in2(N__28828),
            .in3(N__40750),
            .lcout(\uart_pc.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51436),
            .ce(),
            .sr(N__40528));
    defparam \uart_pc.data_Aux_5_LC_10_10_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_5_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_5_LC_10_10_7 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_5_LC_10_10_7  (
            .in0(N__29045),
            .in1(N__40693),
            .in2(N__29074),
            .in3(N__40751),
            .lcout(\uart_pc.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51436),
            .ce(),
            .sr(N__40528));
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_11_2 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_4_LC_10_11_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_pc.data_Aux_RNO_0_4_LC_10_11_2  (
            .in0(N__29990),
            .in1(N__30038),
            .in2(_gnd_net_),
            .in3(N__29941),
            .lcout(\uart_pc.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_11_3 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_5_LC_10_11_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_5_LC_10_11_3  (
            .in0(N__29942),
            .in1(_gnd_net_),
            .in2(N__30046),
            .in3(N__29991),
            .lcout(\uart_pc.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_11_4 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_2_LC_10_11_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_pc.data_Aux_RNO_0_2_LC_10_11_4  (
            .in0(N__29989),
            .in1(N__30037),
            .in2(_gnd_net_),
            .in3(N__29940),
            .lcout(\uart_pc.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_esr_0_LC_10_12_0 .C_ON=1'b0;
    defparam \uart_drone.data_esr_0_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_0_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29893),
            .lcout(uart_drone_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51407),
            .ce(N__29284),
            .sr(N__29266));
    defparam \uart_drone.data_esr_2_LC_10_12_1 .C_ON=1'b0;
    defparam \uart_drone.data_esr_2_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_2_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_2_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30262),
            .lcout(uart_drone_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51407),
            .ce(N__29284),
            .sr(N__29266));
    defparam \uart_drone.data_esr_5_LC_10_12_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_5_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_5_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_5_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30224),
            .lcout(uart_drone_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51407),
            .ce(N__29284),
            .sr(N__29266));
    defparam \uart_drone.data_esr_7_LC_10_12_3 .C_ON=1'b0;
    defparam \uart_drone.data_esr_7_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_7_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_7_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30197),
            .lcout(uart_drone_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51407),
            .ce(N__29284),
            .sr(N__29266));
    defparam \uart_drone.data_esr_3_LC_10_13_2 .C_ON=1'b0;
    defparam \uart_drone.data_esr_3_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_3_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_3_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30248),
            .lcout(uart_drone_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51393),
            .ce(N__29291),
            .sr(N__29267));
    defparam \uart_drone.data_esr_4_LC_10_13_4 .C_ON=1'b0;
    defparam \uart_drone.data_esr_4_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_4_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_4_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30236),
            .lcout(uart_drone_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51393),
            .ce(N__29291),
            .sr(N__29267));
    defparam \uart_drone.data_esr_1_LC_10_13_5 .C_ON=1'b0;
    defparam \uart_drone.data_esr_1_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_1_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_1_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30275),
            .lcout(uart_drone_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51393),
            .ce(N__29291),
            .sr(N__29267));
    defparam \uart_drone.data_esr_6_LC_10_13_6 .C_ON=1'b0;
    defparam \uart_drone.data_esr_6_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_esr_6_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone.data_esr_6_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(uart_drone_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51393),
            .ce(N__29291),
            .sr(N__29267));
    defparam \pid_alt.source_pid_1_10_LC_10_14_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_10_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_10_LC_10_14_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_alt.source_pid_1_10_LC_10_14_0  (
            .in0(N__31854),
            .in1(N__32016),
            .in2(N__32492),
            .in3(N__29144),
            .lcout(throttle_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51379),
            .ce(),
            .sr(N__31774));
    defparam \pid_alt.source_pid_1_6_LC_10_14_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_6_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_6_LC_10_14_2 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_alt.source_pid_1_6_LC_10_14_2  (
            .in0(N__31855),
            .in1(N__29450),
            .in2(N__32672),
            .in3(N__32017),
            .lcout(throttle_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51379),
            .ce(),
            .sr(N__31774));
    defparam \pid_alt.source_pid_1_8_LC_10_14_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_8_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_8_LC_10_14_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_alt.source_pid_1_8_LC_10_14_5  (
            .in0(N__32015),
            .in1(N__31856),
            .in2(N__37794),
            .in3(N__29105),
            .lcout(throttle_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51379),
            .ce(),
            .sr(N__31774));
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_10_15_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI4N6K_2_LC_10_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \dron_frame_decoder_1.state_RNI4N6K_2_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__29238),
            .in2(_gnd_net_),
            .in3(N__29221),
            .lcout(\dron_frame_decoder_1.state_RNI4N6KZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_10_LC_10_16_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_10_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIT3KA1_10_LC_10_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIT3KA1_10_LC_10_16_1  (
            .in0(N__29139),
            .in1(N__30180),
            .in2(N__31807),
            .in3(N__29097),
            .lcout(),
            .ltout(\pid_alt.un1_reset_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_11_LC_10_16_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_11_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFQKS1_11_LC_10_16_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFQKS1_11_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__32046),
            .in2(N__29108),
            .in3(N__29448),
            .lcout(\pid_alt.N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNINTJA1_11_LC_10_16_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNINTJA1_11_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNINTJA1_11_LC_10_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_alt.pid_prereg_esr_RNINTJA1_11_LC_10_16_3  (
            .in0(N__32047),
            .in1(N__30181),
            .in2(N__31574),
            .in3(N__29098),
            .lcout(),
            .ltout(\pid_alt.un1_reset_i_a5_1_10_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIFBU82_6_LC_10_16_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIFBU82_6_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIFBU82_6_LC_10_16_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIFBU82_6_LC_10_16_4  (
            .in0(N__31803),
            .in1(N__30490),
            .in2(N__29453),
            .in3(N__29449),
            .lcout(\pid_alt.un1_reset_i_a5_1_10_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIEKJA1_1_LC_10_16_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIEKJA1_1_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIEKJA1_1_LC_10_16_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIEKJA1_1_LC_10_16_5  (
            .in0(N__30610),
            .in1(N__31495),
            .in2(N__30543),
            .in3(N__31528),
            .lcout(\pid_alt.un1_reset_i_a5_0_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNI8LUI1_6_LC_10_17_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNI8LUI1_6_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNI8LUI1_6_LC_10_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_RNI8LUI1_6_LC_10_17_0  (
            .in0(N__34586),
            .in1(N__34560),
            .in2(N__34200),
            .in3(N__34247),
            .lcout(\pid_side.un1_reset_i_a5_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_10_LC_10_17_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_10_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_10_LC_10_17_5 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \pid_side.pid_prereg_10_LC_10_17_5  (
            .in0(N__34249),
            .in1(N__29417),
            .in2(N__49978),
            .in3(N__29404),
            .lcout(\pid_side.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51347),
            .ce(),
            .sr(N__49556));
    defparam \pid_side.pid_prereg_RNIUDBG1_6_LC_10_17_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIUDBG1_6_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIUDBG1_6_LC_10_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_RNIUDBG1_6_LC_10_17_6  (
            .in0(N__34400),
            .in1(N__34193),
            .in2(N__34594),
            .in3(N__34561),
            .lcout(),
            .ltout(\pid_side.un1_reset_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNIHJND2_10_LC_10_17_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIHJND2_10_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIHJND2_10_LC_10_17_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \pid_side.pid_prereg_RNIHJND2_10_LC_10_17_7  (
            .in0(N__34248),
            .in1(_gnd_net_),
            .in2(N__29372),
            .in3(N__34430),
            .lcout(\pid_side.N_531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNIT3QQ1_17_LC_10_18_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIT3QQ1_17_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIT3QQ1_17_LC_10_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_RNIT3QQ1_17_LC_10_18_3  (
            .in0(N__29368),
            .in1(N__29356),
            .in2(N__29345),
            .in3(N__29326),
            .lcout(\pid_side.m7_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_10_20_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.state_RNI14DT_2_LC_10_20_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \dron_frame_decoder_1.state_RNI14DT_2_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__29315),
            .in2(_gnd_net_),
            .in3(N__49770),
            .lcout(\dron_frame_decoder_1.N_731_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_10_21_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_10_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37010),
            .lcout(drone_H_disp_side_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51317),
            .ce(N__29580),
            .sr(N__49591));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_10_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_10_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36934),
            .lcout(drone_H_disp_side_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51317),
            .ce(N__29580),
            .sr(N__49591));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_10_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_10_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36844),
            .lcout(drone_H_disp_side_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51317),
            .ce(N__29580),
            .sr(N__49591));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_10_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_10_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48433),
            .lcout(drone_H_disp_side_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51317),
            .ce(N__29580),
            .sr(N__49591));
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_22_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_22_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_side_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_3_LC_10_22_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_3_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_3_LC_10_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_3_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29510),
            .lcout(\pid_front.error_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_10_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_3_LC_10_23_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_3_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__39373),
            .in2(_gnd_net_),
            .in3(N__50798),
            .lcout(xy_kp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51310),
            .ce(N__39031),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.aux_3__0__0_LC_11_4_0 .C_ON=1'b0;
    defparam \uart_drone_sync.aux_3__0__0_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.aux_3__0__0_LC_11_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.aux_3__0__0_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29465),
            .lcout(\uart_drone_sync.aux_3__0__0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51501),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_2_LC_11_6_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_2_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_2_LC_11_6_3 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \uart_pc.timer_Count_2_LC_11_6_3  (
            .in0(N__29759),
            .in1(N__48910),
            .in2(N__29692),
            .in3(N__29825),
            .lcout(\uart_pc.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51480),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_7_0 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIRP8S_1_LC_11_7_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_pc.timer_Count_RNIRP8S_1_LC_11_7_0  (
            .in0(N__29717),
            .in1(N__29647),
            .in2(N__29722),
            .in3(_gnd_net_),
            .lcout(\uart_pc.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\uart_pc.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_7_1 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_2_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_2_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__31332),
            .in2(_gnd_net_),
            .in3(N__29753),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_7_2 .C_ON=1'b1;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_3_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_pc.timer_Count_RNO_0_3_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__31303),
            .in2(_gnd_net_),
            .in3(N__29744),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_pc.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_pc.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_7_3 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_4_LC_11_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_4_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__31098),
            .in2(_gnd_net_),
            .in3(N__29741),
            .lcout(\uart_pc.timer_Count_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_7_4 .C_ON=1'b0;
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIGRIF1_2_LC_11_7_4 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \uart_pc.state_RNIGRIF1_2_LC_11_7_4  (
            .in0(N__31099),
            .in1(N__31304),
            .in2(N__30152),
            .in3(N__32172),
            .lcout(\uart_pc.timer_Count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_4_LC_11_7_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_4_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_4_LC_11_7_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_pc.timer_Count_4_LC_11_7_5  (
            .in0(N__29738),
            .in1(N__29820),
            .in2(N__29690),
            .in3(N__48970),
            .lcout(\uart_pc.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51467),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_0_LC_11_7_7 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_0_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_0_LC_11_7_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_pc.timer_Count_0_LC_11_7_7  (
            .in0(N__29721),
            .in1(N__29819),
            .in2(N__29689),
            .in3(N__48969),
            .lcout(\uart_pc.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51467),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIBLRB2_4_LC_11_8_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNIBLRB2_4_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIBLRB2_4_LC_11_8_0 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \uart_pc.state_RNIBLRB2_4_LC_11_8_0  (
            .in0(N__31260),
            .in1(N__30139),
            .in2(N__29732),
            .in3(N__29790),
            .lcout(\uart_pc.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_8_1 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNO_0_1_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_pc.timer_Count_RNO_0_1_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__29723),
            .in2(_gnd_net_),
            .in3(N__29648),
            .lcout(),
            .ltout(\uart_pc.timer_Count_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_1_LC_11_8_2 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_1_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.timer_Count_1_LC_11_8_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.timer_Count_1_LC_11_8_2  (
            .in0(N__48967),
            .in1(N__29691),
            .in2(N__29651),
            .in3(N__29821),
            .lcout(\uart_pc.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51452),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_11_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIDGR31_2_LC_11_8_3 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \uart_drone.timer_Count_RNIDGR31_2_LC_11_8_3  (
            .in0(N__33153),
            .in1(N__33004),
            .in2(N__33091),
            .in3(N__32463),
            .lcout(\uart_drone.data_rdyc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone_sync.Q_0__0_LC_11_8_5 .C_ON=1'b0;
    defparam \uart_drone_sync.Q_0__0_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone_sync.Q_0__0_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_drone_sync.Q_0__0_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29849),
            .lcout(debug_CH0_16A_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51452),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI40411_2_LC_11_8_6 .C_ON=1'b0;
    defparam \uart_drone.state_RNI40411_2_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI40411_2_LC_11_8_6 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \uart_drone.state_RNI40411_2_LC_11_8_6  (
            .in0(N__33005),
            .in1(N__32912),
            .in2(N__32967),
            .in3(N__33075),
            .lcout(\uart_drone.timer_Count_0_sqmuxa ),
            .ltout(\uart_drone.timer_Count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_3_LC_11_8_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_3_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_3_LC_11_8_7 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_3_LC_11_8_7  (
            .in0(N__32438),
            .in1(N__32342),
            .in2(N__29840),
            .in3(N__48968),
            .lcout(\uart_drone.timer_CountZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51452),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNO_0_3_LC_11_9_0 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_3_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_3_LC_11_9_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_pc.state_RNO_0_3_LC_11_9_0  (
            .in0(N__30137),
            .in1(N__31108),
            .in2(N__32189),
            .in3(N__31293),
            .lcout(),
            .ltout(\uart_pc.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_3_LC_11_9_1 .C_ON=1'b0;
    defparam \uart_pc.state_3_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_3_LC_11_9_1 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \uart_pc.state_3_LC_11_9_1  (
            .in0(N__48966),
            .in1(N__29834),
            .in2(N__29837),
            .in3(N__32188),
            .lcout(\uart_pc.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51437),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_11_9_5 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNI5UFA2_3_LC_11_9_5 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \uart_pc.timer_Count_RNI5UFA2_3_LC_11_9_5  (
            .in0(N__31292),
            .in1(N__40575),
            .in2(N__31112),
            .in3(_gnd_net_),
            .lcout(\uart_pc.N_144_1 ),
            .ltout(\uart_pc.N_144_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_4_LC_11_9_6 .C_ON=1'b0;
    defparam \uart_pc.state_4_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_4_LC_11_9_6 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \uart_pc.state_4_LC_11_9_6  (
            .in0(N__30138),
            .in1(N__48965),
            .in2(N__29828),
            .in3(N__29818),
            .lcout(\uart_pc.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51437),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIITIF1_4_LC_11_9_7 .C_ON=1'b0;
    defparam \uart_pc.state_RNIITIF1_4_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIITIF1_4_LC_11_9_7 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \uart_pc.state_RNIITIF1_4_LC_11_9_7  (
            .in0(N__31291),
            .in1(N__29787),
            .in2(N__31111),
            .in3(N__30136),
            .lcout(\uart_pc.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_11_10_0 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNI4U6E1_2_LC_11_10_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_pc.bit_Count_RNI4U6E1_2_LC_11_10_0  (
            .in0(N__29983),
            .in1(N__30030),
            .in2(_gnd_net_),
            .in3(N__29933),
            .lcout(\uart_pc.N_152 ),
            .ltout(\uart_pc.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_RNIUPE73_3_LC_11_10_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNIUPE73_3_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNIUPE73_3_LC_11_10_1 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \uart_pc.state_RNIUPE73_3_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__30088),
            .in2(N__30155),
            .in3(N__30144),
            .lcout(\uart_pc.un1_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_9_LC_11_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_9_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_9_LC_11_11_0 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_9_LC_11_11_0  (
            .in0(N__31414),
            .in1(N__31391),
            .in2(N__46170),
            .in3(N__35641),
            .lcout(\ppm_encoder_1.throttleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51408),
            .ce(),
            .sr(N__49522));
    defparam \uart_pc.bit_Count_0_LC_11_11_2 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_0_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_0_LC_11_11_2 .LUT_INIT=16'b0101001001010000;
    LogicCell40 \uart_pc.bit_Count_0_LC_11_11_2  (
            .in0(N__30097),
            .in1(N__40585),
            .in2(N__29951),
            .in3(N__30151),
            .lcout(\uart_pc.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51408),
            .ce(),
            .sr(N__49522));
    defparam \uart_pc.bit_Count_RNO_0_2_LC_11_11_3 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_pc.bit_Count_RNO_0_2_LC_11_11_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.bit_Count_RNO_0_2_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__29936),
            .in2(_gnd_net_),
            .in3(N__30096),
            .lcout(),
            .ltout(\uart_pc.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.bit_Count_2_LC_11_11_4 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_2_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_2_LC_11_11_4 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uart_pc.bit_Count_2_LC_11_11_4  (
            .in0(N__30077),
            .in1(N__29988),
            .in2(N__30101),
            .in3(N__30036),
            .lcout(\uart_pc.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51408),
            .ce(),
            .sr(N__49522));
    defparam \uart_pc.bit_Count_1_LC_11_11_5 .C_ON=1'b0;
    defparam \uart_pc.bit_Count_1_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_pc.bit_Count_1_LC_11_11_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_pc.bit_Count_1_LC_11_11_5  (
            .in0(N__29954),
            .in1(N__30098),
            .in2(N__30045),
            .in3(N__30076),
            .lcout(\uart_pc.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51408),
            .ce(),
            .sr(N__49522));
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_11_6 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_0_LC_11_11_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_pc.data_Aux_RNO_0_0_LC_11_11_6  (
            .in0(N__29934),
            .in1(N__29984),
            .in2(_gnd_net_),
            .in3(N__30031),
            .lcout(\uart_pc.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_RNO_0_1_LC_11_11_7 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_pc.data_Aux_RNO_0_1_LC_11_11_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uart_pc.data_Aux_RNO_0_1_LC_11_11_7  (
            .in0(N__30032),
            .in1(_gnd_net_),
            .in2(N__29997),
            .in3(N__29935),
            .lcout(\uart_pc.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_0_LC_11_12_0 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_0_LC_11_12_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uart_drone.data_Aux_0_LC_11_12_0  (
            .in0(N__31021),
            .in1(N__30161),
            .in2(N__29894),
            .in3(N__31238),
            .lcout(\uart_drone.data_AuxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_1_LC_11_12_1 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_1_LC_11_12_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_1_LC_11_12_1  (
            .in0(N__31234),
            .in1(N__30274),
            .in2(N__31047),
            .in3(N__30335),
            .lcout(\uart_drone.data_AuxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_2_LC_11_12_2 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_2_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_2_LC_11_12_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_2_LC_11_12_2  (
            .in0(N__31586),
            .in1(N__31025),
            .in2(N__30263),
            .in3(N__31239),
            .lcout(\uart_drone.data_AuxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_3_LC_11_12_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_3_LC_11_12_3 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_3_LC_11_12_3  (
            .in0(N__31235),
            .in1(N__30247),
            .in2(N__31048),
            .in3(N__30326),
            .lcout(\uart_drone.data_AuxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_4_LC_11_12_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_4_LC_11_12_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uart_drone.data_Aux_4_LC_11_12_4  (
            .in0(N__30320),
            .in1(N__30235),
            .in2(N__31046),
            .in3(N__31240),
            .lcout(\uart_drone.data_AuxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_5_LC_11_12_5 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_5_LC_11_12_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_5_LC_11_12_5  (
            .in0(N__31236),
            .in1(N__30223),
            .in2(N__31049),
            .in3(N__30698),
            .lcout(\uart_drone.data_AuxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_6_LC_11_12_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_6_LC_11_12_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_drone.data_Aux_6_LC_11_12_6  (
            .in0(N__30560),
            .in1(N__31026),
            .in2(N__30212),
            .in3(N__31241),
            .lcout(\uart_drone.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \uart_drone.data_Aux_7_LC_11_12_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_7_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.data_Aux_7_LC_11_12_7 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_drone.data_Aux_7_LC_11_12_7  (
            .in0(N__31237),
            .in1(N__30196),
            .in2(N__31050),
            .in3(N__32096),
            .lcout(\uart_drone.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51394),
            .ce(),
            .sr(N__33122));
    defparam \pid_alt.source_pid_1_9_LC_11_13_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_9_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_9_LC_11_13_1 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_alt.source_pid_1_9_LC_11_13_1  (
            .in0(N__31853),
            .in1(N__32030),
            .in2(N__31415),
            .in3(N__30185),
            .lcout(throttle_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51380),
            .ce(),
            .sr(N__31778));
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_13_3 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_0_LC_11_13_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_drone.data_Aux_RNO_0_0_LC_11_13_3  (
            .in0(N__31724),
            .in1(N__31654),
            .in2(_gnd_net_),
            .in3(N__34535),
            .lcout(\uart_drone.data_Auxce_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_13_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_1_LC_11_13_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uart_drone.data_Aux_RNO_0_1_LC_11_13_4  (
            .in0(N__34537),
            .in1(_gnd_net_),
            .in2(N__31663),
            .in3(N__31725),
            .lcout(\uart_drone.data_Auxce_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_3_LC_11_13_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_3_LC_11_13_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_3_LC_11_13_6  (
            .in0(N__34538),
            .in1(_gnd_net_),
            .in2(N__31664),
            .in3(N__31726),
            .lcout(\uart_drone.data_Auxce_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_13_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_4_LC_11_13_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_4_LC_11_13_7  (
            .in0(N__31727),
            .in1(N__31661),
            .in2(_gnd_net_),
            .in3(N__34536),
            .lcout(\uart_drone.data_Auxce_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_esr_13_LC_11_14_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_13_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_13_LC_11_14_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.source_pid_1_esr_13_LC_11_14_2  (
            .in0(N__30410),
            .in1(N__30451),
            .in2(_gnd_net_),
            .in3(N__30505),
            .lcout(throttle_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51367),
            .ce(N__31598),
            .sr(N__31769));
    defparam \pid_alt.source_pid_1_esr_12_LC_11_14_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_12_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_12_LC_11_14_3 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \pid_alt.source_pid_1_esr_12_LC_11_14_3  (
            .in0(N__30506),
            .in1(N__30548),
            .in2(N__30460),
            .in3(N__30409),
            .lcout(throttle_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51367),
            .ce(N__31598),
            .sr(N__31769));
    defparam \pid_alt.source_pid_1_esr_5_LC_11_14_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_5_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_5_LC_11_14_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \pid_alt.source_pid_1_esr_5_LC_11_14_5  (
            .in0(N__31852),
            .in1(_gnd_net_),
            .in2(N__30674),
            .in3(N__30658),
            .lcout(throttle_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51367),
            .ce(N__31598),
            .sr(N__31769));
    defparam \pid_alt.source_pid_1_esr_4_LC_11_14_6 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_esr_4_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_esr_4_LC_11_14_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pid_alt.source_pid_1_esr_4_LC_11_14_6  (
            .in0(N__30659),
            .in1(N__31851),
            .in2(N__30614),
            .in3(N__30670),
            .lcout(throttle_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51367),
            .ce(N__31598),
            .sr(N__31769));
    defparam \pid_alt.pid_prereg_esr_RNIG5AU_0_LC_11_15_2 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIG5AU_0_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIG5AU_0_LC_11_15_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIG5AU_0_LC_11_15_2  (
            .in0(N__30499),
            .in1(N__30638),
            .in2(_gnd_net_),
            .in3(N__31563),
            .lcout(),
            .ltout(\pid_alt.un1_reset_i_a5_0_6_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI2R305_0_LC_11_15_3 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI2R305_0_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI2R305_0_LC_11_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI2R305_0_LC_11_15_3  (
            .in0(N__30314),
            .in1(N__30308),
            .in2(N__30278),
            .in3(N__30685),
            .lcout(),
            .ltout(\pid_alt.un1_reset_i_a5_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI1RJPB_10_LC_11_15_4 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI1RJPB_10_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI1RJPB_10_LC_11_15_4 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI1RJPB_10_LC_11_15_4  (
            .in0(N__30719),
            .in1(N__30713),
            .in2(N__30704),
            .in3(N__30399),
            .lcout(),
            .ltout(\pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI65QMC_24_LC_11_15_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI65QMC_24_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI65QMC_24_LC_11_15_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI65QMC_24_LC_11_15_5  (
            .in0(N__30459),
            .in1(N__32023),
            .in2(N__30701),
            .in3(N__48961),
            .lcout(\pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_15_6 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_5_LC_11_15_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_5_LC_11_15_6  (
            .in0(N__31662),
            .in1(N__34525),
            .in2(_gnd_net_),
            .in3(N__31714),
            .lcout(\uart_drone.data_Auxce_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIJ6482_24_LC_11_16_0 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIJ6482_24_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIJ6482_24_LC_11_16_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIJ6482_24_LC_11_16_0  (
            .in0(N__30492),
            .in1(N__30458),
            .in2(_gnd_net_),
            .in3(N__30686),
            .lcout(\pid_alt.N_535 ),
            .ltout(\pid_alt.N_535_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNI70AB5_4_LC_11_16_1 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNI70AB5_4_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNI70AB5_4_LC_11_16_1 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \pid_alt.pid_prereg_esr_RNI70AB5_4_LC_11_16_1  (
            .in0(N__31833),
            .in1(N__30657),
            .in2(N__30617),
            .in3(N__30609),
            .lcout(\pid_alt.N_472_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_11_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_ctle_14_LC_11_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_ctle_14_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__46157),
            .in2(_gnd_net_),
            .in3(N__49760),
            .lcout(\ppm_encoder_1.pid_altitude_dv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_16_4 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_6_LC_11_16_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_drone.data_Aux_RNO_0_6_LC_11_16_4  (
            .in0(N__31640),
            .in1(N__31703),
            .in2(_gnd_net_),
            .in3(N__34514),
            .lcout(\uart_drone.data_Auxce_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_11_16_5 .C_ON=1'b0;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_11_16_5 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_11_16_5  (
            .in0(N__30536),
            .in1(N__30491),
            .in2(N__30461),
            .in3(N__30408),
            .lcout(\pid_alt.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_7_LC_11_17_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_7_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_7_LC_11_17_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_side.pid_prereg_7_LC_11_17_0  (
            .in0(N__30377),
            .in1(N__30368),
            .in2(N__49977),
            .in3(N__34401),
            .lcout(\pid_side.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \pid_side.state_0_LC_11_17_1 .C_ON=1'b0;
    defparam \pid_side.state_0_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_0_LC_11_17_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.state_0_LC_11_17_1  (
            .in0(N__49926),
            .in1(N__32831),
            .in2(_gnd_net_),
            .in3(N__35867),
            .lcout(\pid_side.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \pid_side.pid_prereg_3_LC_11_17_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_3_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_3_LC_11_17_2 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \pid_side.pid_prereg_3_LC_11_17_2  (
            .in0(N__49930),
            .in1(N__50114),
            .in2(N__35787),
            .in3(N__30932),
            .lcout(\pid_side.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \pid_side.pid_prereg_16_LC_11_17_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_16_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_16_LC_11_17_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_16_LC_11_17_4  (
            .in0(N__30923),
            .in1(N__30890),
            .in2(N__49975),
            .in3(N__34753),
            .lcout(\pid_side.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \pid_side.pid_prereg_5_LC_11_17_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_5_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_5_LC_11_17_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_side.pid_prereg_5_LC_11_17_6  (
            .in0(N__30878),
            .in1(N__30869),
            .in2(N__49976),
            .in3(N__38117),
            .lcout(\pid_side.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \ppm_encoder_1.rudder_6_LC_11_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_6_LC_11_17_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_6_LC_11_17_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.rudder_6_LC_11_17_7  (
            .in0(N__46194),
            .in1(N__31211),
            .in2(_gnd_net_),
            .in3(N__38775),
            .lcout(\ppm_encoder_1.rudderZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51338),
            .ce(),
            .sr(N__49565));
    defparam \pid_side.state_1_LC_11_19_7 .C_ON=1'b0;
    defparam \pid_side.state_1_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.state_1_LC_11_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pid_side.state_1_LC_11_19_7  (
            .in0(N__49974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_side.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51323),
            .ce(),
            .sr(N__49583));
    defparam \pid_side.pid_prereg_13_LC_11_20_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_13_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_13_LC_11_20_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_side.pid_prereg_13_LC_11_20_1  (
            .in0(N__30839),
            .in1(N__30809),
            .in2(N__50039),
            .in3(N__38284),
            .lcout(\pid_side.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51318),
            .ce(),
            .sr(N__49592));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_11_21_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_1_LC_11_21_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_1_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__39641),
            .in2(_gnd_net_),
            .in3(N__50799),
            .lcout(xy_kp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51314),
            .ce(N__39027),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_11_21_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_11_21_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_e_0_6_LC_11_21_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_e_0_6_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__40013),
            .in2(_gnd_net_),
            .in3(N__50800),
            .lcout(xy_kp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51314),
            .ce(N__39027),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_1_LC_11_22_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_1_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_1_LC_11_22_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_front.pid_prereg_1_LC_11_22_1  (
            .in0(N__42802),
            .in1(N__48785),
            .in2(_gnd_net_),
            .in3(N__32216),
            .lcout(\pid_front.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51311),
            .ce(),
            .sr(N__49600));
    defparam \pid_front.state_RNIPKTD_0_LC_11_23_0 .C_ON=1'b0;
    defparam \pid_front.state_RNIPKTD_0_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIPKTD_0_LC_11_23_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \pid_front.state_RNIPKTD_0_LC_11_23_0  (
            .in0(N__42726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49769),
            .lcout(\pid_front.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.state_RNIH1EN_0_LC_12_1_3 .C_ON=1'b0;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIH1EN_0_LC_12_1_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIH1EN_0_LC_12_1_3  (
            .in0(_gnd_net_),
            .in1(N__31163),
            .in2(_gnd_net_),
            .in3(N__49753),
            .lcout(\pid_alt.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_2_LC_12_7_0 .C_ON=1'b0;
    defparam \uart_pc.state_2_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_2_LC_12_7_0 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \uart_pc.state_2_LC_12_7_0  (
            .in0(N__31101),
            .in1(N__31310),
            .in2(N__32135),
            .in3(N__32156),
            .lcout(\uart_pc.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_0_LC_12_7_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_0_LC_12_7_1 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uart_drone.state_RNO_0_0_LC_12_7_1  (
            .in0(N__30943),
            .in1(N__31011),
            .in2(_gnd_net_),
            .in3(N__49778),
            .lcout(),
            .ltout(\uart_drone.state_srsts_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_0_LC_12_7_2 .C_ON=1'b0;
    defparam \uart_drone.state_0_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_0_LC_12_7_2 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \uart_drone.state_0_LC_12_7_2  (
            .in0(N__32362),
            .in1(N__33081),
            .in2(N__30956),
            .in3(N__33171),
            .lcout(\uart_drone.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_4_LC_12_7_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_4_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_4_LC_12_7_7 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \uart_drone.timer_Count_4_LC_12_7_7  (
            .in0(N__48977),
            .in1(N__32423),
            .in2(N__32417),
            .in3(N__32339),
            .lcout(\uart_drone.timer_CountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_2_LC_12_8_1 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_2_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_2_LC_12_8_1 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \uart_drone.timer_Count_2_LC_12_8_1  (
            .in0(N__32447),
            .in1(N__32335),
            .in2(N__32415),
            .in3(N__48980),
            .lcout(\uart_drone.timer_CountZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51435),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_1_LC_12_8_2 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_1_LC_12_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_drone.timer_Count_RNO_0_1_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__32385),
            .in2(_gnd_net_),
            .in3(N__32117),
            .lcout(),
            .ltout(\uart_drone.timer_Count_RNO_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_1_LC_12_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_1_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_1_LC_12_8_3 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \uart_drone.timer_Count_1_LC_12_8_3  (
            .in0(N__32405),
            .in1(N__32334),
            .in2(N__31337),
            .in3(N__48979),
            .lcout(\uart_drone.timer_CountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51435),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_8_6 .C_ON=1'b0;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_pc.timer_Count_RNIVT8S_2_LC_12_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_pc.timer_Count_RNIVT8S_2_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__31333),
            .in2(_gnd_net_),
            .in3(N__31305),
            .lcout(\uart_pc.N_126_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_12_8_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI9E9J_2_LC_12_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_drone.timer_Count_RNI9E9J_2_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__33006),
            .in2(_gnd_net_),
            .in3(N__32464),
            .lcout(\uart_drone.N_126_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_4_LC_12_9_4 .C_ON=1'b0;
    defparam \uart_drone.state_4_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_4_LC_12_9_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \uart_drone.state_4_LC_12_9_4  (
            .in0(N__32908),
            .in1(N__32936),
            .in2(N__32341),
            .in3(N__48978),
            .lcout(\uart_drone.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51422),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI9ADK1_4_LC_12_9_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNI9ADK1_4_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI9ADK1_4_LC_12_9_7 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \uart_drone.state_RNI9ADK1_4_LC_12_9_7  (
            .in0(N__32361),
            .in1(N__32907),
            .in2(N__32105),
            .in3(N__33158),
            .lcout(\uart_drone.un1_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__31204),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\ppm_encoder_1.un1_rudder_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__32245),
            .in2(_gnd_net_),
            .in3(N__31187),
            .lcout(\ppm_encoder_1.un1_rudder_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_6 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_10_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__32269),
            .in2(_gnd_net_),
            .in3(N__31184),
            .lcout(\ppm_encoder_1.un1_rudder_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_7 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_10_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__34978),
            .in2(_gnd_net_),
            .in3(N__31181),
            .lcout(\ppm_encoder_1.un1_rudder_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_8 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_10_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34045),
            .in3(N__31370),
            .lcout(\ppm_encoder_1.un1_rudder_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_9 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_10_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__32638),
            .in2(_gnd_net_),
            .in3(N__31367),
            .lcout(\ppm_encoder_1.un1_rudder_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_10 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_10_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__32299),
            .in2(_gnd_net_),
            .in3(N__31364),
            .lcout(\ppm_encoder_1.un1_rudder_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_11 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_10_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__32584),
            .in2(N__48043),
            .in3(N__31361),
            .lcout(\ppm_encoder_1.un1_rudder_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_rudder_cry_12 ),
            .carryout(\ppm_encoder_1.un1_rudder_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_14_LC_12_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.rudder_esr_14_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__31358),
            .in2(_gnd_net_),
            .in3(N__31349),
            .lcout(\ppm_encoder_1.rudderZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51392),
            .ce(N__36693),
            .sr(N__49527));
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_12_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__44034),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_12_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__35517),
            .in2(N__48040),
            .in3(N__31346),
            .lcout(\ppm_encoder_1.un1_throttle_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_0 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_12_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__32544),
            .in2(_gnd_net_),
            .in3(N__31343),
            .lcout(\ppm_encoder_1.un1_throttle_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_1 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_12_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__32733),
            .in2(N__48041),
            .in3(N__31340),
            .lcout(\ppm_encoder_1.un1_throttle_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_2 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_12_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__46438),
            .in2(_gnd_net_),
            .in3(N__31430),
            .lcout(\ppm_encoder_1.un1_throttle_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_3 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_12_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32701),
            .in3(N__31427),
            .lcout(\ppm_encoder_1.un1_throttle_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_4 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_12_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__32670),
            .in2(N__48042),
            .in3(N__31424),
            .lcout(\ppm_encoder_1.un1_throttle_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_5 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_12_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(N__45534),
            .in2(_gnd_net_),
            .in3(N__31421),
            .lcout(\ppm_encoder_1.un1_throttle_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_6 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_13_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__37795),
            .in2(_gnd_net_),
            .in3(N__31418),
            .lcout(\ppm_encoder_1.un1_throttle_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\ppm_encoder_1.un1_throttle_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_13_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__31407),
            .in2(_gnd_net_),
            .in3(N__31382),
            .lcout(\ppm_encoder_1.un1_throttle_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_8 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_13_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__32490),
            .in2(_gnd_net_),
            .in3(N__31379),
            .lcout(\ppm_encoder_1.un1_throttle_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_9 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_13_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__32616),
            .in2(_gnd_net_),
            .in3(N__31376),
            .lcout(\ppm_encoder_1.un1_throttle_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_10 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_13_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__32752),
            .in2(_gnd_net_),
            .in3(N__31373),
            .lcout(\ppm_encoder_1.un1_throttle_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_11 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_13_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__47885),
            .in2(N__41512),
            .in3(N__31604),
            .lcout(\ppm_encoder_1.un1_throttle_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_throttle_cry_12 ),
            .carryout(\ppm_encoder_1.un1_throttle_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_esr_14_LC_12_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.throttle_esr_14_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31601),
            .lcout(\ppm_encoder_1.throttleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51366),
            .ce(N__36698),
            .sr(N__49542));
    defparam \pid_alt.state_RNIRQ15D_1_LC_12_14_4 .C_ON=1'b0;
    defparam \pid_alt.state_RNIRQ15D_1_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \pid_alt.state_RNIRQ15D_1_LC_12_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_alt.state_RNIRQ15D_1_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__32014),
            .in2(_gnd_net_),
            .in3(N__31768),
            .lcout(\pid_alt.N_72_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_14_5  (
            .in0(N__46667),
            .in1(N__31742),
            .in2(_gnd_net_),
            .in3(N__38657),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_14_7 .C_ON=1'b0;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.data_Aux_RNO_0_2_LC_12_14_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_drone.data_Aux_RNO_0_2_LC_12_14_7  (
            .in0(N__31641),
            .in1(N__31713),
            .in2(_gnd_net_),
            .in3(N__34517),
            .lcout(\uart_drone.data_Auxce_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.source_pid_1_0_LC_12_15_0 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_0_LC_12_15_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \pid_alt.source_pid_1_0_LC_12_15_0  (
            .in0(N__31442),
            .in1(N__31570),
            .in2(N__44038),
            .in3(N__32028),
            .lcout(throttle_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \pid_alt.source_pid_1_1_LC_12_15_1 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_1_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_1_LC_12_15_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \pid_alt.source_pid_1_1_LC_12_15_1  (
            .in0(N__32025),
            .in1(N__31443),
            .in2(N__31535),
            .in3(N__35521),
            .lcout(throttle_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \pid_alt.source_pid_1_2_LC_12_15_2 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_2_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_2_LC_12_15_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \pid_alt.source_pid_1_2_LC_12_15_2  (
            .in0(N__31444),
            .in1(N__31499),
            .in2(N__32546),
            .in3(N__32029),
            .lcout(throttle_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \pid_alt.source_pid_1_3_LC_12_15_3 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_3_LC_12_15_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \pid_alt.source_pid_1_3_LC_12_15_3  (
            .in0(N__32026),
            .in1(N__31465),
            .in2(N__32735),
            .in3(N__31445),
            .lcout(throttle_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \pid_alt.source_pid_1_11_LC_12_15_5 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_11_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_11_LC_12_15_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_alt.source_pid_1_11_LC_12_15_5  (
            .in0(N__32024),
            .in1(N__31842),
            .in2(N__32618),
            .in3(N__32054),
            .lcout(throttle_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \pid_alt.source_pid_1_7_LC_12_15_7 .C_ON=1'b0;
    defparam \pid_alt.source_pid_1_7_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_alt.source_pid_1_7_LC_12_15_7 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_alt.source_pid_1_7_LC_12_15_7  (
            .in0(N__32027),
            .in1(N__31843),
            .in2(N__45544),
            .in3(N__31808),
            .lcout(throttle_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51346),
            .ce(),
            .sr(N__31770));
    defparam \uart_drone.state_RNI62411_4_LC_12_16_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNI62411_4_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI62411_4_LC_12_16_0 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \uart_drone.state_RNI62411_4_LC_12_16_0  (
            .in0(N__33095),
            .in1(N__33027),
            .in2(N__32896),
            .in3(N__33172),
            .lcout(\uart_drone.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_12_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_12_16_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_12_16_5  (
            .in0(N__39152),
            .in1(N__38806),
            .in2(_gnd_net_),
            .in3(N__46788),
            .lcout(\ppm_encoder_1.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_12_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_12_16_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_12_16_6  (
            .in0(N__46787),
            .in1(N__35621),
            .in2(_gnd_net_),
            .in3(N__38429),
            .lcout(\ppm_encoder_1.N_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNI63LK2_3_LC_12_17_1 .C_ON=1'b0;
    defparam \uart_drone.state_RNI63LK2_3_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNI63LK2_3_LC_12_17_1 .LUT_INIT=16'b1100010011000100;
    LogicCell40 \uart_drone.state_RNI63LK2_3_LC_12_17_1  (
            .in0(N__32897),
            .in1(N__34466),
            .in2(N__32092),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_7_0 ),
            .ltout(\uart_drone.un1_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_1_LC_12_17_2 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_1_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_1_LC_12_17_2 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uart_drone.bit_Count_1_LC_12_17_2  (
            .in0(N__34468),
            .in1(N__34516),
            .in2(N__31733),
            .in3(N__31701),
            .lcout(\uart_drone.bit_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51331),
            .ce(),
            .sr(N__49573));
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_17_3 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNIJOJC1_2_LC_12_17_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.bit_Count_RNIJOJC1_2_LC_12_17_3  (
            .in0(N__31700),
            .in1(N__31626),
            .in2(_gnd_net_),
            .in3(N__34502),
            .lcout(\uart_drone.N_152 ),
            .ltout(\uart_drone.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_0_LC_12_17_4 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_0_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_0_LC_12_17_4 .LUT_INIT=16'b0100011001000100;
    LogicCell40 \uart_drone.bit_Count_0_LC_12_17_4  (
            .in0(N__34467),
            .in1(N__34515),
            .in2(N__31730),
            .in3(N__32898),
            .lcout(\uart_drone.bit_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51331),
            .ce(),
            .sr(N__49573));
    defparam \uart_drone.bit_Count_2_LC_12_17_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_2_LC_12_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_drone.bit_Count_2_LC_12_17_5 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \uart_drone.bit_Count_2_LC_12_17_5  (
            .in0(N__31702),
            .in1(N__31627),
            .in2(N__31673),
            .in3(N__34448),
            .lcout(\uart_drone.bit_CountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51331),
            .ce(),
            .sr(N__49573));
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_17_7 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNIU8TV1_3_LC_12_17_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_drone.timer_Count_RNIU8TV1_3_LC_12_17_7  (
            .in0(N__32085),
            .in1(N__33096),
            .in2(_gnd_net_),
            .in3(N__33028),
            .lcout(\uart_drone.N_144_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_0_LC_12_18_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_0_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_0_LC_12_18_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_front.source_pid_1_0_LC_12_18_1  (
            .in0(N__32066),
            .in1(N__33679),
            .in2(N__35731),
            .in3(N__36235),
            .lcout(front_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51322),
            .ce(),
            .sr(N__33533));
    defparam \pid_front.source_pid_1_1_LC_12_18_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_1_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_1_LC_12_18_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \pid_front.source_pid_1_1_LC_12_18_2  (
            .in0(N__33680),
            .in1(N__32067),
            .in2(N__36196),
            .in3(N__32222),
            .lcout(front_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51322),
            .ce(),
            .sr(N__33533));
    defparam \pid_front.source_pid_1_2_LC_12_18_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_2_LC_12_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_2_LC_12_18_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_front.source_pid_1_2_LC_12_18_3  (
            .in0(N__32068),
            .in1(N__33681),
            .in2(N__39250),
            .in3(N__36401),
            .lcout(front_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51322),
            .ce(),
            .sr(N__33533));
    defparam \pid_front.source_pid_1_3_LC_12_18_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_3_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_3_LC_12_18_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \pid_front.source_pid_1_3_LC_12_18_4  (
            .in0(N__38900),
            .in1(N__32069),
            .in2(N__33686),
            .in3(N__36147),
            .lcout(front_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51322),
            .ce(),
            .sr(N__33533));
    defparam \pid_front.pid_prereg_RNI9EOL_10_LC_12_18_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNI9EOL_10_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNI9EOL_10_LC_12_18_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pid_front.pid_prereg_RNI9EOL_10_LC_12_18_6  (
            .in0(N__33401),
            .in1(N__34891),
            .in2(_gnd_net_),
            .in3(N__33730),
            .lcout(\pid_front.N_532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIH2151_21_LC_12_19_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIH2151_21_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIH2151_21_LC_12_19_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIH2151_21_LC_12_19_0  (
            .in0(N__34854),
            .in1(N__48537),
            .in2(_gnd_net_),
            .in3(N__33412),
            .lcout(\pid_front.N_533 ),
            .ltout(\pid_front.N_533_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIC5I03_4_LC_12_19_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIC5I03_4_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIC5I03_4_LC_12_19_1 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \pid_front.pid_prereg_RNIC5I03_4_LC_12_19_1  (
            .in0(N__38937),
            .in1(N__33572),
            .in2(N__32072),
            .in3(N__38973),
            .lcout(\pid_front.N_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIE0SA_1_LC_12_19_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIE0SA_1_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIE0SA_1_LC_12_19_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \pid_front.pid_prereg_RNIE0SA_1_LC_12_19_2  (
            .in0(N__34853),
            .in1(N__38936),
            .in2(_gnd_net_),
            .in3(N__32221),
            .lcout(),
            .ltout(\pid_front.un1_reset_i_a5_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNISBN11_2_LC_12_19_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNISBN11_2_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNISBN11_2_LC_12_19_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_front.pid_prereg_RNISBN11_2_LC_12_19_3  (
            .in0(N__32228),
            .in1(N__33678),
            .in2(N__32231),
            .in3(N__36397),
            .lcout(\pid_front.un1_reset_i_a5_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_RNIJ92F_0_LC_12_19_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIJ92F_0_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIJ92F_0_LC_12_19_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_esr_RNIJ92F_0_LC_12_19_4  (
            .in0(N__38899),
            .in1(N__36454),
            .in2(N__38975),
            .in3(N__36236),
            .lcout(\pid_front.un1_reset_i_a5_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNI75JF_1_LC_12_20_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNI75JF_1_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNI75JF_1_LC_12_20_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_RNI75JF_1_LC_12_20_1  (
            .in0(N__36452),
            .in1(N__36396),
            .in2(N__33685),
            .in3(N__32217),
            .lcout(\pid_front.un1_reset_i_a5_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIQBDL1_12_LC_12_20_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIQBDL1_12_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIQBDL1_12_LC_12_20_5 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \pid_front.pid_prereg_RNIQBDL1_12_LC_12_20_5  (
            .in0(N__36453),
            .in1(N__34642),
            .in2(N__48536),
            .in3(N__34847),
            .lcout(\pid_front.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_21_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_21_5 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36789),
            .lcout(drone_H_disp_front_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51309),
            .ce(N__42519),
            .sr(N__49601));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_23_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_23_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42601),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51306),
            .ce(N__48344),
            .sr(N__49611));
    defparam \uart_pc.state_RNO_0_2_LC_13_7_1 .C_ON=1'b0;
    defparam \uart_pc.state_RNO_0_2_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_pc.state_RNO_0_2_LC_13_7_1 .LUT_INIT=16'b0000000001110010;
    LogicCell40 \uart_pc.state_RNO_0_2_LC_13_7_1  (
            .in0(N__32130),
            .in1(N__40700),
            .in2(N__32179),
            .in3(N__49774),
            .lcout(\uart_pc.state_srsts_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.state_1_LC_13_7_4 .C_ON=1'b0;
    defparam \uart_pc.state_1_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \uart_pc.state_1_LC_13_7_4 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \uart_pc.state_1_LC_13_7_4  (
            .in0(N__49775),
            .in1(N__32150),
            .in2(N__40711),
            .in3(N__32131),
            .lcout(\uart_pc.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51468),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_13_8_0 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNI5A9J_1_LC_13_8_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uart_drone.timer_Count_RNI5A9J_1_LC_13_8_0  (
            .in0(N__32384),
            .in1(N__32116),
            .in2(N__32387),
            .in3(_gnd_net_),
            .lcout(\uart_drone.un1_state_2_0_a3_0 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\uart_drone.un4_timer_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_2_LC_13_8_1 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_2_LC_13_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_2_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__32465),
            .in2(_gnd_net_),
            .in3(N__32441),
            .lcout(\uart_drone.timer_Count_RNO_0_0_2 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_1 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_3_LC_13_8_2 .C_ON=1'b1;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_3_LC_13_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_drone.timer_Count_RNO_0_3_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__33022),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(\uart_drone.timer_Count_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_drone.un4_timer_Count_1_cry_2 ),
            .carryout(\uart_drone.un4_timer_Count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_RNO_0_4_LC_13_8_3 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.timer_Count_RNO_0_4_LC_13_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uart_drone.timer_Count_RNO_0_4_LC_13_8_3  (
            .in0(N__33077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32426),
            .lcout(\uart_drone.timer_Count_RNO_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.timer_Count_0_LC_13_8_6 .C_ON=1'b0;
    defparam \uart_drone.timer_Count_0_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \uart_drone.timer_Count_0_LC_13_8_6 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \uart_drone.timer_Count_0_LC_13_8_6  (
            .in0(N__48957),
            .in1(N__32416),
            .in2(N__32340),
            .in3(N__32386),
            .lcout(\uart_drone.timer_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51453),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIAT1D1_4_LC_13_8_7 .C_ON=1'b0;
    defparam \uart_drone.state_RNIAT1D1_4_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIAT1D1_4_LC_13_8_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uart_drone.state_RNIAT1D1_4_LC_13_8_7  (
            .in0(N__33076),
            .in1(N__48956),
            .in2(N__32363),
            .in3(N__33157),
            .lcout(\uart_drone.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_0_LC_13_10_1 .C_ON=1'b0;
    defparam \pid_front.state_0_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_0_LC_13_10_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_0_LC_13_10_1  (
            .in0(N__42671),
            .in1(N__32834),
            .in2(_gnd_net_),
            .in3(N__33663),
            .lcout(\pid_front.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51423),
            .ce(),
            .sr(N__49528));
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_12_LC_13_10_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_12_LC_13_10_2  (
            .in0(N__32300),
            .in1(N__32285),
            .in2(N__46188),
            .in3(N__34140),
            .lcout(\ppm_encoder_1.rudderZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51423),
            .ce(),
            .sr(N__49528));
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_8_LC_13_10_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_8_LC_13_10_3  (
            .in0(N__32279),
            .in1(N__32273),
            .in2(N__37605),
            .in3(N__46140),
            .lcout(\ppm_encoder_1.rudderZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51423),
            .ce(),
            .sr(N__49528));
    defparam \ppm_encoder_1.rudder_7_LC_13_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_7_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_7_LC_13_10_4 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_7_LC_13_10_4  (
            .in0(N__32255),
            .in1(N__32249),
            .in2(N__46189),
            .in3(N__45954),
            .lcout(\ppm_encoder_1.rudderZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51423),
            .ce(),
            .sr(N__49528));
    defparam \ppm_encoder_1.rudder_11_LC_13_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_11_LC_13_10_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_11_LC_13_10_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_11_LC_13_10_6  (
            .in0(N__32639),
            .in1(N__32624),
            .in2(N__46187),
            .in3(N__35268),
            .lcout(\ppm_encoder_1.rudderZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51423),
            .ce(),
            .sr(N__49528));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_13_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_13_11_1 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_13_11_1  (
            .in0(N__46786),
            .in1(N__49781),
            .in2(N__46666),
            .in3(N__44914),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51409),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_3_LC_13_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_3_LC_13_12_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_3_LC_13_12_0 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.elevator_3_LC_13_12_0  (
            .in0(N__36125),
            .in1(N__36152),
            .in2(N__41971),
            .in3(N__46365),
            .lcout(\ppm_encoder_1.elevatorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51395),
            .ce(),
            .sr(N__49543));
    defparam \pid_front.state_1_LC_13_12_1 .C_ON=1'b0;
    defparam \pid_front.state_1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.state_1_LC_13_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.state_1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42695),
            .lcout(\pid_front.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51395),
            .ce(),
            .sr(N__49543));
    defparam \ppm_encoder_1.throttle_11_LC_13_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_11_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_11_LC_13_12_3 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_11_LC_13_12_3  (
            .in0(N__32617),
            .in1(N__32591),
            .in2(N__46388),
            .in3(N__34001),
            .lcout(\ppm_encoder_1.throttleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51395),
            .ce(),
            .sr(N__49543));
    defparam \ppm_encoder_1.rudder_13_LC_13_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_13_LC_13_12_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.rudder_13_LC_13_12_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.rudder_13_LC_13_12_4  (
            .in0(N__32585),
            .in1(N__32561),
            .in2(N__41691),
            .in3(N__46366),
            .lcout(\ppm_encoder_1.rudderZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51395),
            .ce(),
            .sr(N__49543));
    defparam \ppm_encoder_1.throttle_2_LC_13_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_2_LC_13_12_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_2_LC_13_12_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_2_LC_13_12_7  (
            .in0(N__32552),
            .in1(N__32545),
            .in2(N__46389),
            .in3(N__37737),
            .lcout(\ppm_encoder_1.throttleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51395),
            .ce(),
            .sr(N__49543));
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_13_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.ppm_output_reg_LC_13_13_0 .LUT_INIT=16'b1110010011110100;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_LC_13_13_0  (
            .in0(N__42128),
            .in1(N__42233),
            .in2(N__32515),
            .in3(N__42104),
            .lcout(ppm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.throttle_10_LC_13_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_10_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_10_LC_13_13_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_10_LC_13_13_1  (
            .in0(N__32498),
            .in1(N__32491),
            .in2(N__46304),
            .in3(N__35619),
            .lcout(\ppm_encoder_1.throttleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.throttle_12_LC_13_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_12_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_12_LC_13_13_2 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.throttle_12_LC_13_13_2  (
            .in0(N__32765),
            .in1(N__46242),
            .in2(N__34109),
            .in3(N__32759),
            .lcout(\ppm_encoder_1.throttleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.throttle_3_LC_13_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_3_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_3_LC_13_13_3 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_3_LC_13_13_3  (
            .in0(N__32741),
            .in1(N__32734),
            .in2(N__46305),
            .in3(N__42016),
            .lcout(\ppm_encoder_1.throttleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.throttle_5_LC_13_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_5_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_5_LC_13_13_4 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \ppm_encoder_1.throttle_5_LC_13_13_4  (
            .in0(N__32708),
            .in1(N__46243),
            .in2(N__38017),
            .in3(N__32702),
            .lcout(\ppm_encoder_1.throttleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.throttle_6_LC_13_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_6_LC_13_13_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_6_LC_13_13_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_6_LC_13_13_5  (
            .in0(N__32678),
            .in1(N__32671),
            .in2(N__46306),
            .in3(N__38802),
            .lcout(\ppm_encoder_1.throttleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51381),
            .ce(),
            .sr(N__49548));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_13_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_13_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_13_14_0  (
            .in0(N__43766),
            .in1(N__40895),
            .in2(_gnd_net_),
            .in3(N__34142),
            .lcout(),
            .ltout(\ppm_encoder_1.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_13_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_13_14_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_13_14_1  (
            .in0(N__43880),
            .in1(_gnd_net_),
            .in2(N__32645),
            .in3(N__41207),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_13_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_13_14_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_13_14_2  (
            .in0(N__46766),
            .in1(N__39214),
            .in2(_gnd_net_),
            .in3(N__37741),
            .lcout(),
            .ltout(\ppm_encoder_1.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_14_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__46631),
            .in2(N__32642),
            .in3(N__37718),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_14_4  (
            .in0(N__46765),
            .in1(N__41970),
            .in2(_gnd_net_),
            .in3(N__42015),
            .lcout(\ppm_encoder_1.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_14_6 .C_ON=1'b0;
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \pid_alt.error_i_acumm_esr_13_LC_13_14_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_alt.error_i_acumm_esr_13_LC_13_14_6  (
            .in0(N__33386),
            .in1(N__33347),
            .in2(_gnd_net_),
            .in3(N__33320),
            .lcout(\pid_alt.error_i_acummZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51368),
            .ce(N__33263),
            .sr(N__33226));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_13_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_13_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_13_14_7  (
            .in0(N__38558),
            .in1(N__33110),
            .in2(_gnd_net_),
            .in3(N__46632),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNIOU0N_4_LC_13_15_0 .C_ON=1'b0;
    defparam \uart_drone.state_RNIOU0N_4_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNIOU0N_4_LC_13_15_0 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uart_drone.state_RNIOU0N_4_LC_13_15_0  (
            .in0(N__32895),
            .in1(N__33173),
            .in2(_gnd_net_),
            .in3(N__49765),
            .lcout(\uart_drone.state_RNIOU0NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.state_RNI26LH_1_LC_13_15_1 .C_ON=1'b0;
    defparam \pid_front.state_RNI26LH_1_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNI26LH_1_LC_13_15_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_front.state_RNI26LH_1_LC_13_15_1  (
            .in0(N__42694),
            .in1(N__32832),
            .in2(_gnd_net_),
            .in3(N__33657),
            .lcout(\pid_front.state_ns_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_13_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_13_15_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_13_15_2  (
            .in0(N__38016),
            .in1(N__46767),
            .in2(_gnd_net_),
            .in3(N__39098),
            .lcout(\ppm_encoder_1.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_RNO_0_3_LC_13_15_3 .C_ON=1'b0;
    defparam \uart_drone.state_RNO_0_3_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_drone.state_RNO_0_3_LC_13_15_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \uart_drone.state_RNO_0_3_LC_13_15_3  (
            .in0(N__32894),
            .in1(N__33104),
            .in2(N__33035),
            .in3(N__32968),
            .lcout(),
            .ltout(\uart_drone.N_145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.state_3_LC_13_15_4 .C_ON=1'b0;
    defparam \uart_drone.state_3_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_drone.state_3_LC_13_15_4 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \uart_drone.state_3_LC_13_15_4  (
            .in0(N__32969),
            .in1(N__32932),
            .in2(N__32915),
            .in3(N__49026),
            .lcout(\uart_drone.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51356),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIQ7UK_1_LC_13_15_5 .C_ON=1'b0;
    defparam \pid_side.state_RNIQ7UK_1_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIQ7UK_1_LC_13_15_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.state_RNIQ7UK_1_LC_13_15_5  (
            .in0(N__50012),
            .in1(N__32833),
            .in2(_gnd_net_),
            .in3(N__35897),
            .lcout(),
            .ltout(\pid_side.state_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNINK4U_1_LC_13_15_6 .C_ON=1'b0;
    defparam \pid_side.state_RNINK4U_1_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNINK4U_1_LC_13_15_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \pid_side.state_RNINK4U_1_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33473),
            .in3(N__49025),
            .lcout(\pid_side.state_RNINK4UZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.state_RNIL5IF_0_LC_13_15_7 .C_ON=1'b0;
    defparam \pid_side.state_RNIL5IF_0_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNIL5IF_0_LC_13_15_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \pid_side.state_RNIL5IF_0_LC_13_15_7  (
            .in0(N__49766),
            .in1(_gnd_net_),
            .in2(N__50040),
            .in3(_gnd_net_),
            .lcout(\pid_side.state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_13_16_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_Altitude_esr_0_LC_13_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_Altitude_esr_0_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42571),
            .lcout(drone_altitude_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51348),
            .ce(N__33469),
            .sr(N__49574));
    defparam \pid_front.pid_prereg_esr_RNIQ3AH3_21_LC_13_17_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNIQ3AH3_21_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNIQ3AH3_21_LC_13_17_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \pid_front.pid_prereg_esr_RNIQ3AH3_21_LC_13_17_2  (
            .in0(N__33656),
            .in1(N__49024),
            .in2(N__48535),
            .in3(N__33488),
            .lcout(),
            .ltout(\pid_front.un1_reset_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNI2A6A6_2_LC_13_17_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNI2A6A6_2_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNI2A6A6_2_LC_13_17_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \pid_front.pid_prereg_RNI2A6A6_2_LC_13_17_3  (
            .in0(N__34643),
            .in1(N__33425),
            .in2(N__33416),
            .in3(N__33413),
            .lcout(\pid_front.pid_prereg_RNI2A6A6Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIEQ7C_6_LC_13_18_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIEQ7C_6_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIEQ7C_6_LC_13_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_RNIEQ7C_6_LC_13_18_0  (
            .in0(N__34924),
            .in1(N__42640),
            .in2(N__36521),
            .in3(N__36484),
            .lcout(\pid_front.un1_reset_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_6_LC_13_18_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_6_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_6_LC_13_18_1 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \pid_front.source_pid_1_6_LC_13_18_1  (
            .in0(N__36485),
            .in1(N__39171),
            .in2(N__33598),
            .in3(N__33661),
            .lcout(front_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.source_pid_1_7_LC_13_18_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_7_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_7_LC_13_18_2 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_front.source_pid_1_7_LC_13_18_2  (
            .in0(N__36520),
            .in1(N__33593),
            .in2(N__45601),
            .in3(N__33664),
            .lcout(front_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.source_pid_1_8_LC_13_18_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_8_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_8_LC_13_18_3 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \pid_front.source_pid_1_8_LC_13_18_3  (
            .in0(N__42641),
            .in1(N__37491),
            .in2(N__33599),
            .in3(N__33662),
            .lcout(front_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.source_pid_1_9_LC_13_18_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_9_LC_13_18_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_9_LC_13_18_4 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \pid_front.source_pid_1_9_LC_13_18_4  (
            .in0(N__34925),
            .in1(N__33597),
            .in2(N__36090),
            .in3(N__33665),
            .lcout(front_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.source_pid_1_10_LC_13_18_5 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_10_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_10_LC_13_18_5 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_front.source_pid_1_10_LC_13_18_5  (
            .in0(N__33588),
            .in1(N__33659),
            .in2(N__38465),
            .in3(N__33731),
            .lcout(front_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.source_pid_1_11_LC_13_18_6 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_11_LC_13_18_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_11_LC_13_18_6 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_front.source_pid_1_11_LC_13_18_6  (
            .in0(N__33660),
            .in1(N__33589),
            .in2(N__36333),
            .in3(N__34892),
            .lcout(front_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51332),
            .ce(),
            .sr(N__33519));
    defparam \pid_front.state_RNIVITE6_1_LC_13_18_7 .C_ON=1'b0;
    defparam \pid_front.state_RNIVITE6_1_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVITE6_1_LC_13_18_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIVITE6_1_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__33658),
            .in2(_gnd_net_),
            .in3(N__33510),
            .lcout(\pid_front.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.source_pid_1_esr_5_LC_13_19_1 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_5_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_5_LC_13_19_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_front.source_pid_1_esr_5_LC_13_19_1  (
            .in0(N__33574),
            .in1(N__33553),
            .in2(_gnd_net_),
            .in3(N__38938),
            .lcout(front_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51324),
            .ce(N__33542),
            .sr(N__33526));
    defparam \pid_front.source_pid_1_esr_4_LC_13_19_2 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_4_LC_13_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_4_LC_13_19_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \pid_front.source_pid_1_esr_4_LC_13_19_2  (
            .in0(N__38939),
            .in1(N__33573),
            .in2(N__33554),
            .in3(N__38974),
            .lcout(front_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51324),
            .ce(N__33542),
            .sr(N__33526));
    defparam \pid_front.source_pid_1_esr_12_LC_13_19_3 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_12_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_12_LC_13_19_3 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \pid_front.source_pid_1_esr_12_LC_13_19_3  (
            .in0(N__34855),
            .in1(N__36455),
            .in2(N__48542),
            .in3(N__34640),
            .lcout(front_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51324),
            .ce(N__33542),
            .sr(N__33526));
    defparam \pid_front.source_pid_1_esr_13_LC_13_19_4 .C_ON=1'b0;
    defparam \pid_front.source_pid_1_esr_13_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.source_pid_1_esr_13_LC_13_19_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \pid_front.source_pid_1_esr_13_LC_13_19_4  (
            .in0(N__34641),
            .in1(N__34856),
            .in2(_gnd_net_),
            .in3(N__48538),
            .lcout(front_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51324),
            .ce(N__33542),
            .sr(N__33526));
    defparam \pid_front.pid_prereg_RNI86SO2_1_LC_13_20_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNI86SO2_1_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNI86SO2_1_LC_13_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_front.pid_prereg_RNI86SO2_1_LC_13_20_3  (
            .in0(N__36206),
            .in1(N__33494),
            .in2(N__33743),
            .in3(N__34633),
            .lcout(\pid_front.N_315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_1_LC_13_21_2 .C_ON=1'b0;
    defparam \pid_front.error_axb_1_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_1_LC_13_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_axb_1_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33479),
            .lcout(\pid_front.error_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIO5UD_6_LC_13_22_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIO5UD_6_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIO5UD_6_LC_13_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_RNIO5UD_6_LC_13_22_5  (
            .in0(N__36478),
            .in1(N__42639),
            .in2(N__34917),
            .in3(N__33717),
            .lcout(),
            .ltout(\pid_front.un1_reset_i_a5_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNIPQGQ_7_LC_13_22_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNIPQGQ_7_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNIPQGQ_7_LC_13_22_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_RNIPQGQ_7_LC_13_22_6  (
            .in0(N__34821),
            .in1(N__34877),
            .in2(N__33746),
            .in3(N__36510),
            .lcout(\pid_front.un1_reset_i_a5_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_10_LC_13_23_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_10_LC_13_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_10_LC_13_23_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_front.pid_prereg_10_LC_13_23_7  (
            .in0(N__48266),
            .in1(N__50459),
            .in2(N__42771),
            .in3(N__33723),
            .lcout(\pid_front.pid_preregZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51307),
            .ce(),
            .sr(N__49613));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_24_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33701),
            .lcout(drone_H_disp_front_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNISRMR1_10_LC_14_6_1 .C_ON=1'b0;
    defparam \reset_module_System.count_RNISRMR1_10_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNISRMR1_10_LC_14_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNISRMR1_10_LC_14_6_1  (
            .in0(N__33863),
            .in1(N__33887),
            .in2(N__33839),
            .in3(N__33764),
            .lcout(\reset_module_System.reset6_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI9O1P_2_LC_14_6_2 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI9O1P_2_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI9O1P_2_LC_14_6_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \reset_module_System.count_RNI9O1P_2_LC_14_6_2  (
            .in0(N__33788),
            .in1(N__33809),
            .in2(N__33959),
            .in3(N__35240),
            .lcout(\reset_module_System.reset6_15 ),
            .ltout(\reset_module_System.reset6_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_LC_14_6_3 .C_ON=1'b0;
    defparam \reset_module_System.count_1_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_1_LC_14_6_3 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \reset_module_System.count_1_LC_14_6_3  (
            .in0(N__33692),
            .in1(N__35211),
            .in2(N__33695),
            .in3(N__35018),
            .lcout(\reset_module_System.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51491),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_1_LC_14_6_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNO_0_1_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_1_LC_14_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \reset_module_System.count_RNO_0_1_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__35055),
            .in2(_gnd_net_),
            .in3(N__35126),
            .lcout(\reset_module_System.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_1_cry_1_c_LC_14_7_0 .C_ON=1'b1;
    defparam \reset_module_System.count_1_cry_1_c_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_1_cry_1_c_LC_14_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \reset_module_System.count_1_cry_1_c_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__35125),
            .in2(N__35057),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\reset_module_System.count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNO_0_2_LC_14_7_1 .C_ON=1'b1;
    defparam \reset_module_System.count_RNO_0_2_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNO_0_2_LC_14_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_RNO_0_2_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__35239),
            .in2(_gnd_net_),
            .in3(N__33812),
            .lcout(\reset_module_System.count_1_2 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_1 ),
            .carryout(\reset_module_System.count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_3_LC_14_7_2 .C_ON=1'b1;
    defparam \reset_module_System.count_3_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_3_LC_14_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_3_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__33808),
            .in2(_gnd_net_),
            .in3(N__33797),
            .lcout(\reset_module_System.countZ0Z_3 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_2 ),
            .carryout(\reset_module_System.count_1_cry_3 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_4_LC_14_7_3 .C_ON=1'b1;
    defparam \reset_module_System.count_4_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_4_LC_14_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_4_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__35138),
            .in2(_gnd_net_),
            .in3(N__33794),
            .lcout(\reset_module_System.countZ0Z_4 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_3 ),
            .carryout(\reset_module_System.count_1_cry_4 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_5_LC_14_7_4 .C_ON=1'b1;
    defparam \reset_module_System.count_5_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_5_LC_14_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_5_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__35150),
            .in2(_gnd_net_),
            .in3(N__33791),
            .lcout(\reset_module_System.countZ0Z_5 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_4 ),
            .carryout(\reset_module_System.count_1_cry_5 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_6_LC_14_7_5 .C_ON=1'b1;
    defparam \reset_module_System.count_6_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_6_LC_14_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_6_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__33787),
            .in2(_gnd_net_),
            .in3(N__33776),
            .lcout(\reset_module_System.countZ0Z_6 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_5 ),
            .carryout(\reset_module_System.count_1_cry_6 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_7_LC_14_7_6 .C_ON=1'b1;
    defparam \reset_module_System.count_7_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_7_LC_14_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_7_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__35177),
            .in2(_gnd_net_),
            .in3(N__33773),
            .lcout(\reset_module_System.countZ0Z_7 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_6 ),
            .carryout(\reset_module_System.count_1_cry_7 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_8_LC_14_7_7 .C_ON=1'b1;
    defparam \reset_module_System.count_8_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_8_LC_14_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_8_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__35189),
            .in2(_gnd_net_),
            .in3(N__33770),
            .lcout(\reset_module_System.countZ0Z_8 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_7 ),
            .carryout(\reset_module_System.count_1_cry_8 ),
            .clk(N__51481),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_9_LC_14_8_0 .C_ON=1'b1;
    defparam \reset_module_System.count_9_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_9_LC_14_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_9_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__35164),
            .in2(_gnd_net_),
            .in3(N__33767),
            .lcout(\reset_module_System.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\reset_module_System.count_1_cry_9 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_10_LC_14_8_1 .C_ON=1'b1;
    defparam \reset_module_System.count_10_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_10_LC_14_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_10_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__33760),
            .in2(_gnd_net_),
            .in3(N__33749),
            .lcout(\reset_module_System.countZ0Z_10 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_9 ),
            .carryout(\reset_module_System.count_1_cry_10 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_11_LC_14_8_2 .C_ON=1'b1;
    defparam \reset_module_System.count_11_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_11_LC_14_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_11_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__33883),
            .in2(_gnd_net_),
            .in3(N__33872),
            .lcout(\reset_module_System.countZ0Z_11 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_10 ),
            .carryout(\reset_module_System.count_1_cry_11 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_12_LC_14_8_3 .C_ON=1'b1;
    defparam \reset_module_System.count_12_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_12_LC_14_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_12_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__35068),
            .in2(_gnd_net_),
            .in3(N__33869),
            .lcout(\reset_module_System.countZ0Z_12 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_11 ),
            .carryout(\reset_module_System.count_1_cry_12 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_13_LC_14_8_4 .C_ON=1'b1;
    defparam \reset_module_System.count_13_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_13_LC_14_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_13_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__33899),
            .in2(_gnd_net_),
            .in3(N__33866),
            .lcout(\reset_module_System.countZ0Z_13 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_12 ),
            .carryout(\reset_module_System.count_1_cry_13 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_14_LC_14_8_5 .C_ON=1'b1;
    defparam \reset_module_System.count_14_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_14_LC_14_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_14_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__33859),
            .in2(_gnd_net_),
            .in3(N__33848),
            .lcout(\reset_module_System.countZ0Z_14 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_13 ),
            .carryout(\reset_module_System.count_1_cry_14 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_15_LC_14_8_6 .C_ON=1'b1;
    defparam \reset_module_System.count_15_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_15_LC_14_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_15_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__33923),
            .in2(_gnd_net_),
            .in3(N__33845),
            .lcout(\reset_module_System.countZ0Z_15 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_14 ),
            .carryout(\reset_module_System.count_1_cry_15 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_16_LC_14_8_7 .C_ON=1'b1;
    defparam \reset_module_System.count_16_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_16_LC_14_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_16_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__35090),
            .in2(_gnd_net_),
            .in3(N__33842),
            .lcout(\reset_module_System.countZ0Z_16 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_15 ),
            .carryout(\reset_module_System.count_1_cry_16 ),
            .clk(N__51469),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_17_LC_14_9_0 .C_ON=1'b1;
    defparam \reset_module_System.count_17_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_17_LC_14_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_17_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__33832),
            .in2(_gnd_net_),
            .in3(N__33821),
            .lcout(\reset_module_System.countZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\reset_module_System.count_1_cry_17 ),
            .clk(N__51454),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_18_LC_14_9_1 .C_ON=1'b1;
    defparam \reset_module_System.count_18_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_18_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_18_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__35104),
            .in2(_gnd_net_),
            .in3(N__33818),
            .lcout(\reset_module_System.countZ0Z_18 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_17 ),
            .carryout(\reset_module_System.count_1_cry_18 ),
            .clk(N__51454),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_19_LC_14_9_2 .C_ON=1'b1;
    defparam \reset_module_System.count_19_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_19_LC_14_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \reset_module_System.count_19_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33935),
            .in3(N__33815),
            .lcout(\reset_module_System.countZ0Z_19 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_18 ),
            .carryout(\reset_module_System.count_1_cry_19 ),
            .clk(N__51454),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_20_LC_14_9_3 .C_ON=1'b1;
    defparam \reset_module_System.count_20_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_20_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \reset_module_System.count_20_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__33955),
            .in2(_gnd_net_),
            .in3(N__33941),
            .lcout(\reset_module_System.countZ0Z_20 ),
            .ltout(),
            .carryin(\reset_module_System.count_1_cry_19 ),
            .carryout(\reset_module_System.count_1_cry_20 ),
            .clk(N__51454),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_21_LC_14_9_4 .C_ON=1'b0;
    defparam \reset_module_System.count_21_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_21_LC_14_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \reset_module_System.count_21_LC_14_9_4  (
            .in0(N__33910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33938),
            .lcout(\reset_module_System.countZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51454),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI34OR1_21_LC_14_9_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI34OR1_21_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI34OR1_21_LC_14_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \reset_module_System.count_RNI34OR1_21_LC_14_9_6  (
            .in0(N__33931),
            .in1(N__33922),
            .in2(N__33911),
            .in3(N__33898),
            .lcout(\reset_module_System.reset6_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_14_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNICBN01_6_LC_14_10_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNICBN01_6_LC_14_10_1  (
            .in0(N__40425),
            .in1(N__45140),
            .in2(_gnd_net_),
            .in3(N__44919),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_7_LC_14_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_7_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_7_LC_14_10_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_7_LC_14_10_2  (
            .in0(N__43375),
            .in1(N__37163),
            .in2(N__43241),
            .in3(N__35405),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51438),
            .ce(),
            .sr(N__49535));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_14_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_14_10_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_14_10_4  (
            .in0(N__44920),
            .in1(_gnd_net_),
            .in2(N__45158),
            .in3(N__40962),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_10_5 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_10_5  (
            .in0(N__40963),
            .in1(N__43871),
            .in2(N__45964),
            .in3(N__43782),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_10_6 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_10_6  (
            .in0(N__43870),
            .in1(N__40426),
            .in2(N__43784),
            .in3(N__38780),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_8_LC_14_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_8_LC_14_10_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_8_LC_14_10_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.init_pulses_8_LC_14_10_7  (
            .in0(N__43223),
            .in1(N__43376),
            .in2(N__35396),
            .in3(N__37148),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51438),
            .ce(),
            .sr(N__49535));
    defparam \ppm_encoder_1.rudder_10_LC_14_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_10_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_10_LC_14_11_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.rudder_10_LC_14_11_0  (
            .in0(N__34049),
            .in1(N__34022),
            .in2(N__41148),
            .in3(N__46311),
            .lcout(\ppm_encoder_1.rudderZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51424),
            .ce(),
            .sr(N__49544));
    defparam \ppm_encoder_1.init_pulses_6_LC_14_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_6_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_6_LC_14_11_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_6_LC_14_11_4  (
            .in0(N__43366),
            .in1(N__37190),
            .in2(N__43238),
            .in3(N__35291),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51424),
            .ce(),
            .sr(N__49544));
    defparam \ppm_encoder_1.elevator_0_LC_14_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_0_LC_14_11_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_0_LC_14_11_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.elevator_0_LC_14_11_7  (
            .in0(N__46310),
            .in1(N__35735),
            .in2(_gnd_net_),
            .in3(N__44003),
            .lcout(\ppm_encoder_1.elevatorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51424),
            .ce(),
            .sr(N__49544));
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_12_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_12_0  (
            .in0(N__33999),
            .in1(N__35269),
            .in2(N__45842),
            .in3(N__45933),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_12_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_12_1  (
            .in0(N__35375),
            .in1(_gnd_net_),
            .in2(N__34010),
            .in3(N__34007),
            .lcout(\ppm_encoder_1.elevator_RNIC22D6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_12_2  (
            .in0(N__33969),
            .in1(N__33981),
            .in2(N__45368),
            .in3(N__45500),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_12_3  (
            .in0(N__46745),
            .in1(N__34000),
            .in2(_gnd_net_),
            .in3(N__33970),
            .lcout(),
            .ltout(\ppm_encoder_1.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_12_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__46589),
            .in2(N__33986),
            .in3(N__33982),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_11_LC_14_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_11_LC_14_12_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_11_LC_14_12_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_11_LC_14_12_5  (
            .in0(N__33983),
            .in1(N__34231),
            .in2(N__46367),
            .in3(N__34364),
            .lcout(\ppm_encoder_1.aileronZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51410),
            .ce(),
            .sr(N__49549));
    defparam \ppm_encoder_1.elevator_11_LC_14_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_11_LC_14_12_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_11_LC_14_12_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_11_LC_14_12_6  (
            .in0(N__33971),
            .in1(N__46321),
            .in2(N__36302),
            .in3(N__36335),
            .lcout(\ppm_encoder_1.elevatorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51410),
            .ce(),
            .sr(N__49549));
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_13_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_13_0  (
            .in0(N__34107),
            .in1(N__34141),
            .in2(N__45935),
            .in3(N__45839),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_14_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIH72D6_12_LC_14_13_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIH72D6_12_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__35422),
            .in2(N__34118),
            .in3(N__34115),
            .lcout(\ppm_encoder_1.elevator_RNIH72D6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_13_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_13_2  (
            .in0(N__34065),
            .in1(N__45477),
            .in2(N__34085),
            .in3(N__45366),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_13_3  (
            .in0(N__34067),
            .in1(N__34108),
            .in2(_gnd_net_),
            .in3(N__46782),
            .lcout(),
            .ltout(\ppm_encoder_1.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_13_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_13_4  (
            .in0(N__46630),
            .in1(_gnd_net_),
            .in2(N__34088),
            .in3(N__34083),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_12_LC_14_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_12_LC_14_13_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_12_LC_14_13_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_12_LC_14_13_5  (
            .in0(N__34084),
            .in1(N__37820),
            .in2(N__46307),
            .in3(N__34352),
            .lcout(\ppm_encoder_1.aileronZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51396),
            .ce(),
            .sr(N__49557));
    defparam \ppm_encoder_1.elevator_12_LC_14_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_12_LC_14_13_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_12_LC_14_13_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_12_LC_14_13_6  (
            .in0(N__34066),
            .in1(N__46244),
            .in2(N__36284),
            .in3(N__36260),
            .lcout(\ppm_encoder_1.elevatorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51396),
            .ce(),
            .sr(N__49557));
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__46026),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_14_14_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_14_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__35977),
            .in2(N__47883),
            .in3(N__34052),
            .lcout(\ppm_encoder_1.un1_aileron_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_0 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_14_14_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_14_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__35929),
            .in2(_gnd_net_),
            .in3(N__34169),
            .lcout(\ppm_encoder_1.un1_aileron_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_1 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_14_14_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_14_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__38615),
            .in2(N__47884),
            .in3(N__34166),
            .lcout(\ppm_encoder_1.un1_aileron_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_2 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_14_14_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_14_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__46868),
            .in2(_gnd_net_),
            .in3(N__34163),
            .lcout(\ppm_encoder_1.un1_aileron_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_3 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_14_14_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__38579),
            .in2(_gnd_net_),
            .in3(N__34160),
            .lcout(\ppm_encoder_1.un1_aileron_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_4 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_14_14_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_14_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__47842),
            .in2(N__38698),
            .in3(N__34157),
            .lcout(\ppm_encoder_1.un1_aileron_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_5 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_14_14_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_14_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__45654),
            .in2(_gnd_net_),
            .in3(N__34154),
            .lcout(\ppm_encoder_1.un1_aileron_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_6 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_14_15_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_14_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__37542),
            .in2(_gnd_net_),
            .in3(N__34151),
            .lcout(\ppm_encoder_1.un1_aileron_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\ppm_encoder_1.un1_aileron_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_14_15_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_14_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__38514),
            .in2(_gnd_net_),
            .in3(N__34148),
            .lcout(\ppm_encoder_1.un1_aileron_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_8 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_14_15_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_14_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__36036),
            .in2(_gnd_net_),
            .in3(N__34145),
            .lcout(\ppm_encoder_1.un1_aileron_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_9 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_14_15_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_14_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__34224),
            .in2(_gnd_net_),
            .in3(N__34355),
            .lcout(\ppm_encoder_1.un1_aileron_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_10 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_14_15_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_14_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__37819),
            .in2(_gnd_net_),
            .in3(N__34343),
            .lcout(\ppm_encoder_1.un1_aileron_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_11 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_14_15_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_14_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__47990),
            .in2(N__41621),
            .in3(N__34340),
            .lcout(\ppm_encoder_1.un1_aileron_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_aileron_cry_12 ),
            .carryout(\ppm_encoder_1.un1_aileron_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_14_LC_14_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_14_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_esr_14_LC_14_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.aileron_esr_14_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34337),
            .lcout(\ppm_encoder_1.aileronZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51369),
            .ce(N__36697),
            .sr(N__49575));
    defparam \pid_alt.error_cry_0_c_inv_LC_14_15_7 .C_ON=1'b0;
    defparam \pid_alt.error_cry_0_c_inv_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \pid_alt.error_cry_0_c_inv_LC_14_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_alt.error_cry_0_c_inv_LC_14_15_7  (
            .in0(N__47989),
            .in1(N__34273),
            .in2(_gnd_net_),
            .in3(N__34296),
            .lcout(\pid_alt.drone_altitude_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_10_LC_14_16_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_10_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_10_LC_14_16_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_side.source_pid_1_10_LC_14_16_0  (
            .in0(N__38170),
            .in1(N__35886),
            .in2(N__36041),
            .in3(N__34259),
            .lcout(side_order_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.source_pid_1_11_LC_14_16_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_11_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_11_LC_14_16_1 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_side.source_pid_1_11_LC_14_16_1  (
            .in0(N__35887),
            .in1(N__38171),
            .in2(N__34232),
            .in3(N__34439),
            .lcout(side_order_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.source_pid_1_6_LC_14_16_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_6_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_6_LC_14_16_2 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_side.source_pid_1_6_LC_14_16_2  (
            .in0(N__38172),
            .in1(N__35888),
            .in2(N__38697),
            .in3(N__34208),
            .lcout(side_order_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.source_pid_1_7_LC_14_16_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_7_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_7_LC_14_16_3 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_side.source_pid_1_7_LC_14_16_3  (
            .in0(N__35889),
            .in1(N__38173),
            .in2(N__45658),
            .in3(N__34406),
            .lcout(side_order_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.source_pid_1_8_LC_14_16_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_8_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_8_LC_14_16_4 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \pid_side.source_pid_1_8_LC_14_16_4  (
            .in0(N__38174),
            .in1(N__35890),
            .in2(N__37552),
            .in3(N__34601),
            .lcout(side_order_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.source_pid_1_9_LC_14_16_5 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_9_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_9_LC_14_16_5 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \pid_side.source_pid_1_9_LC_14_16_5  (
            .in0(N__35891),
            .in1(N__38175),
            .in2(N__38524),
            .in3(N__34568),
            .lcout(side_order_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51357),
            .ce(),
            .sr(N__38073));
    defparam \pid_side.state_RNI34HSI_1_LC_14_16_6 .C_ON=1'b0;
    defparam \pid_side.state_RNI34HSI_1_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.state_RNI34HSI_1_LC_14_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_side.state_RNI34HSI_1_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__35885),
            .in2(_gnd_net_),
            .in3(N__38060),
            .lcout(\pid_side.state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNIOB8E3_2_LC_14_17_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIOB8E3_2_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIOB8E3_2_LC_14_17_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pid_side.pid_prereg_RNIOB8E3_2_LC_14_17_0  (
            .in0(N__34664),
            .in1(N__35896),
            .in2(N__34655),
            .in3(N__35956),
            .lcout(\pid_side.un1_reset_i_a5_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIH97T2_21_LC_14_17_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIH97T2_21_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIH97T2_21_LC_14_17_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIH97T2_21_LC_14_17_2  (
            .in0(N__38361),
            .in1(N__36007),
            .in2(_gnd_net_),
            .in3(N__38302),
            .lcout(\pid_side.N_534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_drone.bit_Count_RNO_0_2_LC_14_17_5 .C_ON=1'b0;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_drone.bit_Count_RNO_0_2_LC_14_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_drone.bit_Count_RNO_0_2_LC_14_17_5  (
            .in0(N__34524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34472),
            .lcout(\uart_drone.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNILTAI1_0_LC_14_17_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNILTAI1_0_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNILTAI1_0_LC_14_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_side.pid_prereg_esr_RNILTAI1_0_LC_14_17_6  (
            .in0(N__38246),
            .in1(N__35783),
            .in2(N__38147),
            .in3(N__41919),
            .lcout(\pid_side.un1_reset_i_a5_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNITODS2_7_LC_14_17_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNITODS2_7_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNITODS2_7_LC_14_17_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \pid_side.pid_prereg_RNITODS2_7_LC_14_17_7  (
            .in0(N__34432),
            .in1(N__34402),
            .in2(N__38314),
            .in3(N__34376),
            .lcout(\pid_side.un1_reset_i_a5_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_0_LC_14_18_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_0_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.pid_prereg_esr_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50072),
            .lcout(\pid_front.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51339),
            .ce(N__48481),
            .sr(N__49598));
    defparam \pid_side.pid_prereg_RNI7QS63_14_LC_14_18_3 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNI7QS63_14_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNI7QS63_14_LC_14_18_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_side.pid_prereg_RNI7QS63_14_LC_14_18_3  (
            .in0(N__34805),
            .in1(N__34789),
            .in2(N__34772),
            .in3(N__34757),
            .lcout(\pid_side.N_563 ),
            .ltout(\pid_side.N_563_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNIGPS29_1_LC_14_18_4 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIGPS29_1_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIGPS29_1_LC_14_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \pid_side.pid_prereg_RNIGPS29_1_LC_14_18_4  (
            .in0(N__34739),
            .in1(N__34721),
            .in2(N__34733),
            .in3(N__34730),
            .lcout(),
            .ltout(\pid_side.N_311_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNIQG8J9_21_LC_14_18_5 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIQG8J9_21_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIQG8J9_21_LC_14_18_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIQG8J9_21_LC_14_18_5  (
            .in0(N__38360),
            .in1(N__35878),
            .in2(N__34724),
            .in3(N__49023),
            .lcout(\pid_side.un1_reset_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNIN87D1_1_LC_14_19_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNIN87D1_1_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNIN87D1_1_LC_14_19_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_side.pid_prereg_RNIN87D1_1_LC_14_19_0  (
            .in0(N__37842),
            .in1(N__35948),
            .in2(N__35877),
            .in3(N__49831),
            .lcout(\pid_side.un1_reset_i_a5_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_2_LC_14_19_2 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_2_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_2_LC_14_19_2 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_side.pid_prereg_2_LC_14_19_2  (
            .in0(N__50019),
            .in1(N__34715),
            .in2(N__34682),
            .in3(N__35949),
            .lcout(\pid_side.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51333),
            .ce(),
            .sr(N__49602));
    defparam \pid_side.pid_prereg_RNI2JR61_1_LC_14_19_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNI2JR61_1_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNI2JR61_1_LC_14_19_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \pid_side.pid_prereg_RNI2JR61_1_LC_14_19_6  (
            .in0(N__38138),
            .in1(N__38315),
            .in2(_gnd_net_),
            .in3(N__49830),
            .lcout(\pid_side.un1_reset_i_a5_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_RNI39UK1_0_LC_14_19_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNI39UK1_0_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNI39UK1_0_LC_14_19_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_side.pid_prereg_esr_RNI39UK1_0_LC_14_19_7  (
            .in0(N__35788),
            .in1(N__41920),
            .in2(N__38258),
            .in3(N__37843),
            .lcout(\pid_side.un1_reset_i_a5_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_RNI3CC11_14_LC_14_20_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNI3CC11_14_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNI3CC11_14_LC_14_20_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \pid_front.pid_prereg_RNI3CC11_14_LC_14_20_0  (
            .in0(N__36356),
            .in1(N__34609),
            .in2(N__34961),
            .in3(N__36416),
            .lcout(\pid_front.N_569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_14_LC_14_20_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_14_LC_14_20_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_14_LC_14_20_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_front.pid_prereg_14_LC_14_20_6  (
            .in0(N__50543),
            .in1(N__47768),
            .in2(N__42817),
            .in3(N__34610),
            .lcout(\pid_front.pid_preregZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51325),
            .ce(),
            .sr(N__49606));
    defparam \pid_front.pid_prereg_RNID03J_17_LC_14_21_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_RNID03J_17_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_RNID03J_17_LC_14_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_RNID03J_17_LC_14_21_3  (
            .in0(N__34951),
            .in1(N__36532),
            .in2(N__34940),
            .in3(N__36544),
            .lcout(\pid_front.m7_e_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_9_LC_14_22_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_9_LC_14_22_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_9_LC_14_22_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.elevator_9_LC_14_22_1  (
            .in0(N__36092),
            .in1(N__36062),
            .in2(N__46397),
            .in3(N__35695),
            .lcout(\ppm_encoder_1.elevatorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(N__49614));
    defparam \pid_front.pid_prereg_18_LC_14_22_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_18_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_18_LC_14_22_3 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_18_LC_14_22_3  (
            .in0(N__42800),
            .in1(N__48590),
            .in2(N__50264),
            .in3(N__34952),
            .lcout(\pid_front.pid_preregZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(N__49614));
    defparam \pid_front.pid_prereg_19_LC_14_22_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_19_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_19_LC_14_22_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_19_LC_14_22_5  (
            .in0(N__42801),
            .in1(N__48575),
            .in2(N__51911),
            .in3(N__34939),
            .lcout(\pid_front.pid_preregZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51315),
            .ce(),
            .sr(N__49614));
    defparam \pid_front.pid_prereg_9_LC_14_23_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_9_LC_14_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_9_LC_14_23_3 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pid_front.pid_prereg_9_LC_14_23_3  (
            .in0(N__47591),
            .in1(N__48743),
            .in2(N__34923),
            .in3(N__42776),
            .lcout(\pid_front.pid_preregZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51312),
            .ce(),
            .sr(N__49617));
    defparam \pid_front.pid_prereg_11_LC_14_23_6 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_11_LC_14_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_11_LC_14_23_6 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_front.pid_prereg_11_LC_14_23_6  (
            .in0(N__51797),
            .in1(N__48251),
            .in2(N__42805),
            .in3(N__34884),
            .lcout(\pid_front.pid_preregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51312),
            .ce(),
            .sr(N__49617));
    defparam \pid_front.pid_prereg_13_LC_14_23_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_13_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_13_LC_14_23_7 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pid_front.pid_prereg_13_LC_14_23_7  (
            .in0(N__51863),
            .in1(N__47783),
            .in2(N__34841),
            .in3(N__42775),
            .lcout(\pid_front.pid_preregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51312),
            .ce(),
            .sr(N__49617));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_14_24_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_14_24_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_14_24_4  (
            .in0(N__36620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(drone_H_disp_front_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51308),
            .ce(N__48354),
            .sr(N__49620));
    defparam \reset_module_System.reset_LC_15_6_0 .C_ON=1'b0;
    defparam \reset_module_System.reset_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.reset_LC_15_6_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \reset_module_System.reset_LC_15_6_0  (
            .in0(N__35223),
            .in1(N__35207),
            .in2(_gnd_net_),
            .in3(N__35015),
            .lcout(reset_system),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51502),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_2_LC_15_6_4 .C_ON=1'b0;
    defparam \reset_module_System.count_2_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_2_LC_15_6_4 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \reset_module_System.count_2_LC_15_6_4  (
            .in0(N__35212),
            .in1(N__35246),
            .in2(N__35228),
            .in3(N__35017),
            .lcout(\reset_module_System.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51502),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_0_LC_15_6_5 .C_ON=1'b0;
    defparam \reset_module_System.count_0_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \reset_module_System.count_0_LC_15_6_5 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \reset_module_System.count_0_LC_15_6_5  (
            .in0(N__35016),
            .in1(N__35224),
            .in2(N__35213),
            .in3(N__35056),
            .lcout(\reset_module_System.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51502),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_3 .C_ON=1'b0;
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNI97FD_5_LC_15_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \reset_module_System.count_RNI97FD_5_LC_15_7_3  (
            .in0(N__35188),
            .in1(N__35176),
            .in2(N__35165),
            .in3(N__35149),
            .lcout(\reset_module_System.reset6_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIR9N6_1_LC_15_7_4 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIR9N6_1_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIR9N6_1_LC_15_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \reset_module_System.count_RNIR9N6_1_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__35137),
            .in2(_gnd_net_),
            .in3(N__35124),
            .lcout(),
            .ltout(\reset_module_System.reset6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_5 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIA72I1_16_LC_15_7_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \reset_module_System.count_RNIA72I1_16_LC_15_7_5  (
            .in0(N__35108),
            .in1(N__35089),
            .in2(N__35078),
            .in3(N__35075),
            .lcout(),
            .ltout(\reset_module_System.reset6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_7_6 .C_ON=1'b0;
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \reset_module_System.count_RNIMJ304_12_LC_15_7_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \reset_module_System.count_RNIMJ304_12_LC_15_7_6  (
            .in0(N__35069),
            .in1(N__35054),
            .in2(N__35030),
            .in3(N__35027),
            .lcout(\reset_module_System.reset6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_9_LC_15_8_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_9_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_9_LC_15_8_7 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.rudder_9_LC_15_8_7  (
            .in0(N__35000),
            .in1(N__34985),
            .in2(N__46390),
            .in3(N__35664),
            .lcout(\ppm_encoder_1.rudderZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51482),
            .ce(),
            .sr(N__49529));
    defparam \ppm_encoder_1.init_pulses_11_LC_15_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_11_LC_15_9_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_11_LC_15_9_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_11_LC_15_9_0  (
            .in0(N__43353),
            .in1(N__43237),
            .in2(N__37286),
            .in3(N__35348),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51470),
            .ce(),
            .sr(N__49536));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_15_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_15_9_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_15_9_1  (
            .in0(N__35283),
            .in1(N__45144),
            .in2(_gnd_net_),
            .in3(N__44931),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_15_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_15_9_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_15_9_2  (
            .in0(N__44932),
            .in1(_gnd_net_),
            .in2(N__45159),
            .in3(N__35284),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_9_3  (
            .in0(N__35285),
            .in1(N__43753),
            .in2(_gnd_net_),
            .in3(N__35273),
            .lcout(),
            .ltout(\ppm_encoder_1.N_313_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_9_4 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__41203),
            .in2(N__35249),
            .in3(N__43869),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_12_LC_15_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_12_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_12_LC_15_9_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_12_LC_15_9_5  (
            .in0(N__43236),
            .in1(N__43354),
            .in2(N__37274),
            .in3(N__35330),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51470),
            .ce(),
            .sr(N__49536));
    defparam \ppm_encoder_1.init_pulses_16_LC_15_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_16_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_16_LC_15_10_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_16_LC_15_10_0  (
            .in0(N__43350),
            .in1(N__37247),
            .in2(N__43242),
            .in3(N__35471),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51455),
            .ce(),
            .sr(N__49545));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_15_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_15_10_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_15_10_1  (
            .in0(N__45180),
            .in1(N__45136),
            .in2(_gnd_net_),
            .in3(N__44917),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_17_LC_15_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_17_LC_15_10_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_17_LC_15_10_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_17_LC_15_10_2  (
            .in0(N__43351),
            .in1(N__37232),
            .in2(N__43243),
            .in3(N__35447),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51455),
            .ce(),
            .sr(N__49545));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_15_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_15_10_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_15_10_3  (
            .in0(N__44244),
            .in1(N__45135),
            .in2(_gnd_net_),
            .in3(N__44916),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_15_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_15_10_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_15_10_4  (
            .in0(N__44918),
            .in1(_gnd_net_),
            .in2(N__45157),
            .in3(N__44245),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_18_LC_15_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_18_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_18_LC_15_10_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_18_LC_15_10_5  (
            .in0(N__43221),
            .in1(N__37220),
            .in2(N__43373),
            .in3(N__35432),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51455),
            .ce(),
            .sr(N__49545));
    defparam \ppm_encoder_1.init_pulses_2_LC_15_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_2_LC_15_10_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_2_LC_15_10_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ppm_encoder_1.init_pulses_2_LC_15_10_6  (
            .in0(N__43352),
            .in1(N__43222),
            .in2(N__37214),
            .in3(N__35309),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51455),
            .ce(),
            .sr(N__49545));
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_15_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI87N01_2_LC_15_10_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI87N01_2_LC_15_10_7  (
            .in0(N__40911),
            .in1(N__45134),
            .in2(_gnd_net_),
            .in3(N__44915),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_11_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNINSH16_0_LC_15_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNINSH16_0_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__42045),
            .in2(N__37655),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_11_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__37921),
            .in2(N__37910),
            .in3(N__35312),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_11_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__37687),
            .in2(N__37673),
            .in3(N__35303),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_11_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__41996),
            .in2(N__41939),
            .in3(N__35300),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_11_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__40789),
            .in2(N__38033),
            .in3(N__35297),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_11_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__44122),
            .in2(N__37982),
            .in3(N__35294),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_11_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__38743),
            .in2(N__38723),
            .in3(N__35408),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_11_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__45727),
            .in2(N__45707),
            .in3(N__35399),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_12_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__44077),
            .in2(N__37571),
            .in3(N__35384),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_8 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_12_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__44146),
            .in2(N__35486),
            .in3(N__35381),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_12_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__35587),
            .in2(N__35573),
            .in3(N__35378),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_12_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__35371),
            .in2(N__35357),
            .in3(N__35339),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_12_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__35336),
            .in2(N__35423),
            .in3(N__35321),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_12_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__41659),
            .in2(N__41645),
            .in3(N__35318),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_12_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__41851),
            .in2(N__41837),
            .in3(N__35315),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_12_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__37409),
            .in2(N__37361),
            .in3(N__35474),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_13_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__44597),
            .in2(_gnd_net_),
            .in3(N__35462),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_16 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_13_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35459),
            .in3(N__35438),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_0_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_13_2  (
            .in0(N__40859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35435),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_13_3  (
            .in0(N__46795),
            .in1(N__37947),
            .in2(_gnd_net_),
            .in3(N__37893),
            .lcout(\ppm_encoder_1.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_13_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_13_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_15_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_10_LC_15_13_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_10_LC_15_13_5  (
            .in0(N__41166),
            .in1(N__45148),
            .in2(_gnd_net_),
            .in3(N__44909),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_15_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_15_13_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_15_13_6  (
            .in0(N__44910),
            .in1(_gnd_net_),
            .in2(N__45160),
            .in3(N__40887),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_15_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_15_13_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_15_13_7  (
            .in0(N__37445),
            .in1(N__45152),
            .in2(_gnd_net_),
            .in3(N__44911),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_15_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_15_14_0 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_15_14_0  (
            .in0(N__43881),
            .in1(N__44105),
            .in2(N__37613),
            .in3(N__43728),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_14_3  (
            .in0(N__46663),
            .in1(N__35546),
            .in2(_gnd_net_),
            .in3(N__37966),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_1_LC_15_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_1_LC_15_14_4 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_1_LC_15_14_4 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.aileron_1_LC_15_14_4  (
            .in0(N__37967),
            .in1(N__35540),
            .in2(N__46308),
            .in3(N__35978),
            .lcout(\ppm_encoder_1.aileronZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51397),
            .ce(),
            .sr(N__49576));
    defparam \ppm_encoder_1.elevator_1_LC_15_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_1_LC_15_14_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_1_LC_15_14_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \ppm_encoder_1.elevator_1_LC_15_14_5  (
            .in0(N__36167),
            .in1(N__36197),
            .in2(N__37952),
            .in3(N__46255),
            .lcout(\ppm_encoder_1.elevatorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51397),
            .ce(),
            .sr(N__49576));
    defparam \ppm_encoder_1.throttle_1_LC_15_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_1_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_1_LC_15_14_6 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.throttle_1_LC_15_14_6  (
            .in0(N__35534),
            .in1(N__35522),
            .in2(N__46309),
            .in3(N__37894),
            .lcout(\ppm_encoder_1.throttleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51397),
            .ce(),
            .sr(N__49576));
    defparam \ppm_encoder_1.aileron_2_LC_15_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_2_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_2_LC_15_14_7 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_2_LC_15_14_7  (
            .in0(N__37714),
            .in1(N__46248),
            .in2(N__35930),
            .in3(N__35495),
            .lcout(\ppm_encoder_1.aileronZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51397),
            .ce(),
            .sr(N__49576));
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_15_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIGN7O2_9_LC_15_15_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNIGN7O2_9_LC_15_15_0  (
            .in0(N__35701),
            .in1(N__38485),
            .in2(N__45498),
            .in3(N__45367),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_15_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIV9PO6_9_LC_15_15_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIV9PO6_9_LC_15_15_1  (
            .in0(N__44150),
            .in1(_gnd_net_),
            .in2(N__35489),
            .in3(N__35627),
            .lcout(\ppm_encoder_1.throttle_RNIV9PO6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_15_2  (
            .in0(N__46665),
            .in1(N__35681),
            .in2(_gnd_net_),
            .in3(N__38486),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_15_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_15_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_15_15_3  (
            .in0(N__35648),
            .in1(N__46807),
            .in2(_gnd_net_),
            .in3(N__35702),
            .lcout(\ppm_encoder_1.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_15_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_15_15_4 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_15_15_4  (
            .in0(N__35666),
            .in1(N__43711),
            .in2(N__43886),
            .in3(N__44177),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_9_LC_15_15_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_9_LC_15_15_5  (
            .in0(N__44498),
            .in1(_gnd_net_),
            .in2(N__35675),
            .in3(N__35672),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51382),
            .ce(N__44410),
            .sr(N__49584));
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_15_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNI04QV2_9_LC_15_15_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNI04QV2_9_LC_15_15_6  (
            .in0(N__35665),
            .in1(N__35647),
            .in2(N__45832),
            .in3(N__45897),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_15_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_15_15_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_15_15_7  (
            .in0(N__43710),
            .in1(N__43882),
            .in2(_gnd_net_),
            .in3(N__41416),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_15_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGUOT2_10_LC_15_16_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIGUOT2_10_LC_15_16_1  (
            .in0(N__35620),
            .in1(N__41149),
            .in2(N__45841),
            .in3(N__45905),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_15_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI7T1D6_10_LC_15_16_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNI7T1D6_10_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__35594),
            .in2(N__35576),
            .in3(N__35561),
            .lcout(\ppm_encoder_1.elevator_RNI7T1D6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_15_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI02LH2_10_LC_15_16_3 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNI02LH2_10_LC_15_16_3  (
            .in0(N__38424),
            .in1(N__36018),
            .in2(N__45494),
            .in3(N__45353),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_16_5  (
            .in0(N__46664),
            .in1(N__35555),
            .in2(_gnd_net_),
            .in3(N__36019),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_10_LC_15_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_10_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_10_LC_15_16_6 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.aileron_10_LC_15_16_6  (
            .in0(N__36020),
            .in1(N__46256),
            .in2(N__36050),
            .in3(N__36037),
            .lcout(\ppm_encoder_1.aileronZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51370),
            .ce(),
            .sr(N__49593));
    defparam \pid_side.pid_prereg_esr_RNIAA5MI_21_LC_15_17_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIAA5MI_21_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIAA5MI_21_LC_15_17_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \pid_side.pid_prereg_esr_RNIAA5MI_21_LC_15_17_0  (
            .in0(N__38389),
            .in1(N__36008),
            .in2(N__35993),
            .in3(N__35984),
            .lcout(\pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_0_LC_15_17_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_0_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_0_LC_15_17_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_side.source_pid_1_0_LC_15_17_1  (
            .in0(N__35747),
            .in1(N__35892),
            .in2(N__46030),
            .in3(N__41921),
            .lcout(side_order_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51358),
            .ce(),
            .sr(N__38075));
    defparam \pid_side.source_pid_1_1_LC_15_17_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_1_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_1_LC_15_17_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \pid_side.source_pid_1_1_LC_15_17_2  (
            .in0(N__35893),
            .in1(N__35748),
            .in2(N__49835),
            .in3(N__35976),
            .lcout(side_order_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51358),
            .ce(),
            .sr(N__38075));
    defparam \pid_side.source_pid_1_2_LC_15_17_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_2_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_2_LC_15_17_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \pid_side.source_pid_1_2_LC_15_17_3  (
            .in0(N__35749),
            .in1(N__35894),
            .in2(N__35928),
            .in3(N__35957),
            .lcout(side_order_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51358),
            .ce(),
            .sr(N__38075));
    defparam \pid_side.source_pid_1_3_LC_15_17_4 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_3_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_3_LC_15_17_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \pid_side.source_pid_1_3_LC_15_17_4  (
            .in0(N__35895),
            .in1(N__35750),
            .in2(N__35792),
            .in3(N__38614),
            .lcout(side_order_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51358),
            .ce(),
            .sr(N__38075));
    defparam \pid_side.pid_prereg_esr_RNIIK254_21_LC_15_17_6 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_RNIIK254_21_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_esr_RNIIK254_21_LC_15_17_6 .LUT_INIT=16'b0000110100000101;
    LogicCell40 \pid_side.pid_prereg_esr_RNIIK254_21_LC_15_17_6  (
            .in0(N__38388),
            .in1(N__38316),
            .in2(N__38370),
            .in3(N__37855),
            .lcout(\pid_side.N_291 ),
            .ltout(\pid_side.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_RNISEFQ7_4_LC_15_17_7 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_RNISEFQ7_4_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \pid_side.pid_prereg_RNISEFQ7_4_LC_15_17_7 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \pid_side.pid_prereg_RNISEFQ7_4_LC_15_17_7  (
            .in0(N__38256),
            .in1(N__38123),
            .in2(N__35753),
            .in3(N__38191),
            .lcout(\pid_side.N_451_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_15_18_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__35727),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_15_18_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_15_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__36192),
            .in2(N__48084),
            .in3(N__36158),
            .lcout(\ppm_encoder_1.un1_elevator_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_0 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_15_18_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_15_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__39246),
            .in2(_gnd_net_),
            .in3(N__36155),
            .lcout(\ppm_encoder_1.un1_elevator_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_1 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_15_18_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_15_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__36148),
            .in2(N__48085),
            .in3(N__36110),
            .lcout(\ppm_encoder_1.un1_elevator_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_2 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_15_18_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__46831),
            .in2(_gnd_net_),
            .in3(N__36107),
            .lcout(\ppm_encoder_1.un1_elevator_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_3 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_15_18_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_15_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__39127),
            .in2(_gnd_net_),
            .in3(N__36104),
            .lcout(\ppm_encoder_1.un1_elevator_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_4 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_15_18_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_15_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__39172),
            .in2(N__48086),
            .in3(N__36101),
            .lcout(\ppm_encoder_1.un1_elevator_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_5 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_15_18_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_15_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__45597),
            .in2(_gnd_net_),
            .in3(N__36098),
            .lcout(\ppm_encoder_1.un1_elevator_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_6 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_15_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_15_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__37498),
            .in2(_gnd_net_),
            .in3(N__36095),
            .lcout(\ppm_encoder_1.un1_elevator_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\ppm_encoder_1.un1_elevator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_15_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_15_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__36091),
            .in2(_gnd_net_),
            .in3(N__36341),
            .lcout(\ppm_encoder_1.un1_elevator_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_8 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_15_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_15_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__38464),
            .in2(_gnd_net_),
            .in3(N__36338),
            .lcout(\ppm_encoder_1.un1_elevator_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_9 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_15_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_15_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__36334),
            .in2(_gnd_net_),
            .in3(N__36287),
            .lcout(\ppm_encoder_1.un1_elevator_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_10 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_15_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_15_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__36277),
            .in2(_gnd_net_),
            .in3(N__36245),
            .lcout(\ppm_encoder_1.un1_elevator_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_11 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_15_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_15_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__41560),
            .in2(N__48087),
            .in3(N__36242),
            .lcout(\ppm_encoder_1.un1_elevator_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_elevator_cry_12 ),
            .carryout(\ppm_encoder_1.un1_elevator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_esr_14_LC_15_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_esr_14_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_esr_14_LC_15_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.elevator_esr_14_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36239),
            .lcout(\ppm_encoder_1.elevatorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51340),
            .ce(N__36692),
            .sr(N__49607));
    defparam \pid_front.pid_prereg_esr_RNI5QBD_0_LC_15_20_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_RNI5QBD_0_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.pid_prereg_esr_RNI5QBD_0_LC_15_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \pid_front.pid_prereg_esr_RNI5QBD_0_LC_15_20_7  (
            .in0(N__38955),
            .in1(N__38886),
            .in2(N__38925),
            .in3(N__36231),
            .lcout(\pid_front.un1_reset_i_a5_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_15_21_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_15_21_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_15_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36970),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51326),
            .ce(N__42526),
            .sr(N__49615));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_15_21_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_15_21_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_15_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36880),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51326),
            .ce(N__42526),
            .sr(N__49615));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_15_21_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_15_21_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_15_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48448),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51326),
            .ce(N__42526),
            .sr(N__49615));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_15_21_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_15_21_4 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_15_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36605),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51326),
            .ce(N__42526),
            .sr(N__49615));
    defparam \pid_front.pid_prereg_17_LC_15_22_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_17_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_17_LC_15_22_1 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \pid_front.pid_prereg_17_LC_15_22_1  (
            .in0(N__42791),
            .in1(N__47729),
            .in2(N__36548),
            .in3(N__51569),
            .lcout(\pid_front.pid_preregZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51319),
            .ce(),
            .sr(N__49618));
    defparam \pid_front.pid_prereg_20_LC_15_22_2 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_20_LC_15_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_20_LC_15_22_2 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_20_LC_15_22_2  (
            .in0(N__42798),
            .in1(N__48560),
            .in2(N__51722),
            .in3(N__36533),
            .lcout(\pid_front.pid_preregZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51319),
            .ce(),
            .sr(N__49618));
    defparam \pid_front.pid_prereg_7_LC_15_22_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_7_LC_15_22_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_7_LC_15_22_4 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pid_front.pid_prereg_7_LC_15_22_4  (
            .in0(N__42799),
            .in1(N__50417),
            .in2(N__36516),
            .in3(N__47612),
            .lcout(\pid_front.pid_preregZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51319),
            .ce(),
            .sr(N__49618));
    defparam \pid_front.pid_prereg_6_LC_15_22_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_6_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_6_LC_15_22_5 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_front.pid_prereg_6_LC_15_22_5  (
            .in0(N__47627),
            .in1(N__50312),
            .in2(N__42816),
            .in3(N__36477),
            .lcout(\pid_front.pid_preregZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51319),
            .ce(),
            .sr(N__49618));
    defparam \pid_front.pid_prereg_12_LC_15_22_7 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_12_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_12_LC_15_22_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_front.pid_prereg_12_LC_15_22_7  (
            .in0(N__51767),
            .in1(N__47798),
            .in2(N__42815),
            .in3(N__36440),
            .lcout(\pid_front.pid_preregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51319),
            .ce(),
            .sr(N__49618));
    defparam \pid_front.pid_prereg_16_LC_15_23_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_16_LC_15_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_16_LC_15_23_1 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_front.pid_prereg_16_LC_15_23_1  (
            .in0(N__47741),
            .in1(N__50345),
            .in2(N__42804),
            .in3(N__36415),
            .lcout(\pid_front.pid_preregZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51316),
            .ce(),
            .sr(N__49621));
    defparam \pid_front.pid_prereg_2_LC_15_23_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_2_LC_15_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_2_LC_15_23_3 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_2_LC_15_23_3  (
            .in0(N__42764),
            .in1(N__48709),
            .in2(N__47699),
            .in3(N__36386),
            .lcout(\pid_front.pid_preregZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51316),
            .ce(),
            .sr(N__49621));
    defparam \pid_front.pid_prereg_15_LC_15_23_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_15_LC_15_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_15_LC_15_23_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pid_front.pid_prereg_15_LC_15_23_5  (
            .in0(N__47753),
            .in1(N__51827),
            .in2(N__42803),
            .in3(N__36355),
            .lcout(\pid_front.pid_preregZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51316),
            .ce(),
            .sr(N__49621));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_15_24_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_15_24_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_15_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37129),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51313),
            .ce(N__48355),
            .sr(N__49623));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_15_24_1 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_15_24_1 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_15_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37048),
            .lcout(drone_H_disp_front_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51313),
            .ce(N__48355),
            .sr(N__49623));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_15_24_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_15_24_2 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_15_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36971),
            .lcout(drone_H_disp_front_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51313),
            .ce(N__48355),
            .sr(N__49623));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_15_24_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_15_24_3 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_15_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36884),
            .lcout(drone_H_disp_front_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51313),
            .ce(N__48355),
            .sr(N__49623));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_15_24_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_15_24_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_15_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36809),
            .lcout(\dron_frame_decoder_1.drone_H_disp_front_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51313),
            .ce(N__48355),
            .sr(N__49623));
    defparam \ppm_encoder_1.rudder_esr_4_LC_16_7_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_4_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_4_LC_16_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_4_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36731),
            .lcout(\ppm_encoder_1.rudderZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51503),
            .ce(N__36688),
            .sr(N__49530));
    defparam \ppm_encoder_1.rudder_esr_5_LC_16_7_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_5_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.rudder_esr_5_LC_16_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.rudder_esr_5_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36713),
            .lcout(\ppm_encoder_1.rudderZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51503),
            .ce(N__36688),
            .sr(N__49530));
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_16_8_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_16_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__41288),
            .in2(N__37346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_16_8_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_1_LC_16_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_1_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__37388),
            .in2(_gnd_net_),
            .in3(N__36635),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_0 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_16_8_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_2_LC_16_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_2_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__40484),
            .in2(N__40442),
            .in3(N__37202),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_1 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_16_8_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_3_LC_16_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_3_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40826),
            .in3(N__37199),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_2 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_16_8_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_4_LC_16_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_4_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__40769),
            .in2(_gnd_net_),
            .in3(N__37196),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_3 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_16_8_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_5_LC_16_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_5_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__40478),
            .in2(_gnd_net_),
            .in3(N__37193),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_4 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_16_8_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_6_LC_16_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_6_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__40490),
            .in2(N__40412),
            .in3(N__37178),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_5 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_16_8_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_7_LC_16_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_7_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__37175),
            .in2(_gnd_net_),
            .in3(N__37151),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_6 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_16_9_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_8_LC_16_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_8_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__37376),
            .in2(_gnd_net_),
            .in3(N__37136),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_8 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_16_9_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_9_LC_16_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_9_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37370),
            .in3(N__37133),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_8 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_16_9_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_10_LC_16_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_10_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__37622),
            .in2(_gnd_net_),
            .in3(N__37295),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_9 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_16_9_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_11_LC_16_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_11_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__37292),
            .in2(_gnd_net_),
            .in3(N__37277),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_10 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_16_9_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_12_LC_16_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_12_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__40865),
            .in2(_gnd_net_),
            .in3(N__37265),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_11 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_16_9_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_13_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_13_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__40496),
            .in2(N__40451),
            .in3(N__37262),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_12 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_16_9_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_14_LC_16_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_14_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__37304),
            .in2(_gnd_net_),
            .in3(N__37259),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_13 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_16_9_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_15_LC_16_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_15_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__44054),
            .in2(_gnd_net_),
            .in3(N__37256),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_14 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_16_10_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_16_LC_16_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_16_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__37253),
            .in2(_gnd_net_),
            .in3(N__37241),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_16 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_16_10_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_17_LC_16_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_17_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__37238),
            .in2(_gnd_net_),
            .in3(N__37226),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_init_pulses_3_cry_16 ),
            .carryout(\ppm_encoder_1.un1_init_pulses_3_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_16_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_18_LC_16_10_2 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_18_LC_16_10_2  (
            .in0(N__45240),
            .in1(N__44835),
            .in2(N__45133),
            .in3(N__37223),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_16_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_16_10_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_16_10_3  (
            .in0(N__44833),
            .in1(_gnd_net_),
            .in2(N__45089),
            .in3(N__44101),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_16_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_16_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_16_10_4  (
            .in0(N__44170),
            .in1(N__45028),
            .in2(_gnd_net_),
            .in3(N__44834),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_16_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_16_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_16_10_5  (
            .in0(N__45029),
            .in1(N__44202),
            .in2(N__44912),
            .in3(N__41443),
            .lcout(\ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_16_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_16_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__45024),
            .in2(_gnd_net_),
            .in3(N__44832),
            .lcout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1 ),
            .ltout(\ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_16_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNILVE13_0_LC_16_10_7 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNILVE13_0_LC_16_10_7  (
            .in0(N__44839),
            .in1(N__41409),
            .in2(N__37349),
            .in3(N__41345),
            .lcout(\ppm_encoder_1.init_pulses_RNILVE13Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_13_LC_16_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_13_LC_16_11_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_13_LC_16_11_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_13_LC_16_11_0  (
            .in0(N__43358),
            .in1(N__37334),
            .in2(N__43239),
            .in3(N__37325),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51456),
            .ce(),
            .sr(N__49558));
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_11_1 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_11_1  (
            .in0(N__40464),
            .in1(_gnd_net_),
            .in2(N__45131),
            .in3(N__44899),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_14_LC_16_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_14_LC_16_11_2 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_14_LC_16_11_2 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_14_LC_16_11_2  (
            .in0(N__43359),
            .in1(N__37319),
            .in2(N__43240),
            .in3(N__37310),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51456),
            .ce(),
            .sr(N__49558));
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_11_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_11_4  (
            .in0(N__44898),
            .in1(N__45078),
            .in2(_gnd_net_),
            .in3(N__37440),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_11_5 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_11_5  (
            .in0(N__37441),
            .in1(N__43757),
            .in2(N__43852),
            .in3(N__41467),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_11_6 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_11_6  (
            .in0(N__41693),
            .in1(N__43835),
            .in2(N__43776),
            .in3(N__40465),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_15_LC_16_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_15_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_15_LC_16_11_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_15_LC_16_11_7  (
            .in0(N__43175),
            .in1(N__37424),
            .in2(N__43374),
            .in3(N__37415),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51456),
            .ce(),
            .sr(N__49558));
    defparam \ppm_encoder_1.init_pulses_0_LC_16_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_0_LC_16_12_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_0_LC_16_12_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.init_pulses_0_LC_16_12_0  (
            .in0(N__43176),
            .in1(N__42032),
            .in2(N__41381),
            .in3(N__43361),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51439),
            .ce(),
            .sr(N__49566));
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_16_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI65N01_0_LC_16_12_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI65N01_0_LC_16_12_1  (
            .in0(N__41405),
            .in1(N__45052),
            .in2(_gnd_net_),
            .in3(N__44858),
            .lcout(\ppm_encoder_1.un1_init_pulses_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_16_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_16_12_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_16_12_2  (
            .in0(N__44861),
            .in1(_gnd_net_),
            .in2(N__45122),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_1_LC_16_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_1_LC_16_12_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_1_LC_16_12_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_1_LC_16_12_3  (
            .in0(N__43360),
            .in1(N__37403),
            .in2(N__43220),
            .in3(N__37394),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51439),
            .ce(),
            .sr(N__49566));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_12_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_12_4  (
            .in0(N__44859),
            .in1(_gnd_net_),
            .in2(N__45121),
            .in3(N__40941),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_16_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_16_12_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_16_12_5  (
            .in0(N__40942),
            .in1(N__45051),
            .in2(_gnd_net_),
            .in3(N__44857),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_10_LC_16_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_10_LC_16_12_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_10_LC_16_12_6 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \ppm_encoder_1.init_pulses_10_LC_16_12_6  (
            .in0(N__43177),
            .in1(N__37640),
            .in2(N__37631),
            .in3(N__43362),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51439),
            .ce(),
            .sr(N__49566));
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_16_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_16_12_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_16_12_7  (
            .in0(N__41167),
            .in1(N__45056),
            .in2(_gnd_net_),
            .in3(N__44860),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_16_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIU1QV2_8_LC_16_13_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIU1QV2_8_LC_16_13_0  (
            .in0(N__37755),
            .in1(N__37606),
            .in2(N__45932),
            .in3(N__45829),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_16_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_16_13_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__44078),
            .in2(N__37574),
            .in3(N__37562),
            .lcout(\ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_16_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIEL7O2_8_LC_16_13_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNIEL7O2_8_LC_16_13_2  (
            .in0(N__37458),
            .in1(N__37512),
            .in2(N__45361),
            .in3(N__45476),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_16_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_16_13_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_16_13_3  (
            .in0(N__37460),
            .in1(N__37756),
            .in2(N__46813),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ppm_encoder_1.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_16_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_16_13_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__46601),
            .in2(N__37556),
            .in3(N__37513),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_8_LC_16_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_8_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_8_LC_16_13_5 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_8_LC_16_13_5  (
            .in0(N__37514),
            .in1(N__37553),
            .in2(N__46387),
            .in3(N__37526),
            .lcout(\ppm_encoder_1.aileronZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51425),
            .ce(),
            .sr(N__49577));
    defparam \ppm_encoder_1.elevator_8_LC_16_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_8_LC_16_13_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_8_LC_16_13_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_8_LC_16_13_6  (
            .in0(N__37459),
            .in1(N__37502),
            .in2(N__46396),
            .in3(N__37472),
            .lcout(\ppm_encoder_1.elevatorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51425),
            .ce(),
            .sr(N__49577));
    defparam \ppm_encoder_1.throttle_8_LC_16_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_8_LC_16_13_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_8_LC_16_13_7 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.throttle_8_LC_16_13_7  (
            .in0(N__37799),
            .in1(N__37757),
            .in2(N__37769),
            .in3(N__46386),
            .lcout(\ppm_encoder_1.throttleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51425),
            .ce(),
            .sr(N__49577));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_0 .LUT_INIT=16'b1100111111011100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_0  (
            .in0(N__45156),
            .in1(N__49784),
            .in2(N__44930),
            .in3(N__41723),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51411),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_14_1 .LUT_INIT=16'b0101010110000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_14_1  (
            .in0(N__43701),
            .in1(N__46806),
            .in2(N__46662),
            .in3(N__41261),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_14_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_14_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_14_2  (
            .in0(N__41262),
            .in1(N__49783),
            .in2(N__37745),
            .in3(N__44786),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51411),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_3  (
            .in0(N__46642),
            .in1(N__44900),
            .in2(N__49797),
            .in3(N__41746),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51411),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_14_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_14_4  (
            .in0(N__37742),
            .in1(N__37710),
            .in2(N__45360),
            .in3(N__45802),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_14_5 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_14_5  (
            .in0(N__37694),
            .in1(N__39207),
            .in2(N__37676),
            .in3(N__45454),
            .lcout(\ppm_encoder_1.elevator_RNIPVQ05Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_14_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_14_6  (
            .in0(N__37661),
            .in1(N__49785),
            .in2(N__40993),
            .in3(N__44787),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51411),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_14_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_14_7 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_14_7  (
            .in0(N__44011),
            .in1(N__45453),
            .in2(N__42059),
            .in3(N__41699),
            .lcout(\ppm_encoder_1.elevator_RNIHNQ05Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_15_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__41720),
            .in2(_gnd_net_),
            .in3(N__41741),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_16_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_16_15_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_16_15_1  (
            .in0(N__44668),
            .in1(N__41113),
            .in2(N__43739),
            .in3(N__49015),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51398),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_16_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI077O2_1_LC_16_15_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI077O2_1_LC_16_15_2  (
            .in0(N__37965),
            .in1(N__45314),
            .in2(N__37951),
            .in3(N__45440),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_16_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIUINC6_1_LC_16_15_3 .LUT_INIT=16'b1110111111101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIUINC6_1_LC_16_15_3  (
            .in0(N__45890),
            .in1(N__37871),
            .in2(N__37928),
            .in3(N__37925),
            .lcout(\ppm_encoder_1.throttle_RNIUINC6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_16_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_16_15_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_16_15_4  (
            .in0(N__37865),
            .in1(N__49014),
            .in2(N__41117),
            .in3(N__44669),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51398),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_15_5 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_15_5  (
            .in0(N__41721),
            .in1(_gnd_net_),
            .in2(N__41747),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_16_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIEES71_1_LC_16_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIEES71_1_LC_16_15_6  (
            .in0(N__37895),
            .in1(N__42175),
            .in2(N__37874),
            .in3(N__44667),
            .lcout(\ppm_encoder_1.throttle_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_16_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_16_15_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__37864),
            .in2(_gnd_net_),
            .in3(N__40983),
            .lcout(\ppm_encoder_1.N_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.source_pid_1_esr_12_LC_16_16_0 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_12_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_12_LC_16_16_0 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \pid_side.source_pid_1_esr_12_LC_16_16_0  (
            .in0(N__38318),
            .in1(N__38398),
            .in2(N__38375),
            .in3(N__37856),
            .lcout(side_order_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51383),
            .ce(N__38090),
            .sr(N__38074));
    defparam \pid_side.source_pid_1_esr_13_LC_16_16_1 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_13_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_13_LC_16_16_1 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \pid_side.source_pid_1_esr_13_LC_16_16_1  (
            .in0(N__38399),
            .in1(N__38371),
            .in2(_gnd_net_),
            .in3(N__38317),
            .lcout(side_order_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51383),
            .ce(N__38090),
            .sr(N__38074));
    defparam \pid_side.source_pid_1_esr_4_LC_16_16_2 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_4_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_4_LC_16_16_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pid_side.source_pid_1_esr_4_LC_16_16_2  (
            .in0(N__38142),
            .in1(N__38200),
            .in2(N__38180),
            .in3(N__38257),
            .lcout(side_order_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51383),
            .ce(N__38090),
            .sr(N__38074));
    defparam \pid_side.source_pid_1_esr_5_LC_16_16_3 .C_ON=1'b0;
    defparam \pid_side.source_pid_1_esr_5_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \pid_side.source_pid_1_esr_5_LC_16_16_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \pid_side.source_pid_1_esr_5_LC_16_16_3  (
            .in0(N__38201),
            .in1(N__38179),
            .in2(_gnd_net_),
            .in3(N__38143),
            .lcout(side_order_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51383),
            .ce(N__38090),
            .sr(N__38074));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_16_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_16_16_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_16_16_4  (
            .in0(N__41263),
            .in1(N__41087),
            .in2(N__41367),
            .in3(N__44666),
            .lcout(\ppm_encoder_1.init_pulses_3_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_16_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_16_16_5 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_16_16_5  (
            .in0(N__45785),
            .in1(N__46415),
            .in2(N__38039),
            .in3(N__41041),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_16_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIFISN6_4_LC_16_16_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIFISN6_4_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__40793),
            .in2(N__38036),
            .in3(N__46889),
            .lcout(\ppm_encoder_1.elevator_RNIFISN6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_16_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_16_16_7 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_16_16_7  (
            .in0(N__38018),
            .in1(N__43642),
            .in2(N__45813),
            .in3(N__45889),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_16_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI8F7O2_5_LC_16_17_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \ppm_encoder_1.elevator_RNI8F7O2_5_LC_16_17_0  (
            .in0(N__39087),
            .in1(N__45423),
            .in2(N__38550),
            .in3(N__45310),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_16_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIKNSN6_5_LC_16_17_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.elevator_RNIKNSN6_5_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__44126),
            .in2(N__37991),
            .in3(N__37988),
            .lcout(\ppm_encoder_1.elevator_RNIKNSN6Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_16_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIQTPV2_6_LC_16_17_2 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIQTPV2_6_LC_16_17_2  (
            .in0(N__38807),
            .in1(N__38776),
            .in2(N__45840),
            .in3(N__45898),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_16_17_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGQOO6_6_LC_16_17_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.throttle_RNIGQOO6_6_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__38750),
            .in2(N__38726),
            .in3(N__38708),
            .lcout(\ppm_encoder_1.throttle_RNIGQOO6Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_16_17_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIAH7O2_6_LC_16_17_4 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.elevator_RNIAH7O2_6_LC_16_17_4  (
            .in0(N__39144),
            .in1(N__45422),
            .in2(N__38653),
            .in3(N__45309),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_6_LC_16_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_6_LC_16_17_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_6_LC_16_17_7 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ppm_encoder_1.aileron_6_LC_16_17_7  (
            .in0(N__38652),
            .in1(N__46328),
            .in2(N__38702),
            .in3(N__38669),
            .lcout(\ppm_encoder_1.aileronZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51371),
            .ce(),
            .sr(N__49603));
    defparam \ppm_encoder_1.aileron_3_LC_16_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_3_LC_16_18_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_3_LC_16_18_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \ppm_encoder_1.aileron_3_LC_16_18_0  (
            .in0(N__38630),
            .in1(N__38613),
            .in2(N__46374),
            .in3(N__42277),
            .lcout(\ppm_encoder_1.aileronZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.aileron_5_LC_16_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_5_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_5_LC_16_18_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.aileron_5_LC_16_18_1  (
            .in0(N__38594),
            .in1(N__38578),
            .in2(N__38554),
            .in3(N__46340),
            .lcout(\ppm_encoder_1.aileronZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.aileron_9_LC_16_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_9_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_9_LC_16_18_2 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.aileron_9_LC_16_18_2  (
            .in0(N__38525),
            .in1(N__38498),
            .in2(N__46375),
            .in3(N__38479),
            .lcout(\ppm_encoder_1.aileronZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.elevator_10_LC_16_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_10_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_10_LC_16_18_3 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \ppm_encoder_1.elevator_10_LC_16_18_3  (
            .in0(N__38460),
            .in1(N__38435),
            .in2(N__38428),
            .in3(N__46341),
            .lcout(\ppm_encoder_1.elevatorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.elevator_2_LC_16_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_2_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_2_LC_16_18_4 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.elevator_2_LC_16_18_4  (
            .in0(N__46332),
            .in1(N__39251),
            .in2(N__39215),
            .in3(N__39221),
            .lcout(\ppm_encoder_1.elevatorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.elevator_6_LC_16_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_6_LC_16_18_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_6_LC_16_18_5 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ppm_encoder_1.elevator_6_LC_16_18_5  (
            .in0(N__39185),
            .in1(N__39148),
            .in2(N__39179),
            .in3(N__46342),
            .lcout(\ppm_encoder_1.elevatorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \ppm_encoder_1.elevator_5_LC_16_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_5_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_5_LC_16_18_6 .LUT_INIT=16'b0111001011011000;
    LogicCell40 \ppm_encoder_1.elevator_5_LC_16_18_6  (
            .in0(N__46333),
            .in1(N__39128),
            .in2(N__39097),
            .in3(N__39104),
            .lcout(\ppm_encoder_1.elevatorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51359),
            .ce(),
            .sr(N__49608));
    defparam \Commands_frame_decoder.source_xy_kp_1_e_0_4_LC_16_19_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_xy_kp_1_e_0_4_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_xy_kp_1_e_0_4_LC_16_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_xy_kp_1_e_0_4_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__40255),
            .in2(_gnd_net_),
            .in3(N__50797),
            .lcout(xy_kp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51349),
            .ce(N__39032),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_4_LC_16_20_5 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_4_LC_16_20_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_4_LC_16_20_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_4_LC_16_20_5  (
            .in0(N__42814),
            .in1(N__48626),
            .in2(N__47663),
            .in3(N__38961),
            .lcout(\pid_front.pid_preregZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51341),
            .ce(),
            .sr(N__49616));
    defparam \pid_front.pid_prereg_5_LC_16_21_1 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_5_LC_16_21_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_5_LC_16_21_1 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pid_front.pid_prereg_5_LC_16_21_1  (
            .in0(N__42810),
            .in1(N__48671),
            .in2(N__47645),
            .in3(N__38924),
            .lcout(\pid_front.pid_preregZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51334),
            .ce(),
            .sr(N__49619));
    defparam \pid_front.pid_prereg_3_LC_16_21_3 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_3_LC_16_21_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_3_LC_16_21_3 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pid_front.pid_prereg_3_LC_16_21_3  (
            .in0(N__42809),
            .in1(N__50384),
            .in2(N__47681),
            .in3(N__38892),
            .lcout(\pid_front.pid_preregZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51334),
            .ce(),
            .sr(N__49619));
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_16_22_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_alt_ki_6_LC_16_22_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Commands_frame_decoder.source_alt_ki_6_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__40139),
            .in2(_gnd_net_),
            .in3(N__50796),
            .lcout(alt_ki_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51327),
            .ce(N__38855),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_16_22_3 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_16_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43468),
            .lcout(drone_H_disp_front_i_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_16_22_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_16_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39794),
            .lcout(drone_H_disp_front_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_16_22_5 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_16_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39788),
            .lcout(drone_H_disp_front_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_16_22_6 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_16_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39782),
            .lcout(drone_H_disp_front_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_16_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_16_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39776),
            .lcout(drone_H_disp_front_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_16_23_0 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_0_LC_16_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_0_LC_16_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39760),
            .lcout(front_command_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_16_23_1 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_16_23_1 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_1_LC_16_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_1_LC_16_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39651),
            .lcout(front_command_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_16_23_2 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_16_23_2 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_2_LC_16_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_2_LC_16_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39512),
            .lcout(front_command_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_16_23_3 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_16_23_3 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_3_LC_16_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_3_LC_16_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39363),
            .lcout(front_command_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_16_23_4 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_16_23_4 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_4_LC_16_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_4_LC_16_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40403),
            .lcout(front_command_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_16_23_5 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_16_23_5 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_5_LC_16_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_5_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40256),
            .lcout(front_command_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_16_23_6 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_16_23_6 .SEQ_MODE=4'b1000;
    defparam \Commands_frame_decoder.source_CH3data_esr_6_LC_16_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_esr_6_LC_16_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40140),
            .lcout(front_command_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_16_23_7 .C_ON=1'b0;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_16_23_7 .SEQ_MODE=4'b1001;
    defparam \Commands_frame_decoder.source_CH3data_ess_7_LC_16_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Commands_frame_decoder.source_CH3data_ess_7_LC_16_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39993),
            .lcout(front_command_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51320),
            .ce(N__39884),
            .sr(N__49624));
    defparam \pid_front.error_axb_7_LC_16_24_0 .C_ON=1'b0;
    defparam \pid_front.error_axb_7_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_7_LC_16_24_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \pid_front.error_axb_7_LC_16_24_0  (
            .in0(N__39853),
            .in1(N__39844),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pid_front.error_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_16_24_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_16_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_16_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39866),
            .lcout(drone_H_disp_front_i_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_16_24_4 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_16_24_4 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_16_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_16_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39860),
            .lcout(drone_H_disp_front_i_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_axb_8_l_ofx_LC_16_24_6 .C_ON=1'b0;
    defparam \pid_front.error_axb_8_l_ofx_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_axb_8_l_ofx_LC_16_24_6 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \pid_front.error_axb_8_l_ofx_LC_16_24_6  (
            .in0(N__39854),
            .in1(N__39845),
            .in2(_gnd_net_),
            .in3(N__43518),
            .lcout(\pid_front.error_axb_8_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_pc.data_Aux_6_LC_17_8_0 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_6_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_6_LC_17_8_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \uart_pc.data_Aux_6_LC_17_8_0  (
            .in0(N__39836),
            .in1(N__40707),
            .in2(N__39811),
            .in3(N__40759),
            .lcout(\uart_pc.data_AuxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51504),
            .ce(),
            .sr(N__40532));
    defparam \uart_pc.data_Aux_7_LC_17_8_1 .C_ON=1'b0;
    defparam \uart_pc.data_Aux_7_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_pc.data_Aux_7_LC_17_8_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \uart_pc.data_Aux_7_LC_17_8_1  (
            .in0(N__40760),
            .in1(N__40543),
            .in2(N__40712),
            .in3(N__40589),
            .lcout(\uart_pc.data_AuxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51504),
            .ce(),
            .sr(N__40532));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_17_8_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_17_8_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_17_8_4  (
            .in0(N__44926),
            .in1(_gnd_net_),
            .in2(N__41344),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_17_8_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_17_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__41337),
            .in2(_gnd_net_),
            .in3(N__44925),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_17_8_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_17_8_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__41372),
            .in2(_gnd_net_),
            .in3(N__42182),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_17_9_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_17_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__41325),
            .in2(_gnd_net_),
            .in3(N__44848),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_9_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_9_1  (
            .in0(N__44849),
            .in1(N__43903),
            .in2(_gnd_net_),
            .in3(N__45124),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_17_9_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_17_9_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_17_9_2  (
            .in0(N__41441),
            .in1(N__41326),
            .in2(N__40472),
            .in3(N__44853),
            .lcout(\ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_9_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_9_3  (
            .in0(N__41327),
            .in1(N__40924),
            .in2(N__44913),
            .in3(N__41439),
            .lcout(\ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_9_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_9_4  (
            .in0(N__41440),
            .in1(N__41328),
            .in2(N__44933),
            .in3(N__40433),
            .lcout(\ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_17_9_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_17_9_5 .LUT_INIT=16'b1101110011011110;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_17_9_5  (
            .in0(N__44852),
            .in1(N__49782),
            .in2(N__46582),
            .in3(N__45127),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNELZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51492),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_9_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_9_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_9_6  (
            .in0(N__45125),
            .in1(N__40888),
            .in2(_gnd_net_),
            .in3(N__44850),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_17_9_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_2_18_LC_17_9_7 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_2_18_LC_17_9_7  (
            .in0(N__44851),
            .in1(N__41442),
            .in2(N__45253),
            .in3(N__45126),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_3_LC_17_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_3_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.init_pulses_3_LC_17_10_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_3_LC_17_10_0  (
            .in0(N__43308),
            .in1(N__40847),
            .in2(N__43219),
            .in3(N__40838),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51483),
            .ce(),
            .sr(N__49559));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_17_10_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_17_10_1 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_17_10_1  (
            .in0(N__44842),
            .in1(N__41221),
            .in2(N__45090),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_17_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNI98N01_3_LC_17_10_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNI98N01_3_LC_17_10_2  (
            .in0(N__41220),
            .in1(N__45031),
            .in2(_gnd_net_),
            .in3(N__44841),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_4_LC_17_10_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_4_LC_17_10_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_4_LC_17_10_3 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \ppm_encoder_1.init_pulses_4_LC_17_10_3  (
            .in0(N__40814),
            .in1(N__40802),
            .in2(N__43244),
            .in3(N__43309),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51483),
            .ce(),
            .sr(N__49559));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_17_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_17_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_17_10_4  (
            .in0(N__41052),
            .in1(N__45030),
            .in2(_gnd_net_),
            .in3(N__44840),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_10_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_10_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_10_5  (
            .in0(N__44843),
            .in1(_gnd_net_),
            .in2(N__45091),
            .in3(N__41053),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_10_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_10_6  (
            .in0(N__41054),
            .in1(N__43839),
            .in2(N__43783),
            .in3(N__41042),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_5_LC_17_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_10_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_5_LC_17_10_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \ppm_encoder_1.init_pulses_5_LC_17_10_7  (
            .in0(N__41018),
            .in1(N__43178),
            .in2(N__41006),
            .in3(N__43310),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51483),
            .ce(),
            .sr(N__49559));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_17_11_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_17_11_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_17_11_0  (
            .in0(N__46752),
            .in1(N__41270),
            .in2(_gnd_net_),
            .in3(N__42219),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_17_11_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_17_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__41077),
            .in2(_gnd_net_),
            .in3(N__40994),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_11_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_11_2 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__40967),
            .in2(N__40946),
            .in3(N__44896),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_17_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_17_11_3 .LUT_INIT=16'b1101110111010001;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_17_11_3  (
            .in0(N__41192),
            .in1(N__43831),
            .in2(N__43777),
            .in3(N__40943),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_17_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_17_11_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_17_11_4  (
            .in0(N__46754),
            .in1(N__43762),
            .in2(N__46645),
            .in3(N__45085),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_ns_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_17_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_17_11_5 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_17_11_5  (
            .in0(N__42220),
            .in1(_gnd_net_),
            .in2(N__41276),
            .in3(N__46753),
            .lcout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux ),
            .ltout(\ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_17_11_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_17_11_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_17_11_6  (
            .in0(N__43832),
            .in1(N__43761),
            .in2(N__40928),
            .in3(N__40925),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_17_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_17_11_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_17_11_7  (
            .in0(N__44897),
            .in1(N__45211),
            .in2(_gnd_net_),
            .in3(N__41323),
            .lcout(\ppm_encoder_1.un1_init_pulses_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_12_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_12_0 .LUT_INIT=16'b1001011001011010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_12_0  (
            .in0(N__41447),
            .in1(N__41324),
            .in2(N__41417),
            .in3(N__44846),
            .lcout(\ppm_encoder_1.un1_init_pulses_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_17_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_17_12_1 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_17_12_1  (
            .in0(N__45023),
            .in1(N__41081),
            .in2(N__41274),
            .in3(N__41368),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1 ),
            .ltout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_17_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_17_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41291),
            .in3(N__44844),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_17_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_17_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_17_12_3  (
            .in0(N__41083),
            .in1(N__43954),
            .in2(N__41275),
            .in3(N__42221),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_153_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_17_12_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_17_12_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__49764),
            .in2(_gnd_net_),
            .in3(N__44845),
            .lcout(\ppm_encoder_1.N_1818_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_12_5 .LUT_INIT=16'b1100111110001011;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_12_5  (
            .in0(N__41225),
            .in1(N__43834),
            .in2(N__41202),
            .in3(N__43749),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_12_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_12_6  (
            .in0(N__43833),
            .in1(N__41168),
            .in2(N__43772),
            .in3(N__41150),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_17_12_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_17_12_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_17_12_7  (
            .in0(N__44847),
            .in1(N__49010),
            .in2(N__41107),
            .in3(N__41082),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51457),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_17_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIM4PT2_13_LC_17_13_0 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \ppm_encoder_1.throttle_RNIM4PT2_13_LC_17_13_0  (
            .in0(N__41692),
            .in1(N__45924),
            .in2(N__41486),
            .in3(N__45830),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_17_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIMC2D6_13_LC_17_13_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ppm_encoder_1.elevator_RNIMC2D6_13_LC_17_13_1  (
            .in0(N__41663),
            .in1(_gnd_net_),
            .in2(N__41648),
            .in3(N__41630),
            .lcout(\ppm_encoder_1.elevator_RNIMC2D6Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_17_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI68LH2_13_LC_17_13_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.elevator_RNI68LH2_13_LC_17_13_2  (
            .in0(N__41529),
            .in1(N__41580),
            .in2(N__45362),
            .in3(N__45478),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_17_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_17_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_17_13_3  (
            .in0(N__41484),
            .in1(N__46805),
            .in2(_gnd_net_),
            .in3(N__41530),
            .lcout(),
            .ltout(\ppm_encoder_1.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_17_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_17_13_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_17_13_4  (
            .in0(N__46583),
            .in1(_gnd_net_),
            .in2(N__41624),
            .in3(N__41581),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_13_LC_17_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_13_LC_17_13_5 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_13_LC_17_13_5 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ppm_encoder_1.aileron_13_LC_17_13_5  (
            .in0(N__41582),
            .in1(N__46376),
            .in2(N__41620),
            .in3(N__41594),
            .lcout(\ppm_encoder_1.aileronZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51440),
            .ce(),
            .sr(N__49585));
    defparam \ppm_encoder_1.elevator_13_LC_17_13_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_13_LC_17_13_6 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.elevator_13_LC_17_13_6 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.elevator_13_LC_17_13_6  (
            .in0(N__41531),
            .in1(N__41570),
            .in2(N__46394),
            .in3(N__41546),
            .lcout(\ppm_encoder_1.elevatorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51440),
            .ce(),
            .sr(N__49585));
    defparam \ppm_encoder_1.throttle_13_LC_17_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_13_LC_17_13_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_13_LC_17_13_7 .LUT_INIT=16'b1100101000111010;
    LogicCell40 \ppm_encoder_1.throttle_13_LC_17_13_7  (
            .in0(N__41485),
            .in1(N__41519),
            .in2(N__46395),
            .in3(N__41495),
            .lcout(\ppm_encoder_1.throttleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51440),
            .ce(),
            .sr(N__49585));
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_17_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_17_14_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_17_14_0  (
            .in0(N__41815),
            .in1(N__41468),
            .in2(N__45831),
            .in3(N__45925),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_17_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_17_14_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__41858),
            .in2(N__41840),
            .in3(N__41822),
            .lcout(\ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_17_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_17_14_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_17_14_2  (
            .in0(N__41797),
            .in1(N__41779),
            .in2(N__45499),
            .in3(N__45352),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_17_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_17_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_17_14_3  (
            .in0(N__46814),
            .in1(N__41816),
            .in2(_gnd_net_),
            .in3(N__41798),
            .lcout(),
            .ltout(\ppm_encoder_1.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_14_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_14_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_14_4  (
            .in0(N__46643),
            .in1(_gnd_net_),
            .in2(N__41783),
            .in3(N__41780),
            .lcout(),
            .ltout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_17_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_14_LC_17_14_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_14_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__44473),
            .in2(N__41765),
            .in3(N__41762),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51426),
            .ce(N__44408),
            .sr(N__49594));
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_14_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_14_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_14_6  (
            .in0(N__47501),
            .in1(N__44188),
            .in2(N__47474),
            .in3(N__41753),
            .lcout(\ppm_encoder_1.counter24_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_17_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_17_15_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_17_15_0  (
            .in0(N__41745),
            .in1(N__41722),
            .in2(N__44725),
            .in3(N__42174),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_0 ),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_17_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIGCMK2_0_LC_17_15_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.throttle_RNIGCMK2_0_LC_17_15_1  (
            .in0(N__43979),
            .in1(N__45993),
            .in2(N__41702),
            .in3(N__45304),
            .lcout(\ppm_encoder_1.un2_throttle_iv_0_0 ),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_15_2 .LUT_INIT=16'b0010111111010000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_15_2  (
            .in0(N__45448),
            .in1(N__44012),
            .in2(N__42062),
            .in3(N__42058),
            .lcout(\ppm_encoder_1.un1_init_pulses_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_17_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_17_15_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_17_15_3  (
            .in0(N__44722),
            .in1(N__46644),
            .in2(N__49799),
            .in3(N__43953),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51412),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_17_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_17_15_5 .LUT_INIT=16'b1111010111110010;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_17_15_5  (
            .in0(N__44723),
            .in1(N__45161),
            .in2(N__49798),
            .in3(N__42217),
            .lcout(\ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51412),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_17_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNIMIMK2_3_LC_17_15_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \ppm_encoder_1.throttle_RNIMIMK2_3_LC_17_15_6  (
            .in0(N__42020),
            .in1(N__42278),
            .in2(N__45338),
            .in3(N__45786),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_17_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNIT3R05_3_LC_17_15_7 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \ppm_encoder_1.elevator_RNIT3R05_3_LC_17_15_7  (
            .in0(N__41995),
            .in1(N__41975),
            .in2(N__41942),
            .in3(N__45447),
            .lcout(\ppm_encoder_1.elevator_RNIT3R05Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.pid_prereg_esr_0_LC_17_16_1 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_esr_0_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_esr_0_LC_17_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_side.pid_prereg_esr_0_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48296),
            .lcout(\pid_side.pid_preregZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51399),
            .ce(N__41890),
            .sr(N__49604));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_17_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_17_16_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_17_16_2  (
            .in0(N__42173),
            .in1(N__43946),
            .in2(N__42218),
            .in3(N__42420),
            .lcout(),
            .ltout(\ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_17_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_17_16_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_17_16_3  (
            .in0(N__47173),
            .in1(_gnd_net_),
            .in2(N__41861),
            .in3(_gnd_net_),
            .lcout(\ppm_encoder_1.init_pulses_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_17_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_17_16_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__42419),
            .in2(_gnd_net_),
            .in3(N__42086),
            .lcout(\ppm_encoder_1.PPM_STATE_53_d ),
            .ltout(\ppm_encoder_1.PPM_STATE_53_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_17_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_17_16_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_17_16_5  (
            .in0(N__43944),
            .in1(N__42204),
            .in2(N__42236),
            .in3(N__42171),
            .lcout(\ppm_encoder_1.init_pulses_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_16_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(N__47174),
            .in2(_gnd_net_),
            .in3(N__42421),
            .lcout(\ppm_encoder_1.N_134_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_17_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_17_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_17_16_7  (
            .in0(N__43945),
            .in1(N__42205),
            .in2(N__44724),
            .in3(N__42172),
            .lcout(\ppm_encoder_1.init_pulses_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_17_17_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_17_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_17_17_0  (
            .in0(N__42829),
            .in1(N__42068),
            .in2(N__42854),
            .in3(N__47086),
            .lcout(\ppm_encoder_1.N_232 ),
            .ltout(\ppm_encoder_1.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_17_17_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_17_17_1 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_17_17_1  (
            .in0(N__49038),
            .in1(N__47163),
            .in2(N__42146),
            .in3(N__42423),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_17_17_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_1_LC_17_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_1_LC_17_17_2  (
            .in0(N__42830),
            .in1(N__47087),
            .in2(N__42395),
            .in3(N__42853),
            .lcout(\ppm_encoder_1.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_0_LC_17_17_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_17_17_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_0_LC_17_17_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \ppm_encoder_1.PPM_STATE_0_LC_17_17_6  (
            .in0(N__42424),
            .in1(N__42112),
            .in2(N__47172),
            .in3(N__42097),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51384),
            .ce(),
            .sr(N__49609));
    defparam \ppm_encoder_1.PPM_STATE_1_LC_17_17_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.PPM_STATE_1_LC_17_17_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ppm_encoder_1.PPM_STATE_1_LC_17_17_7  (
            .in0(N__42113),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42425),
            .lcout(\ppm_encoder_1.PPM_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51384),
            .ce(),
            .sr(N__49609));
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_17_18_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_17_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_17_18_0  (
            .in0(N__47364),
            .in1(N__46977),
            .in2(N__46958),
            .in3(N__42087),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_17_18_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.ppm_output_reg_RNO_2_LC_17_18_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \ppm_encoder_1.ppm_output_reg_RNO_2_LC_17_18_1  (
            .in0(N__46978),
            .in1(N__47365),
            .in2(N__46954),
            .in3(N__42422),
            .lcout(\ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_18_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_18_2  (
            .in0(N__42359),
            .in1(N__47363),
            .in2(N__42341),
            .in3(N__46946),
            .lcout(\ppm_encoder_1.counter24_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_2_LC_17_18_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_2_LC_17_18_3  (
            .in0(N__42386),
            .in1(N__44490),
            .in2(_gnd_net_),
            .in3(N__42371),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51372),
            .ce(N__44411),
            .sr(N__49612));
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_18_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_3_LC_17_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_3_LC_17_18_4  (
            .in0(N__44488),
            .in1(N__42242),
            .in2(_gnd_net_),
            .in3(N__42353),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51372),
            .ce(N__44411),
            .sr(N__49612));
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_17_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_17_18_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_0_LC_17_18_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_0_LC_17_18_5  (
            .in0(N__43919),
            .in1(N__44489),
            .in2(_gnd_net_),
            .in3(N__42332),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51372),
            .ce(N__44411),
            .sr(N__49612));
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_17_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_17_18_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_17_18_6  (
            .in0(N__42320),
            .in1(N__46976),
            .in2(N__42287),
            .in3(N__46995),
            .lcout(\ppm_encoder_1.counter24_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_17_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_17_18_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_1_LC_17_18_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_1_LC_17_18_7  (
            .in0(N__42314),
            .in1(N__42302),
            .in2(_gnd_net_),
            .in3(N__44491),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51372),
            .ce(N__44411),
            .sr(N__49612));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_17_19_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_17_19_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_17_19_1  (
            .in0(N__42276),
            .in1(_gnd_net_),
            .in2(N__46655),
            .in3(N__42257),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_17_19_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIUS1G_4_LC_17_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNIUS1G_4_LC_17_19_4  (
            .in0(N__47298),
            .in1(N__47320),
            .in2(N__47275),
            .in3(N__47341),
            .lcout(),
            .ltout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_17_19_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIAEV01_8_LC_17_19_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ppm_encoder_1.counter_RNIAEV01_8_LC_17_19_5  (
            .in0(N__42836),
            .in1(N__47547),
            .in2(N__42857),
            .in3(N__47244),
            .lcout(\ppm_encoder_1.N_139_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_17_19_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_17_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44826),
            .lcout(\ppm_encoder_1.N_1818_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_17_20_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIDBJ8_13_LC_17_20_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ppm_encoder_1.counter_RNIDBJ8_13_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__47496),
            .in2(_gnd_net_),
            .in3(N__47523),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_17_20_2 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_17_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43525),
            .lcout(drone_H_disp_front_i_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7  (
            .in0(N__47418),
            .in1(N__47442),
            .in2(N__47393),
            .in3(N__47466),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_8_LC_17_21_0 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_8_LC_17_21_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_8_LC_17_21_0 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pid_front.pid_prereg_8_LC_17_21_0  (
            .in0(N__47600),
            .in1(N__50495),
            .in2(N__42818),
            .in3(N__42630),
            .lcout(\pid_front.pid_preregZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51342),
            .ce(),
            .sr(N__49622));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_17_22_7 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_17_22_7 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_17_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42610),
            .lcout(drone_H_disp_front_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51335),
            .ce(N__42527),
            .sr(N__49625));
    defparam \pid_front.error_cry_0_c_inv_LC_17_23_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_inv_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_inv_LC_17_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pid_front.error_cry_0_c_inv_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__42461),
            .in2(_gnd_net_),
            .in3(N__42472),
            .lcout(\pid_front.error_axb_0 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\pid_front.error_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_17_23_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_c_RNIC7KB_LC_17_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_0_c_RNIC7KB_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__42455),
            .in2(_gnd_net_),
            .in3(N__42428),
            .lcout(\pid_front.error_1 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0 ),
            .carryout(\pid_front.error_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_17_23_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_c_RNIEALB_LC_17_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_1_c_RNIEALB_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__43088),
            .in2(_gnd_net_),
            .in3(N__43064),
            .lcout(\pid_front.error_2 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1 ),
            .carryout(\pid_front.error_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_17_23_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_c_RNIGDMB_LC_17_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_2_c_RNIGDMB_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__43061),
            .in2(_gnd_net_),
            .in3(N__43031),
            .lcout(\pid_front.error_3 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2 ),
            .carryout(\pid_front.error_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_17_23_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_c_RNIABAG_LC_17_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_c_RNIABAG_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__43028),
            .in2(N__43022),
            .in3(N__42998),
            .lcout(\pid_front.error_4 ),
            .ltout(),
            .carryin(\pid_front.error_cry_3 ),
            .carryout(\pid_front.error_cry_0_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_17_23_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_0_0_c_RNIOQKB_LC_17_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_0_0_c_RNIOQKB_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__42995),
            .in2(N__42989),
            .in3(N__42965),
            .lcout(\pid_front.error_5 ),
            .ltout(),
            .carryin(\pid_front.error_cry_0_0 ),
            .carryout(\pid_front.error_cry_1_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_17_23_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_1_0_c_RNIR0RF_LC_17_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_1_0_c_RNIR0RF_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(N__42962),
            .in2(N__42956),
            .in3(N__42932),
            .lcout(\pid_front.error_6 ),
            .ltout(),
            .carryin(\pid_front.error_cry_1_0 ),
            .carryout(\pid_front.error_cry_2_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_17_23_7 .C_ON=1'b1;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_17_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_2_0_c_RNIU61K_LC_17_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_2_0_c_RNIU61K_LC_17_23_7  (
            .in0(_gnd_net_),
            .in1(N__42929),
            .in2(N__42923),
            .in3(N__42899),
            .lcout(\pid_front.error_7 ),
            .ltout(),
            .carryin(\pid_front.error_cry_2_0 ),
            .carryout(\pid_front.error_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_17_24_0 .C_ON=1'b1;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_17_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_3_0_c_RNI1D7O_LC_17_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_3_0_c_RNI1D7O_LC_17_24_0  (
            .in0(_gnd_net_),
            .in1(N__42896),
            .in2(N__42890),
            .in3(N__42860),
            .lcout(\pid_front.error_8 ),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(\pid_front.error_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_17_24_1 .C_ON=1'b1;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_17_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_4_c_RNILNBG_LC_17_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_4_c_RNILNBG_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__43625),
            .in2(N__43619),
            .in3(N__43598),
            .lcout(\pid_front.error_9 ),
            .ltout(),
            .carryin(\pid_front.error_cry_4 ),
            .carryout(\pid_front.error_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_17_24_2 .C_ON=1'b1;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_5_c_RNIVNFF_LC_17_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_5_c_RNIVNFF_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__43595),
            .in2(N__43586),
            .in3(N__43562),
            .lcout(\pid_front.error_10 ),
            .ltout(),
            .carryin(\pid_front.error_cry_5 ),
            .carryout(\pid_front.error_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_17_24_3 .C_ON=1'b1;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_17_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_6_c_RNI3VJG_LC_17_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pid_front.error_cry_6_c_RNI3VJG_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(N__43559),
            .in2(_gnd_net_),
            .in3(N__43538),
            .lcout(\pid_front.error_11 ),
            .ltout(),
            .carryin(\pid_front.error_cry_6 ),
            .carryout(\pid_front.error_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_17_24_4 .C_ON=1'b1;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_17_24_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_7_c_RNIAPPM_LC_17_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_7_c_RNIAPPM_LC_17_24_4  (
            .in0(_gnd_net_),
            .in1(N__43535),
            .in2(N__43529),
            .in3(N__43484),
            .lcout(\pid_front.error_12 ),
            .ltout(),
            .carryin(\pid_front.error_cry_7 ),
            .carryout(\pid_front.error_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_17_24_5 .C_ON=1'b1;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_17_24_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_8_c_RNIAC2E_LC_17_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_8_c_RNIAC2E_LC_17_24_5  (
            .in0(_gnd_net_),
            .in1(N__43481),
            .in2(N__43472),
            .in3(N__43436),
            .lcout(\pid_front.error_13 ),
            .ltout(),
            .carryin(\pid_front.error_cry_8 ),
            .carryout(\pid_front.error_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_17_24_6 .C_ON=1'b1;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_17_24_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_9_c_RNIDG3E_LC_17_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pid_front.error_cry_9_c_RNIDG3E_LC_17_24_6  (
            .in0(_gnd_net_),
            .in1(N__43433),
            .in2(N__48371),
            .in3(N__43409),
            .lcout(\pid_front.error_14 ),
            .ltout(),
            .carryin(\pid_front.error_cry_9 ),
            .carryout(\pid_front.error_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_17_24_7 .C_ON=1'b0;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.error_cry_10_c_RNINTDI_LC_17_24_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \pid_front.error_cry_10_c_RNINTDI_LC_17_24_7  (
            .in0(N__43406),
            .in1(N__48370),
            .in2(_gnd_net_),
            .in3(N__43394),
            .lcout(\pid_front.error_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_9_LC_18_10_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_9_LC_18_10_0 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.init_pulses_9_LC_18_10_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \ppm_encoder_1.init_pulses_9_LC_18_10_0  (
            .in0(N__43372),
            .in1(N__43256),
            .in2(N__43218),
            .in3(N__43100),
            .lcout(\ppm_encoder_1.init_pulsesZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51493),
            .ce(),
            .sr(N__49567));
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_18_10_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_18_10_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_18_10_2  (
            .in0(N__44163),
            .in1(N__45061),
            .in2(_gnd_net_),
            .in3(N__44922),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_10_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_10_4  (
            .in0(N__43902),
            .in1(N__45060),
            .in2(_gnd_net_),
            .in3(N__44921),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_18_10_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_18_10_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_18_10_6  (
            .in0(N__44100),
            .in1(N__45062),
            .in2(_gnd_net_),
            .in3(N__44923),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_10_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_10_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_10_7  (
            .in0(N__44924),
            .in1(_gnd_net_),
            .in2(N__45123),
            .in3(N__44215),
            .lcout(\ppm_encoder_1.un1_init_pulses_3_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_0_LC_18_11_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_0_LC_18_11_3 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.throttle_0_LC_18_11_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \ppm_encoder_1.throttle_0_LC_18_11_3  (
            .in0(N__43978),
            .in1(N__46190),
            .in2(_gnd_net_),
            .in3(N__44042),
            .lcout(\ppm_encoder_1.throttleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51484),
            .ce(),
            .sr(N__49578));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_18_11_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_18_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_18_11_4  (
            .in0(N__44010),
            .in1(N__43977),
            .in2(_gnd_net_),
            .in3(N__43958),
            .lcout(),
            .ltout(\ppm_encoder_1.N_286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_18_11_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_18_11_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__46538),
            .in2(N__43922),
            .in3(N__46001),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_11_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_11_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_11_7  (
            .in0(N__43904),
            .in1(N__43840),
            .in2(N__43778),
            .in3(N__43646),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_18_12_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_4_LC_18_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_4_LC_18_12_1  (
            .in0(N__44501),
            .in1(N__46466),
            .in2(_gnd_net_),
            .in3(N__44357),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51471),
            .ce(N__44404),
            .sr(N__49586));
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_18_12_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_5_LC_18_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_5_LC_18_12_2  (
            .in0(N__44348),
            .in1(N__44342),
            .in2(_gnd_net_),
            .in3(N__44503),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51471),
            .ce(N__44404),
            .sr(N__49586));
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_12_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_10_LC_18_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_10_LC_18_12_3  (
            .in0(N__44499),
            .in1(N__44327),
            .in2(_gnd_net_),
            .in3(N__44315),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51471),
            .ce(N__44404),
            .sr(N__49586));
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_12_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_11_LC_18_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_11_LC_18_12_5  (
            .in0(N__44500),
            .in1(N__44309),
            .in2(_gnd_net_),
            .in3(N__44300),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51471),
            .ce(N__44404),
            .sr(N__49586));
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_12_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_12_LC_18_12_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_12_LC_18_12_6  (
            .in0(N__44288),
            .in1(N__44502),
            .in2(_gnd_net_),
            .in3(N__44276),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51471),
            .ce(N__44404),
            .sr(N__49586));
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_18_13_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_18_13_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_18_13_0  (
            .in0(N__44260),
            .in1(N__47420),
            .in2(N__44230),
            .in3(N__47444),
            .lcout(\ppm_encoder_1.counter24_0_I_51_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_16_LC_18_13_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_16_LC_18_13_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_16_LC_18_13_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_16_LC_18_13_1  (
            .in0(N__45182),
            .in1(N__44261),
            .in2(N__45221),
            .in3(N__44831),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51458),
            .ce(),
            .sr(N__49595));
    defparam \ppm_encoder_1.pulses2count_17_LC_18_13_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_17_LC_18_13_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_17_LC_18_13_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_17_LC_18_13_2  (
            .in0(N__44828),
            .in1(N__45218),
            .in2(N__44231),
            .in3(N__44252),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51458),
            .ce(),
            .sr(N__49595));
    defparam \ppm_encoder_1.pulses2count_15_LC_18_13_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_15_LC_18_13_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_15_LC_18_13_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ppm_encoder_1.pulses2count_15_LC_18_13_3  (
            .in0(N__44216),
            .in1(N__44189),
            .in2(N__45220),
            .in3(N__44830),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51458),
            .ce(),
            .sr(N__49595));
    defparam \ppm_encoder_1.pulses2count_18_LC_18_13_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_18_LC_18_13_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_18_LC_18_13_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ppm_encoder_1.pulses2count_18_LC_18_13_4  (
            .in0(N__44829),
            .in1(N__45254),
            .in2(N__45194),
            .in3(N__45219),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51458),
            .ce(),
            .sr(N__49595));
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_18_13_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_18_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_18_13_5  (
            .in0(N__47392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45190),
            .lcout(\ppm_encoder_1.counter24_0_I_57_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_18_13_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_18_13_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_18_13_7  (
            .in0(N__45181),
            .in1(N__45132),
            .in2(_gnd_net_),
            .in3(N__44827),
            .lcout(\ppm_encoder_1.un1_init_pulses_0_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_14_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_14_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_14_0  (
            .in0(N__44564),
            .in1(N__47276),
            .in2(N__44543),
            .in3(N__47300),
            .lcout(\ppm_encoder_1.counter24_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_14_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_6_LC_18_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_6_LC_18_14_1  (
            .in0(N__44492),
            .in1(N__44588),
            .in2(_gnd_net_),
            .in3(N__44579),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51441),
            .ce(N__44409),
            .sr(N__49599));
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_14_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_14_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_7_LC_18_14_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_7_LC_18_14_2  (
            .in0(N__45683),
            .in1(N__44494),
            .in2(_gnd_net_),
            .in3(N__44558),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51441),
            .ce(N__44409),
            .sr(N__49599));
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_18_14_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_13_LC_18_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_13_LC_18_14_3  (
            .in0(N__44493),
            .in1(N__44534),
            .in2(_gnd_net_),
            .in3(N__44522),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51441),
            .ce(N__44409),
            .sr(N__49599));
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_18_14_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_18_14_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.pulses2count_esr_8_LC_18_14_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_8_LC_18_14_5  (
            .in0(N__44516),
            .in1(_gnd_net_),
            .in2(N__44504),
            .in3(N__44420),
            .lcout(\ppm_encoder_1.pulses2countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51441),
            .ce(N__44409),
            .sr(N__49599));
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_18_15_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNISVPV2_7_LC_18_15_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.throttle_RNISVPV2_7_LC_18_15_0  (
            .in0(N__45510),
            .in1(N__45965),
            .in2(N__45934),
            .in3(N__45803),
            .lcout(),
            .ltout(\ppm_encoder_1.un2_throttle_iv_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_18_15_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.throttle_RNILVOO6_7_LC_18_15_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \ppm_encoder_1.throttle_RNILVOO6_7_LC_18_15_1  (
            .in0(N__45731),
            .in1(_gnd_net_),
            .in2(N__45710),
            .in3(N__45692),
            .lcout(\ppm_encoder_1.throttle_RNILVOO6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_18_15_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNICJ7O2_7_LC_18_15_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \ppm_encoder_1.elevator_RNICJ7O2_7_LC_18_15_2  (
            .in0(N__45570),
            .in1(N__45627),
            .in2(N__45339),
            .in3(N__45424),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_18_15_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_18_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_18_15_3  (
            .in0(N__46812),
            .in1(N__45511),
            .in2(_gnd_net_),
            .in3(N__45571),
            .lcout(),
            .ltout(\ppm_encoder_1.N_293_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_18_15_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_18_15_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_18_15_4  (
            .in0(N__46584),
            .in1(_gnd_net_),
            .in2(N__45686),
            .in3(N__45628),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_7_LC_18_15_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_7_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_7_LC_18_15_5 .LUT_INIT=16'b0011110010101010;
    LogicCell40 \ppm_encoder_1.aileron_7_LC_18_15_5  (
            .in0(N__45629),
            .in1(N__45677),
            .in2(N__45662),
            .in3(N__46155),
            .lcout(\ppm_encoder_1.aileronZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51427),
            .ce(),
            .sr(N__49605));
    defparam \ppm_encoder_1.elevator_7_LC_18_15_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_7_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_7_LC_18_15_6 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.elevator_7_LC_18_15_6  (
            .in0(N__45572),
            .in1(N__45617),
            .in2(N__46193),
            .in3(N__45605),
            .lcout(\ppm_encoder_1.elevatorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51427),
            .ce(),
            .sr(N__49605));
    defparam \ppm_encoder_1.throttle_7_LC_18_15_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_7_LC_18_15_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_7_LC_18_15_7 .LUT_INIT=16'b0101101011001100;
    LogicCell40 \ppm_encoder_1.throttle_7_LC_18_15_7  (
            .in0(N__45560),
            .in1(N__45512),
            .in2(N__45545),
            .in3(N__46156),
            .lcout(\ppm_encoder_1.throttleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51427),
            .ce(),
            .sr(N__49605));
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_18_16_0 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.elevator_RNI6D7O2_4_LC_18_16_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \ppm_encoder_1.elevator_RNI6D7O2_4_LC_18_16_0  (
            .in0(N__46677),
            .in1(N__46476),
            .in2(N__45452),
            .in3(N__45308),
            .lcout(\ppm_encoder_1.un2_throttle_iv_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.aileron_4_LC_18_16_1 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_4_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.aileron_4_LC_18_16_1 .LUT_INIT=16'b0011101011001010;
    LogicCell40 \ppm_encoder_1.aileron_4_LC_18_16_1  (
            .in0(N__46478),
            .in1(N__46880),
            .in2(N__46191),
            .in3(N__46867),
            .lcout(\ppm_encoder_1.aileronZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51413),
            .ce(),
            .sr(N__49610));
    defparam \ppm_encoder_1.elevator_4_LC_18_16_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.elevator_4_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.elevator_4_LC_18_16_2 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \ppm_encoder_1.elevator_4_LC_18_16_2  (
            .in0(N__46679),
            .in1(N__46151),
            .in2(N__46850),
            .in3(N__46835),
            .lcout(\ppm_encoder_1.elevatorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51413),
            .ce(),
            .sr(N__49610));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_18_16_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_18_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_18_16_3  (
            .in0(N__46811),
            .in1(N__46413),
            .in2(_gnd_net_),
            .in3(N__46678),
            .lcout(),
            .ltout(\ppm_encoder_1.N_290_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_18_16_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_18_16_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__46585),
            .in2(N__46481),
            .in3(N__46477),
            .lcout(\ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.throttle_4_LC_18_16_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.throttle_4_LC_18_16_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.throttle_4_LC_18_16_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \ppm_encoder_1.throttle_4_LC_18_16_5  (
            .in0(N__46457),
            .in1(N__46442),
            .in2(N__46192),
            .in3(N__46414),
            .lcout(\ppm_encoder_1.throttleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51413),
            .ce(),
            .sr(N__49610));
    defparam \ppm_encoder_1.aileron_0_LC_18_16_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.aileron_0_LC_18_16_7 .SEQ_MODE=4'b1001;
    defparam \ppm_encoder_1.aileron_0_LC_18_16_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \ppm_encoder_1.aileron_0_LC_18_16_7  (
            .in0(N__46144),
            .in1(N__46031),
            .in2(_gnd_net_),
            .in3(N__45997),
            .lcout(\ppm_encoder_1.aileronZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51413),
            .ce(),
            .sr(N__49610));
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_17_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_1_c_LC_18_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_1_c_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__45977),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_17_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_9_c_LC_18_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_9_c_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__45971),
            .in2(N__48176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_0 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_17_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_LC_18_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__47126),
            .in2(N__48104),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_1 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_17_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_21_c_LC_18_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_21_c_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__46928),
            .in2(N__48173),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_2 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_17_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_LC_18_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__47054),
            .in2(N__48105),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_3 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_17_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_LC_18_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__47093),
            .in2(N__48174),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_4 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_17_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_LC_18_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__47021),
            .in2(N__48106),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_5 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_17_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_45_c_LC_18_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_45_c_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__46919),
            .in2(N__48175),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_6 ),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_18_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_51_c_LC_18_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_51_c_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__46910),
            .in2(N__48210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_18_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_57_c_LC_18_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ppm_encoder_1.counter24_0_I_57_c_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__46898),
            .in2(N__48161),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ppm_encoder_1.counter24_0_data_tmp_8 ),
            .carryout(\ppm_encoder_1.counter24_0_N_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_18_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47177),
            .lcout(\ppm_encoder_1.counter24_0_N_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_18_18_3 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_18_18_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_18_18_3  (
            .in0(N__47319),
            .in1(N__47150),
            .in2(N__47141),
            .in3(N__47340),
            .lcout(\ppm_encoder_1.counter24_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_18_4 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_18_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_18_4  (
            .in0(N__47120),
            .in1(N__47575),
            .in2(N__47108),
            .in3(N__47197),
            .lcout(\ppm_encoder_1.counter24_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_18_18_5 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter_RNIK1KG_0_LC_18_18_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \ppm_encoder_1.counter_RNIK1KG_0_LC_18_18_5  (
            .in0(N__47222),
            .in1(N__46996),
            .in2(N__47201),
            .in3(N__47576),
            .lcout(\ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_18_18_6 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_18_18_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_18_18_6  (
            .in0(N__47078),
            .in1(N__47221),
            .in2(N__47069),
            .in3(N__47246),
            .lcout(\ppm_encoder_1.counter24_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_18_7 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_18_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_18_7  (
            .in0(N__47525),
            .in1(N__47048),
            .in2(N__47036),
            .in3(N__47549),
            .lcout(\ppm_encoder_1.counter24_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ppm_encoder_1.counter_0_LC_18_19_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_0_LC_18_19_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_0_LC_18_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_0_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__46997),
            .in2(N__47014),
            .in3(N__47015),
            .lcout(\ppm_encoder_1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_1_LC_18_19_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_1_LC_18_19_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_1_LC_18_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_1_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__46979),
            .in2(_gnd_net_),
            .in3(N__46961),
            .lcout(\ppm_encoder_1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_0 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_2_LC_18_19_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_2_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_2_LC_18_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_2_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__46953),
            .in2(_gnd_net_),
            .in3(N__47369),
            .lcout(\ppm_encoder_1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_1 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_3_LC_18_19_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_3_LC_18_19_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_3_LC_18_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_3_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__47366),
            .in2(_gnd_net_),
            .in3(N__47345),
            .lcout(\ppm_encoder_1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_2 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_4_LC_18_19_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_4_LC_18_19_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_4_LC_18_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_4_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__47342),
            .in2(_gnd_net_),
            .in3(N__47324),
            .lcout(\ppm_encoder_1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_3 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_5_LC_18_19_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_5_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_5_LC_18_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_5_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__47321),
            .in2(_gnd_net_),
            .in3(N__47303),
            .lcout(\ppm_encoder_1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_4 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_6_LC_18_19_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_6_LC_18_19_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_6_LC_18_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_6_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__47299),
            .in2(_gnd_net_),
            .in3(N__47279),
            .lcout(\ppm_encoder_1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_5 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_7_LC_18_19_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_7_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_7_LC_18_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_7_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__47271),
            .in2(_gnd_net_),
            .in3(N__47249),
            .lcout(\ppm_encoder_1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_6 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_7 ),
            .clk(N__51373),
            .ce(),
            .sr(N__47714));
    defparam \ppm_encoder_1.counter_8_LC_18_20_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_8_LC_18_20_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_8_LC_18_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_8_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__47245),
            .in2(_gnd_net_),
            .in3(N__47225),
            .lcout(\ppm_encoder_1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_9_LC_18_20_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_9_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_9_LC_18_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_9_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__47220),
            .in2(_gnd_net_),
            .in3(N__47204),
            .lcout(\ppm_encoder_1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_8 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_10_LC_18_20_2 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_10_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_10_LC_18_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_10_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__47196),
            .in2(_gnd_net_),
            .in3(N__47180),
            .lcout(\ppm_encoder_1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_9 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_11_LC_18_20_3 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_11_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_11_LC_18_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_11_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__47574),
            .in2(_gnd_net_),
            .in3(N__47552),
            .lcout(\ppm_encoder_1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_10 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_12_LC_18_20_4 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_12_LC_18_20_4 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_12_LC_18_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_12_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__47548),
            .in2(_gnd_net_),
            .in3(N__47528),
            .lcout(\ppm_encoder_1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_11 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_13_LC_18_20_5 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_13_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_13_LC_18_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_13_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__47524),
            .in2(_gnd_net_),
            .in3(N__47504),
            .lcout(\ppm_encoder_1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_12 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_14_LC_18_20_6 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_14_LC_18_20_6 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_14_LC_18_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_14_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__47497),
            .in2(_gnd_net_),
            .in3(N__47477),
            .lcout(\ppm_encoder_1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_13 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_15_LC_18_20_7 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_15_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_15_LC_18_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_15_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__47467),
            .in2(_gnd_net_),
            .in3(N__47447),
            .lcout(\ppm_encoder_1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_14 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_15 ),
            .clk(N__51360),
            .ce(),
            .sr(N__47713));
    defparam \ppm_encoder_1.counter_16_LC_18_21_0 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_16_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_16_LC_18_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_16_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__47443),
            .in2(_gnd_net_),
            .in3(N__47423),
            .lcout(\ppm_encoder_1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .clk(N__51350),
            .ce(),
            .sr(N__47712));
    defparam \ppm_encoder_1.counter_17_LC_18_21_1 .C_ON=1'b1;
    defparam \ppm_encoder_1.counter_17_LC_18_21_1 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_17_LC_18_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ppm_encoder_1.counter_17_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__47419),
            .in2(_gnd_net_),
            .in3(N__47399),
            .lcout(\ppm_encoder_1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\ppm_encoder_1.un1_counter_13_cry_16 ),
            .carryout(\ppm_encoder_1.un1_counter_13_cry_17 ),
            .clk(N__51350),
            .ce(),
            .sr(N__47712));
    defparam \ppm_encoder_1.counter_18_LC_18_21_2 .C_ON=1'b0;
    defparam \ppm_encoder_1.counter_18_LC_18_21_2 .SEQ_MODE=4'b1000;
    defparam \ppm_encoder_1.counter_18_LC_18_21_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ppm_encoder_1.counter_18_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__47391),
            .in2(_gnd_net_),
            .in3(N__47396),
            .lcout(\ppm_encoder_1.counterZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51350),
            .ce(),
            .sr(N__47712));
    defparam \pid_front.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_18_22_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_18_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pid_front.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__48784),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_18_22_1 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_18_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__48710),
            .in2(_gnd_net_),
            .in3(N__47684),
            .lcout(\pid_front.un1_pid_prereg_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_1 ),
            .carryout(\pid_front.un1_pid_prereg_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_18_22_2 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_18_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__50377),
            .in2(_gnd_net_),
            .in3(N__47666),
            .lcout(\pid_front.un1_pid_prereg_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_2 ),
            .carryout(\pid_front.un1_pid_prereg_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_18_22_3 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_18_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__48625),
            .in2(_gnd_net_),
            .in3(N__47648),
            .lcout(\pid_front.un1_pid_prereg_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_3 ),
            .carryout(\pid_front.un1_pid_prereg_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_18_22_4 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_18_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(N__48667),
            .in2(N__48207),
            .in3(N__47630),
            .lcout(\pid_front.un1_pid_prereg_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_4 ),
            .carryout(\pid_front.un1_pid_prereg_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_18_22_5 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_18_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(N__48165),
            .in2(N__50311),
            .in3(N__47615),
            .lcout(\pid_front.un1_pid_prereg_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_5 ),
            .carryout(\pid_front.un1_pid_prereg_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_18_22_6 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_18_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(N__48169),
            .in2(N__50416),
            .in3(N__47603),
            .lcout(\pid_front.un1_pid_prereg_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_6 ),
            .carryout(\pid_front.un1_pid_prereg_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_18_22_7 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_18_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(N__50491),
            .in2(N__48209),
            .in3(N__47594),
            .lcout(\pid_front.un1_pid_prereg_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_7 ),
            .carryout(\pid_front.un1_pid_prereg_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_18_23_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_18_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__48739),
            .in2(N__48208),
            .in3(N__47579),
            .lcout(\pid_front.un1_pid_prereg_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_18_23_1 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_18_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__50452),
            .in2(N__48232),
            .in3(N__48254),
            .lcout(\pid_front.un1_pid_prereg_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_9 ),
            .carryout(\pid_front.un1_pid_prereg_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_18_23_2 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_18_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__51796),
            .in2(_gnd_net_),
            .in3(N__48239),
            .lcout(\pid_front.un1_pid_prereg_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_10 ),
            .carryout(\pid_front.un1_pid_prereg_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_18_23_3 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_18_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__51760),
            .in2(N__48231),
            .in3(N__47786),
            .lcout(\pid_front.un1_pid_prereg_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_11 ),
            .carryout(\pid_front.un1_pid_prereg_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_18_23_4 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_18_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__51856),
            .in2(_gnd_net_),
            .in3(N__47771),
            .lcout(\pid_front.un1_pid_prereg_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_12 ),
            .carryout(\pid_front.un1_pid_prereg_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_18_23_5 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_18_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__50539),
            .in2(_gnd_net_),
            .in3(N__47756),
            .lcout(\pid_front.un1_pid_prereg_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_13 ),
            .carryout(\pid_front.un1_pid_prereg_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_18_23_6 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_18_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__51823),
            .in2(_gnd_net_),
            .in3(N__47744),
            .lcout(\pid_front.un1_pid_prereg_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_14 ),
            .carryout(\pid_front.un1_pid_prereg_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_18_23_7 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_18_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__50341),
            .in2(_gnd_net_),
            .in3(N__47732),
            .lcout(\pid_front.un1_pid_prereg_cry_15_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_15 ),
            .carryout(\pid_front.un1_pid_prereg_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_18_24_0 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_18_24_0 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_18_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_18_24_0  (
            .in0(_gnd_net_),
            .in1(N__51562),
            .in2(_gnd_net_),
            .in3(N__47717),
            .lcout(\pid_front.un1_pid_prereg_cry_16_THRU_CO ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\pid_front.un1_pid_prereg_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_18_24_1 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_18_24_1 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_18_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(N__50251),
            .in2(_gnd_net_),
            .in3(N__48578),
            .lcout(\pid_front.un1_pid_prereg_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_17 ),
            .carryout(\pid_front.un1_pid_prereg_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_18_24_2 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_18_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_18_24_2  (
            .in0(_gnd_net_),
            .in1(N__51907),
            .in2(_gnd_net_),
            .in3(N__48563),
            .lcout(\pid_front.un1_pid_prereg_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_18 ),
            .carryout(\pid_front.un1_pid_prereg_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_18_24_3 .C_ON=1'b1;
    defparam \pid_front.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_18_24_3 .SEQ_MODE=4'b0000;
    defparam \pid_front.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_18_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pid_front.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_18_24_3  (
            .in0(_gnd_net_),
            .in1(N__51711),
            .in2(_gnd_net_),
            .in3(N__48548),
            .lcout(\pid_front.un1_pid_prereg_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\pid_front.un1_pid_prereg_cry_19 ),
            .carryout(\pid_front.un1_pid_prereg_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.pid_prereg_esr_21_LC_18_24_4 .C_ON=1'b0;
    defparam \pid_front.pid_prereg_esr_21_LC_18_24_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.pid_prereg_esr_21_LC_18_24_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pid_front.pid_prereg_esr_21_LC_18_24_4  (
            .in0(N__51712),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48545),
            .lcout(\pid_front.pid_preregZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51328),
            .ce(N__48482),
            .sr(N__49627));
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_18_25_0 .C_ON=1'b0;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_18_25_0 .SEQ_MODE=4'b1000;
    defparam \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_18_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_18_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48455),
            .lcout(drone_H_disp_front_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51321),
            .ce(N__48359),
            .sr(N__49628));
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.C_ON=1'b0;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49746),
            .lcout(GB_BUFFER_reset_system_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_side.error_p_reg_0_LC_20_15_5 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_0_LC_20_15_5 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_0_LC_20_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_side.error_p_reg_0_LC_20_15_5  (
            .in0(N__48289),
            .in1(N__48308),
            .in2(_gnd_net_),
            .in3(N__50178),
            .lcout(\pid_side.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51460),
            .ce(),
            .sr(N__50697));
    defparam \pid_side.error_p_reg_1_LC_20_15_6 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_1_LC_20_15_6 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_1_LC_20_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_1_LC_20_15_6  (
            .in0(N__50177),
            .in1(N__49854),
            .in2(_gnd_net_),
            .in3(N__48278),
            .lcout(\pid_side.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51460),
            .ce(),
            .sr(N__50697));
    defparam \pid_side.error_p_reg_3_LC_20_15_7 .C_ON=1'b0;
    defparam \pid_side.error_p_reg_3_LC_20_15_7 .SEQ_MODE=4'b1000;
    defparam \pid_side.error_p_reg_3_LC_20_15_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_side.error_p_reg_3_LC_20_15_7  (
            .in0(N__50179),
            .in1(N__50095),
            .in2(_gnd_net_),
            .in3(N__50126),
            .lcout(\pid_side.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51460),
            .ce(),
            .sr(N__50697));
    defparam \pid_front.error_p_reg_0_LC_20_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_0_LC_20_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_0_LC_20_23_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_0_LC_20_23_0  (
            .in0(N__51658),
            .in1(N__50059),
            .in2(_gnd_net_),
            .in3(N__50081),
            .lcout(\pid_front.error_p_regZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51351),
            .ce(),
            .sr(N__50690));
    defparam \pid_side.pid_prereg_1_LC_21_19_0 .C_ON=1'b0;
    defparam \pid_side.pid_prereg_1_LC_21_19_0 .SEQ_MODE=4'b1000;
    defparam \pid_side.pid_prereg_1_LC_21_19_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \pid_side.pid_prereg_1_LC_21_19_0  (
            .in0(N__50048),
            .in1(N__49867),
            .in2(_gnd_net_),
            .in3(N__49821),
            .lcout(\pid_side.pid_preregZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51415),
            .ce(),
            .sr(N__49626));
    defparam \pid_front.state_RNIVIRQ_1_LC_21_20_2 .C_ON=1'b0;
    defparam \pid_front.state_RNIVIRQ_1_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \pid_front.state_RNIVIRQ_1_LC_21_20_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \pid_front.state_RNIVIRQ_1_LC_21_20_2  (
            .in0(_gnd_net_),
            .in1(N__49064),
            .in2(_gnd_net_),
            .in3(N__49046),
            .lcout(\pid_front.state_RNIVIRQZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pid_front.error_p_reg_1_LC_21_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_1_LC_21_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_1_LC_21_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_1_LC_21_23_6  (
            .in0(N__51657),
            .in1(N__48774),
            .in2(_gnd_net_),
            .in3(N__48794),
            .lcout(\pid_front.error_p_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51361),
            .ce(),
            .sr(N__50691));
    defparam \pid_front.error_p_reg_9_LC_22_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_9_LC_22_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_9_LC_22_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_9_LC_22_23_1  (
            .in0(N__51660),
            .in1(N__48738),
            .in2(_gnd_net_),
            .in3(N__48755),
            .lcout(\pid_front.error_p_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51375),
            .ce(),
            .sr(N__50692));
    defparam \pid_front.error_p_reg_2_LC_22_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_2_LC_22_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_2_LC_22_23_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_2_LC_22_23_7  (
            .in0(N__51659),
            .in1(N__48702),
            .in2(_gnd_net_),
            .in3(N__48719),
            .lcout(\pid_front.error_p_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51375),
            .ce(),
            .sr(N__50692));
    defparam \pid_front.error_p_reg_5_LC_23_23_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_5_LC_23_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_5_LC_23_23_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \pid_front.error_p_reg_5_LC_23_23_3  (
            .in0(N__48660),
            .in1(_gnd_net_),
            .in2(N__51680),
            .in3(N__48683),
            .lcout(\pid_front.error_p_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51386),
            .ce(),
            .sr(N__50693));
    defparam \pid_front.error_p_reg_4_LC_23_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_4_LC_23_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_4_LC_23_23_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_p_reg_4_LC_23_23_4  (
            .in0(N__48612),
            .in1(N__51671),
            .in2(_gnd_net_),
            .in3(N__48638),
            .lcout(\pid_front.error_p_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51386),
            .ce(),
            .sr(N__50693));
    defparam \pid_front.error_p_reg_14_LC_24_22_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_14_LC_24_22_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_14_LC_24_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_front.error_p_reg_14_LC_24_22_0  (
            .in0(N__50552),
            .in1(N__51665),
            .in2(_gnd_net_),
            .in3(N__50523),
            .lcout(\pid_front.error_p_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51416),
            .ce(),
            .sr(N__50696));
    defparam \pid_front.error_p_reg_8_LC_24_22_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_8_LC_24_22_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_8_LC_24_22_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_8_LC_24_22_1  (
            .in0(N__51663),
            .in1(N__50484),
            .in2(_gnd_net_),
            .in3(N__50504),
            .lcout(\pid_front.error_p_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51416),
            .ce(),
            .sr(N__50696));
    defparam \pid_front.error_p_reg_10_LC_24_22_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_10_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_10_LC_24_22_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_front.error_p_reg_10_LC_24_22_2  (
            .in0(N__50468),
            .in1(N__51664),
            .in2(_gnd_net_),
            .in3(N__50445),
            .lcout(\pid_front.error_p_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51416),
            .ce(),
            .sr(N__50696));
    defparam \pid_front.error_p_reg_7_LC_24_22_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_7_LC_24_22_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_7_LC_24_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_7_LC_24_22_3  (
            .in0(N__51662),
            .in1(N__50409),
            .in2(_gnd_net_),
            .in3(N__50426),
            .lcout(\pid_front.error_p_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51416),
            .ce(),
            .sr(N__50696));
    defparam \pid_front.error_p_reg_3_LC_24_22_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_3_LC_24_22_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_3_LC_24_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_3_LC_24_22_7  (
            .in0(N__51661),
            .in1(N__50373),
            .in2(_gnd_net_),
            .in3(N__50390),
            .lcout(\pid_front.error_p_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51416),
            .ce(),
            .sr(N__50696));
    defparam \pid_front.error_p_reg_16_LC_24_23_0 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_16_LC_24_23_0 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_16_LC_24_23_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_16_LC_24_23_0  (
            .in0(N__51668),
            .in1(N__50334),
            .in2(_gnd_net_),
            .in3(N__50354),
            .lcout(\pid_front.error_p_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_6_LC_24_23_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_6_LC_24_23_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_6_LC_24_23_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_p_reg_6_LC_24_23_1  (
            .in0(N__50292),
            .in1(N__51670),
            .in2(_gnd_net_),
            .in3(N__50318),
            .lcout(\pid_front.error_p_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_18_LC_24_23_2 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_18_LC_24_23_2 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_18_LC_24_23_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \pid_front.error_p_reg_18_LC_24_23_2  (
            .in0(N__50273),
            .in1(N__51676),
            .in2(_gnd_net_),
            .in3(N__50244),
            .lcout(\pid_front.error_p_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_19_LC_24_23_3 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_19_LC_24_23_3 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_19_LC_24_23_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_p_reg_19_LC_24_23_3  (
            .in0(N__51891),
            .in1(N__51669),
            .in2(_gnd_net_),
            .in3(N__51920),
            .lcout(\pid_front.error_p_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_13_LC_24_23_4 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_13_LC_24_23_4 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_13_LC_24_23_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_13_LC_24_23_4  (
            .in0(N__51667),
            .in1(N__51855),
            .in2(_gnd_net_),
            .in3(N__51872),
            .lcout(\pid_front.error_p_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_15_LC_24_23_5 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_15_LC_24_23_5 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_15_LC_24_23_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_15_LC_24_23_5  (
            .in0(N__51675),
            .in1(N__51822),
            .in2(_gnd_net_),
            .in3(N__51836),
            .lcout(\pid_front.error_p_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_11_LC_24_23_6 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_11_LC_24_23_6 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_11_LC_24_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \pid_front.error_p_reg_11_LC_24_23_6  (
            .in0(N__51666),
            .in1(N__51795),
            .in2(_gnd_net_),
            .in3(N__51803),
            .lcout(\pid_front.error_p_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_12_LC_24_23_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_12_LC_24_23_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_12_LC_24_23_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pid_front.error_p_reg_12_LC_24_23_7  (
            .in0(N__51677),
            .in1(N__51776),
            .in2(_gnd_net_),
            .in3(N__51750),
            .lcout(\pid_front.error_p_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51401),
            .ce(),
            .sr(N__50695));
    defparam \pid_front.error_p_reg_20_LC_24_24_1 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_20_LC_24_24_1 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_20_LC_24_24_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \pid_front.error_p_reg_20_LC_24_24_1  (
            .in0(N__51699),
            .in1(N__51731),
            .in2(_gnd_net_),
            .in3(N__51679),
            .lcout(\pid_front.error_p_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51387),
            .ce(),
            .sr(N__50694));
    defparam \pid_front.error_p_reg_17_LC_24_24_7 .C_ON=1'b0;
    defparam \pid_front.error_p_reg_17_LC_24_24_7 .SEQ_MODE=4'b1000;
    defparam \pid_front.error_p_reg_17_LC_24_24_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \pid_front.error_p_reg_17_LC_24_24_7  (
            .in0(N__51561),
            .in1(N__51678),
            .in2(_gnd_net_),
            .in3(N__51575),
            .lcout(\pid_front.error_p_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__51387),
            .ce(),
            .sr(N__50694));
endmodule // Pc2drone
