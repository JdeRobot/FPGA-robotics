-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Apr 22 2019 18:24:36

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_pc : in std_logic;
    debug_CH5_31B : out std_logic;
    debug_CH3_20A : out std_logic;
    debug_CH0_16A : out std_logic;
    uart_input_drone : in std_logic;
    ppm_output : out std_logic;
    debug_CH6_5B : out std_logic;
    debug_CH2_18A : out std_logic;
    debug_CH4_2A : out std_logic;
    debug_CH1_0A : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46800\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45792\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45112\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40568\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_1\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_16\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_0\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_2\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_17\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_1\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_3\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_18\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_2\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_4\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_19\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_3\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_5\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_20\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_4\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_6\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_21\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_5\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_22\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_7\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_6\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_7\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_23\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_8\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_9\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_8\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_10\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_9\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_11\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_10\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_12\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_11\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_13\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_12\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_14\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_13\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_15\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_14\ : std_logic;
signal \pid_alt.un1_error_d_reg_add_1_cry_15\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_24\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_16\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \pid_alt.O_10\ : std_logic;
signal \pid_alt.un1_error_d_reg_2_0\ : std_logic;
signal \pid_alt.un1_error_d_reg_1_15\ : std_logic;
signal \pid_alt.O_13\ : std_logic;
signal \pid_alt.O_11\ : std_logic;
signal \pid_alt.O_5\ : std_logic;
signal \pid_alt.O_14\ : std_logic;
signal \pid_alt.O_6\ : std_logic;
signal \pid_alt.O_12\ : std_logic;
signal \pid_alt.O_9\ : std_logic;
signal \pid_alt.O_7\ : std_logic;
signal \pid_alt.O_1_4\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_0\ : std_logic;
signal \pid_alt.error_filt\ : std_logic;
signal \pid_alt.O_2_5\ : std_logic;
signal \pid_alt.error_filt_0\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \pid_alt.O_3_6\ : std_logic;
signal \pid_alt.O_2_6\ : std_logic;
signal \pid_alt.error_filt_cry_0\ : std_logic;
signal \pid_alt.O_3_7\ : std_logic;
signal \pid_alt.O_2_7\ : std_logic;
signal \pid_alt.error_filt_cry_1\ : std_logic;
signal \pid_alt.O_3_8\ : std_logic;
signal \pid_alt.O_2_8\ : std_logic;
signal \pid_alt.error_filt_cry_2\ : std_logic;
signal \pid_alt.O_3_9\ : std_logic;
signal \pid_alt.O_2_9\ : std_logic;
signal \pid_alt.error_filt_cry_3\ : std_logic;
signal \pid_alt.O_2_10\ : std_logic;
signal \pid_alt.O_3_10\ : std_logic;
signal \pid_alt.error_filt_cry_4\ : std_logic;
signal \pid_alt.O_3_11\ : std_logic;
signal \pid_alt.O_2_11\ : std_logic;
signal \pid_alt.error_filt_cry_5\ : std_logic;
signal \pid_alt.O_2_12\ : std_logic;
signal \pid_alt.O_3_12\ : std_logic;
signal \pid_alt.error_filt_cry_6\ : std_logic;
signal \pid_alt.error_filt_cry_7\ : std_logic;
signal \pid_alt.O_3_13\ : std_logic;
signal \pid_alt.O_2_13\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal \pid_alt.O_3_14\ : std_logic;
signal \pid_alt.O_2_14\ : std_logic;
signal \pid_alt.error_filt_cry_8\ : std_logic;
signal \pid_alt.O_1_15\ : std_logic;
signal \pid_alt.error_filt_cry_9\ : std_logic;
signal \pid_alt.O_1_16\ : std_logic;
signal \pid_alt.error_filt_cry_10\ : std_logic;
signal \pid_alt.O_1_17\ : std_logic;
signal \pid_alt.error_filt_cry_11\ : std_logic;
signal \pid_alt.O_1_18\ : std_logic;
signal \pid_alt.error_filt_cry_12\ : std_logic;
signal \pid_alt.O_1_19\ : std_logic;
signal \pid_alt.error_filt_cry_13\ : std_logic;
signal \pid_alt.O_1_20\ : std_logic;
signal \pid_alt.error_filt_cry_14\ : std_logic;
signal \pid_alt.error_filt_cry_15\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \pid_alt.error_filt_cry_16\ : std_logic;
signal \pid_alt.error_filt_cry_17\ : std_logic;
signal \pid_alt.error_filt_cry_18\ : std_logic;
signal \pid_alt.error_filt_cry_19\ : std_logic;
signal \pid_alt.error_filt_cry_20\ : std_logic;
signal \pid_alt.O_1_21\ : std_logic;
signal \pid_alt.error_filt_cry_21\ : std_logic;
signal \pid_alt.O_1_11\ : std_logic;
signal \pid_alt.O_1_12\ : std_logic;
signal \pid_alt.O_1_10\ : std_logic;
signal \pid_alt.O_0_17\ : std_logic;
signal \pid_alt.O_0_20\ : std_logic;
signal \pid_alt.O_0_23\ : std_logic;
signal \pid_alt.O_1_13\ : std_logic;
signal \pid_alt.O_0_21\ : std_logic;
signal \pid_alt.O_0_24\ : std_logic;
signal \pid_alt.O_0_18\ : std_logic;
signal \pid_alt.O_0_19\ : std_logic;
signal \pid_alt.error_p_regZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_17\ : std_logic;
signal \pid_alt.error_d_regZ0Z_17\ : std_logic;
signal alt_kd_2 : std_logic;
signal alt_kd_3 : std_logic;
signal alt_kd_7 : std_logic;
signal alt_kd_1 : std_logic;
signal alt_kd_0 : std_logic;
signal \pid_alt.g0_0_0_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_19\ : std_logic;
signal \pid_alt.error_p_regZ0Z_19\ : std_logic;
signal \pid_alt.O_1_6\ : std_logic;
signal \pid_alt.O_1_5\ : std_logic;
signal \pid_alt.O_1_14\ : std_logic;
signal alt_kp_3 : std_logic;
signal alt_kp_1 : std_logic;
signal alt_kp_7 : std_logic;
signal alt_kp_2 : std_logic;
signal \pid_alt.O_0_22\ : std_logic;
signal alt_kd_6 : std_logic;
signal alt_kd_5 : std_logic;
signal \pid_alt.O_4\ : std_logic;
signal \pid_alt.N_1074_0\ : std_logic;
signal \pid_alt.N_5_0\ : std_logic;
signal \pid_alt.g1_1\ : std_logic;
signal \pid_alt.N_1080_0_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_fastZ0Z_1\ : std_logic;
signal \pid_alt.N_3_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0\ : std_logic;
signal \pid_alt.N_1078_0\ : std_logic;
signal \pid_alt.error_p_regZ0Z_1\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_1\ : std_logic;
signal \pid_alt.error_d_regZ0Z_1\ : std_logic;
signal \pid_alt.N_1074_1\ : std_logic;
signal \pid_alt.N_3_1_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2\ : std_logic;
signal \pid_alt.g1_0\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_20\ : std_logic;
signal \pid_alt.error_d_regZ0Z_20\ : std_logic;
signal \pid_alt.O_1_7\ : std_logic;
signal alt_kp_0 : std_logic;
signal alt_kp_6 : std_logic;
signal alt_kp_5 : std_logic;
signal \pid_alt.O_0_16\ : std_logic;
signal alt_kd_4 : std_logic;
signal \Commands_frame_decoder.source_alt_kd_1_sqmuxa\ : std_logic;
signal \pid_alt.g0_4_0\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_2\ : std_logic;
signal \pid_alt.error_p_regZ0Z_2\ : std_logic;
signal \pid_alt.error_d_regZ0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2\ : std_logic;
signal \pid_alt.error_p_regZ0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_3\ : std_logic;
signal \pid_alt.error_d_regZ0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\ : std_logic;
signal \pid_alt.error_p_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_12\ : std_logic;
signal \pid_alt.error_d_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_13\ : std_logic;
signal \pid_alt.O_0_15\ : std_logic;
signal \dron_frame_decoder_1.WDT10lto9_3_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt12_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i_1\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt12_0\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0\ : std_logic;
signal \pid_alt.state_1_0_0\ : std_logic;
signal \pid_alt.error_p_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_11\ : std_logic;
signal \pid_alt.error_d_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_16\ : std_logic;
signal \pid_alt.error_d_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_7\ : std_logic;
signal \pid_alt.error_d_regZ0Z_7\ : std_logic;
signal \pid_alt.error_p_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_0\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_15\ : std_logic;
signal \pid_alt.error_d_regZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\ : std_logic;
signal \pid_alt.error_p_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_22\ : std_logic;
signal \pid_alt.error_d_regZ0Z_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_23\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_23\ : std_logic;
signal \pid_alt.O_1_8\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_8\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_11\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_12\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_14\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.N_188_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_188_4\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_1\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1\ : std_logic;
signal \pid_alt.error_p_regZ0Z_0\ : std_logic;
signal \pid_alt.error_d_regZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.state_RNO_1Z0Z_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_i_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\ : std_logic;
signal \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_4\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_5\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_6\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_7\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_8\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\ : std_logic;
signal \pid_alt.pid_preregZ0Z_16\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\ : std_logic;
signal \pid_alt.pid_preregZ0Z_17\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\ : std_logic;
signal \pid_alt.pid_preregZ0Z_18\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\ : std_logic;
signal \pid_alt.pid_preregZ0Z_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_20\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_21\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_23\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_24\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_25\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_26\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_27\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_28\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_29\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26\ : std_logic;
signal \pid_alt.un1_pid_prereg_296_1_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26\ : std_logic;
signal \pid_alt.error_d_regZ0Z_27\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_27\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \pid_alt.error_1\ : std_logic;
signal \pid_alt.error_cry_0\ : std_logic;
signal \pid_alt.error_2\ : std_logic;
signal \pid_alt.error_cry_1\ : std_logic;
signal \pid_alt.error_3\ : std_logic;
signal \pid_alt.error_cry_2\ : std_logic;
signal \pid_alt.error_4\ : std_logic;
signal \pid_alt.error_cry_3\ : std_logic;
signal alt_command_1 : std_logic;
signal \pid_alt.error_5\ : std_logic;
signal \pid_alt.error_cry_4\ : std_logic;
signal alt_command_2 : std_logic;
signal \pid_alt.error_6\ : std_logic;
signal \pid_alt.error_cry_5\ : std_logic;
signal alt_command_3 : std_logic;
signal \pid_alt.error_7\ : std_logic;
signal \pid_alt.error_cry_6\ : std_logic;
signal \pid_alt.error_cry_7\ : std_logic;
signal \pid_alt.error_8\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \pid_alt.error_9\ : std_logic;
signal \pid_alt.error_cry_8\ : std_logic;
signal \pid_alt.error_10\ : std_logic;
signal \pid_alt.error_cry_9\ : std_logic;
signal \pid_alt.error_11\ : std_logic;
signal \pid_alt.error_cry_10\ : std_logic;
signal \pid_alt.error_12\ : std_logic;
signal \pid_alt.error_cry_11\ : std_logic;
signal \pid_alt.error_13\ : std_logic;
signal \pid_alt.error_cry_12\ : std_logic;
signal \pid_alt.error_14\ : std_logic;
signal \pid_alt.error_cry_13\ : std_logic;
signal \pid_alt.error_cry_14\ : std_logic;
signal \pid_alt.error_15\ : std_logic;
signal alt_command_4 : std_logic;
signal alt_command_5 : std_logic;
signal alt_command_6 : std_logic;
signal alt_command_7 : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27\ : std_logic;
signal \pid_alt.un1_pid_prereg_296_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27\ : std_logic;
signal \pid_alt.N_410_0\ : std_logic;
signal \uart_drone_sync.aux_1__0__0_0\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0__0_0\ : std_logic;
signal \Commands_frame_decoder.WDT8lto13_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.WDT8lto9_3_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT8lt12_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxacf1\ : std_logic;
signal \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\ : std_logic;
signal \uart_drone_sync.aux_2__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_3__0__0_0\ : std_logic;
signal \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_322_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_RNIF38SZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.N_354\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_8\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_7\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \pid_alt.un9lto29_i_a2\ : std_logic;
signal \pid_alt.un9lto29_i_a2_0\ : std_logic;
signal \pid_alt.un9lto29_i_a2_1\ : std_logic;
signal \pid_alt.un9lto29_i_a2_2\ : std_logic;
signal \pid_alt.un9lto29_i_a2_3\ : std_logic;
signal \pid_alt.un9lto29_i_a2_4\ : std_logic;
signal \pid_alt.N_232_i\ : std_logic;
signal \pid_alt.un9lto29_i_a2_5\ : std_logic;
signal \pid_alt.un9lto29_i_a2_6\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_22\ : std_logic;
signal \pid_alt.pid_preregZ0Z_21\ : std_logic;
signal \pid_alt.pid_preregZ0Z_23\ : std_logic;
signal \pid_alt.pid_preregZ0Z_20\ : std_logic;
signal \pid_alt.source_pid10lt4_0\ : std_logic;
signal \pid_alt.un9lto29_i_a2_2_and\ : std_logic;
signal \pid_alt.pid_preregZ0Z_28\ : std_logic;
signal \pid_alt.pid_preregZ0Z_15\ : std_logic;
signal \pid_alt.pid_preregZ0Z_29\ : std_logic;
signal \pid_alt.pid_preregZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\ : std_logic;
signal \pid_alt.error_p_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_10\ : std_logic;
signal \pid_alt.error_d_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\ : std_logic;
signal \pid_alt.error_p_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_9\ : std_logic;
signal \pid_alt.error_d_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\ : std_logic;
signal \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_26\ : std_logic;
signal \pid_alt.error_d_regZ0Z_26\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_21\ : std_logic;
signal \pid_alt.error_d_regZ0Z_21\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20\ : std_logic;
signal \pid_alt.drone_altitude_i_0\ : std_logic;
signal \pid_alt.error_axbZ0Z_3\ : std_logic;
signal drone_altitude_i_10 : std_logic;
signal drone_altitude_i_11 : std_logic;
signal \pid_alt.error_axbZ0Z_1\ : std_logic;
signal \pid_alt.error_axbZ0Z_12\ : std_logic;
signal \pid_alt.error_axbZ0Z_13\ : std_logic;
signal \pid_alt.error_axbZ0Z_14\ : std_logic;
signal \pid_alt.error_axbZ0Z_2\ : std_logic;
signal alt_ki_0 : std_logic;
signal drone_altitude_i_9 : std_logic;
signal alt_command_0 : std_logic;
signal \pid_alt.O_1_9\ : std_logic;
signal uart_input_pc_c : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \Commands_frame_decoder.N_327\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0\ : std_logic;
signal \Commands_frame_decoder.N_358_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \pid_alt.un9lto29_i_a2_3_and\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_0\ : std_logic;
signal \pid_alt.un9lto29_i_a2_4_and\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_5\ : std_logic;
signal \pid_alt.N_123_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_12\ : std_logic;
signal \pid_alt.N_123\ : std_logic;
signal \pid_alt.N_106_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0\ : std_logic;
signal \pid_alt.N_100\ : std_logic;
signal \pid_alt.N_91_1_cascade_\ : std_logic;
signal \pid_alt.un1_reset_0_i_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_26\ : std_logic;
signal \pid_alt.pid_preregZ0Z_25\ : std_logic;
signal \pid_alt.pid_preregZ0Z_27\ : std_logic;
signal \pid_alt.pid_preregZ0Z_24\ : std_logic;
signal \pid_alt.un9lto29_i_a2_5_and\ : std_logic;
signal \pid_alt.pid_preregZ0Z_13\ : std_logic;
signal \pid_alt.N_124\ : std_logic;
signal \pid_alt.pid_preregZ0Z_8\ : std_logic;
signal \pid_alt.N_12_i\ : std_logic;
signal \pid_alt.un9lto29_i_a2_0_and\ : std_logic;
signal \pid_alt.N_96\ : std_logic;
signal \pid_alt.pid_preregZ0Z_5\ : std_logic;
signal \pid_alt.pid_preregZ0Z_4\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_4\ : std_logic;
signal \pid_alt.state_RNIFCSD1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\ : std_logic;
signal \pid_alt.error_p_regZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_25\ : std_logic;
signal \pid_alt.error_d_regZ0Z_25\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_24\ : std_logic;
signal \pid_alt.error_d_regZ0Z_24\ : std_logic;
signal \pid_alt.error_p_regZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24\ : std_logic;
signal \pid_alt.error_p_regZ0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_6\ : std_logic;
signal \pid_alt.error_d_regZ0Z_6\ : std_logic;
signal drone_altitude_0 : std_logic;
signal drone_altitude_1 : std_logic;
signal drone_altitude_2 : std_logic;
signal drone_altitude_3 : std_logic;
signal \dron_frame_decoder_1.N_392_0\ : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.N_358\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_4\ : std_logic;
signal drone_altitude_i_4 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_5\ : std_logic;
signal drone_altitude_i_5 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_6\ : std_logic;
signal drone_altitude_i_6 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_7\ : std_logic;
signal drone_altitude_i_7 : std_logic;
signal drone_altitude_i_8 : std_logic;
signal uart_drone_data_2 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_10\ : std_logic;
signal uart_drone_data_4 : std_logic;
signal drone_altitude_12 : std_logic;
signal uart_drone_data_5 : std_logic;
signal drone_altitude_13 : std_logic;
signal uart_drone_data_6 : std_logic;
signal drone_altitude_14 : std_logic;
signal uart_drone_data_7 : std_logic;
signal drone_altitude_15 : std_logic;
signal uart_drone_data_0 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_8\ : std_logic;
signal uart_drone_data_1 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_9\ : std_logic;
signal \pid_alt.stateZ0Z_0\ : std_logic;
signal \pid_alt.state_0_0\ : std_logic;
signal \uart_pc_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.un1_state53_iZ0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxacf0\ : std_logic;
signal \Commands_frame_decoder.preinitZ0\ : std_logic;
signal \Commands_frame_decoder.count_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a4_0_1_1\ : std_logic;
signal \Commands_frame_decoder.N_320_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a4_0_3_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.N_364\ : std_logic;
signal \Commands_frame_decoder.N_360_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_359\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_0_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_6\ : std_logic;
signal alt_kp_4 : std_logic;
signal \Commands_frame_decoder.stateZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_1\ : std_logic;
signal \pid_alt.pid_preregZ0Z_2\ : std_logic;
signal \pid_alt.N_91_1\ : std_logic;
signal \pid_alt.pid_preregZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\ : std_logic;
signal \pid_alt.error_p_regZ0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_5\ : std_logic;
signal \pid_alt.error_d_regZ0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8lt7_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23\ : std_logic;
signal uart_drone_data_3 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_11\ : std_logic;
signal \dron_frame_decoder_1.N_384_0\ : std_logic;
signal \uart_pc_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4\ : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.N_330\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a4_2_0_0\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_1\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\ : std_logic;
signal \uart_drone.data_rdyc_1_0\ : std_logic;
signal \uart_pc.data_rdyc_1\ : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \frame_decoder_OFF3data_7\ : std_logic;
signal \frame_decoder_CH3data_7\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \frame_decoder_OFF3data_1\ : std_logic;
signal \frame_decoder_CH3data_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH3data_2\ : std_logic;
signal \frame_decoder_OFF3data_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH3data_3\ : std_logic;
signal \frame_decoder_OFF3data_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH3data_4\ : std_logic;
signal \frame_decoder_OFF3data_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH3data_5\ : std_logic;
signal \frame_decoder_OFF3data_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH3data_6\ : std_logic;
signal \frame_decoder_OFF3data_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7\ : std_logic;
signal \scaler_3.N_1239_i_l_ofxZ0\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8\ : std_logic;
signal \pid_alt.pid_preregZ0Z_7\ : std_logic;
signal \pid_alt.pid_preregZ0Z_11\ : std_logic;
signal \pid_alt.pid_preregZ0Z_10\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_4\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_9\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \scaler_4.N_1251_i_l_ofxZ0\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_16\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_15\ : std_logic;
signal \pid_alt.m7_e_4_cascade_\ : std_logic;
signal \pid_alt.N_238_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_18\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_19\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_14\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_17\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_20\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \uart_pc.N_126_li_cascade_\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa_cascade_\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.N_145_cascade_\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal uart_pc_data_0 : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \frame_decoder_CH2data_1\ : std_logic;
signal \frame_decoder_OFF2data_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH2data_2\ : std_logic;
signal \frame_decoder_OFF2data_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH2data_3\ : std_logic;
signal \frame_decoder_OFF2data_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH2data_4\ : std_logic;
signal \frame_decoder_OFF2data_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH2data_5\ : std_logic;
signal \frame_decoder_OFF2data_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH2data_6\ : std_logic;
signal \frame_decoder_OFF2data_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8\ : std_logic;
signal \frame_decoder_OFF2data_7\ : std_logic;
signal \frame_decoder_CH2data_7\ : std_logic;
signal \scaler_2.N_1227_i_l_ofxZ0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_30\ : std_logic;
signal \pid_alt.N_106\ : std_logic;
signal \pid_alt.pid_preregZ0Z_9\ : std_logic;
signal \pid_alt.N_96_i_1\ : std_logic;
signal \pid_alt.un1_reset_0_i\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1_c_RNO_0\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2_c_RNI780L\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_9\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNO_1\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal \pid_alt.un1_reset_1_0_i_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm7lto4\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_2\ : std_logic;
signal \pid_alt.m21_e_8\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_3\ : std_logic;
signal \pid_alt.m21_e_2\ : std_logic;
signal \pid_alt.m21_e_10_cascade_\ : std_logic;
signal \pid_alt.N_138\ : std_logic;
signal \pid_alt.m35_e_3\ : std_logic;
signal \pid_alt.N_62_mux_cascade_\ : std_logic;
signal \pid_alt.N_129\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_1\ : std_logic;
signal \pid_alt.m21_e_0_cascade_\ : std_logic;
signal \pid_alt.m21_e_9\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_8\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_10\ : std_logic;
signal \pid_alt.m35_e_2\ : std_logic;
signal \pid_alt.N_62_mux\ : std_logic;
signal \pid_alt.error_i_acumm7lto5\ : std_logic;
signal \pid_alt.error_i_acumm7lto12\ : std_logic;
signal \pid_alt.N_9_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_7\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \uart_pc.data_AuxZ1Z_0\ : std_logic;
signal \uart_pc.data_AuxZ1Z_1\ : std_logic;
signal \uart_pc.data_AuxZ1Z_2\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \frame_decoder_OFF2data_0\ : std_logic;
signal \frame_decoder_CH2data_0\ : std_logic;
signal \scaler_3.un2_source_data_0\ : std_logic;
signal \frame_decoder_OFF3data_0\ : std_logic;
signal \frame_decoder_CH3data_0\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal scaler_2_data_4 : std_logic;
signal scaler_2_data_5 : std_logic;
signal scaler_3_data_4 : std_logic;
signal scaler_3_data_5 : std_logic;
signal scaler_4_data_5 : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3\ : std_logic;
signal throttle_command_5 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal throttle_command_2 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\ : std_logic;
signal throttle_command_1 : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_6\ : std_logic;
signal uart_drone_data_rdy : std_logic;
signal \debug_CH1_0A_c\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal scaler_4_data_4 : std_logic;
signal ppm_output_c : std_logic;
signal throttle_command_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\ : std_logic;
signal throttle_command_4 : std_logic;
signal scaler_4_data_6 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal scaler_3_data_8 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal scaler_3_data_14 : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_0\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_1\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_4\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_3\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_5\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_7\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_8\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_9\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_10\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_10\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_12\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_11\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_12\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_13\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_15\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_16\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_17\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\ : std_logic;
signal \debug_CH3_20A_c\ : std_logic;
signal \debug_CH3_20A_c_0\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_pc.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.state_srsts_0_0_0\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_drone.N_126_li_cascade_\ : std_logic;
signal \debug_CH2_18A_c\ : std_logic;
signal \uart_pc.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal \uart_drone.data_rdyc_1\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal \debug_CH0_16A_c\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \uart_pc.CO0_cascade_\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_0\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.N_152_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7_cascade_\ : std_logic;
signal \ppm_encoder_1.N_299_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal scaler_3_data_7 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal throttle_command_7 : std_logic;
signal \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \scaler_2.un2_source_data_0\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_9\ : std_logic;
signal \debug_CH3_20A_c_0_g\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9\ : std_logic;
signal \ppm_encoder_1.N_301_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal scaler_3_data_9 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal throttle_command_9 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal scaler_3_data_12 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal throttle_command_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal throttle_command_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal scaler_3_data_11 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_320_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal scaler_3_data_10 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal reset_system : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.N_145\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_21\ : std_logic;
signal \pid_alt.error_i_acumm7lto13\ : std_logic;
signal \pid_alt.N_238\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_13\ : std_logic;
signal \pid_alt.N_96_i_0\ : std_logic;
signal uart_pc_data_6 : std_logic;
signal alt_ki_6 : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_6\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_6\ : std_logic;
signal \pid_alt.N_96_i\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_11\ : std_logic;
signal \pid_alt.N_128\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_11\ : std_logic;
signal \pid_alt.un1_reset_1_0_i\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_0\ : std_logic;
signal \pid_alt.state_0_g_0\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal \reset_module_System.reset6_13_cascade_\ : std_logic;
signal \reset_module_System.reset6_3\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.reset6_17\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.N_145_cascade_\ : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_304\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\ : std_logic;
signal \ppm_encoder_1.N_227_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.N_296_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6\ : std_logic;
signal \ppm_encoder_1.N_298_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal scaler_3_data_6 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\ : std_logic;
signal throttle_command_6 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal throttle_command_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13\ : std_logic;
signal scaler_3_data_13 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal throttle_command_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \ppm_encoder_1.N_305_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_303_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_319_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_302\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_145_17\ : std_logic;
signal \ppm_encoder_1.N_145_17_cascade_\ : std_logic;
signal \ppm_encoder_1.N_238\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \pid_alt.O_0_5\ : std_logic;
signal \pid_alt.error_i_regZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \ppm_encoder_1.N_297_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\ : std_logic;
signal throttle_command_3 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_3\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal scaler_2_data_6 : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal scaler_2_data_7 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal scaler_2_data_8 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal scaler_2_data_9 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal scaler_2_data_10 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal scaler_2_data_12 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal scaler_2_data_13 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal scaler_2_data_14 : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.pid_altitude_dv_0\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal scaler_2_data_11 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_1330_i\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_322_g\ : std_logic;
signal uart_pc_data_2 : std_logic;
signal alt_ki_2 : std_logic;
signal \pid_alt.O_0_6\ : std_logic;
signal \pid_alt.error_i_regZ0Z_2\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \uart_drone.un1_state_4_0_cascade_\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cascade_\ : std_logic;
signal pid_altitude_dv : std_logic;
signal throttle_command_0 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.throttle_RNIN3352Z0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIALN65Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.throttle_RNI5V123Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.throttle_RNI82223Z0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.throttle_RNIJII96Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \ppm_encoder_1.throttle_RNIONI96Z0Z_8\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNITSI96Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_306\ : std_logic;
signal \pid_alt.un9_error_filt_1_15\ : std_logic;
signal \pid_alt.un9_error_filt_2_0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_axbZ0Z_0\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \pid_alt.un9_error_filt_1_16\ : std_logic;
signal \pid_alt.un9_error_filt_2_1\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_1_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_0\ : std_logic;
signal \pid_alt.un9_error_filt_1_17\ : std_logic;
signal \pid_alt.un9_error_filt_2_2\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_2_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_1\ : std_logic;
signal \pid_alt.un9_error_filt_1_18\ : std_logic;
signal \pid_alt.un9_error_filt_2_3\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_3_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_2\ : std_logic;
signal \pid_alt.un9_error_filt_2_4\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_4_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_3\ : std_logic;
signal \pid_alt.un9_error_filt_2_5\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_5_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_4\ : std_logic;
signal \pid_alt.un9_error_filt_2_6\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_6_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_5\ : std_logic;
signal \pid_alt.un9_error_filt_2_7\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_7_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_6\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_7\ : std_logic;
signal \pid_alt.un9_error_filt_2_8\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \pid_alt.un9_error_filt_2_9\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_9_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_8\ : std_logic;
signal \pid_alt.un9_error_filt_2_10\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_10_sZ0\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_9\ : std_logic;
signal \pid_alt.un9_error_filt_1_19\ : std_logic;
signal \pid_alt.un9_error_filt_2_11\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_cry_10\ : std_logic;
signal \pid_alt.un9_error_filt_add_1_sZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_140_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_300\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_159_d\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \pid_alt.O_0_4\ : std_logic;
signal \pid_alt.error_i_regZ0Z_0\ : std_logic;
signal \pid_alt.O_0_7\ : std_logic;
signal \pid_alt.error_i_regZ0Z_3\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.N_227\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_59_d\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \ppm_encoder_1.N_1330_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \pid_alt.error_filt_21\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_21\ : std_logic;
signal uart_pc_data_5 : std_logic;
signal alt_ki_5 : std_logic;
signal reset_system_g : std_logic;
signal \GB_BUFFER_reset_system_g_THRU_CO\ : std_logic;
signal uart_pc_data_3 : std_logic;
signal alt_ki_3 : std_logic;
signal \pid_alt.O_0_8\ : std_logic;
signal \pid_alt.error_i_regZ0Z_4\ : std_logic;
signal \pid_alt.O_0_9\ : std_logic;
signal \pid_alt.error_i_regZ0Z_5\ : std_logic;
signal \pid_alt.O_0_12\ : std_logic;
signal \pid_alt.error_i_regZ0Z_8\ : std_logic;
signal uart_pc_data_4 : std_logic;
signal alt_ki_4 : std_logic;
signal uart_pc_data_1 : std_logic;
signal alt_ki_1 : std_logic;
signal \pid_alt.error_filt_19\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_19\ : std_logic;
signal uart_pc_data_7 : std_logic;
signal alt_ki_7 : std_logic;
signal \Commands_frame_decoder.state_RNIQRI31Z0Z_10\ : std_logic;
signal \pid_alt.O_0_14\ : std_logic;
signal \pid_alt.error_i_regZ0Z_10\ : std_logic;
signal \pid_alt.O_15\ : std_logic;
signal \pid_alt.error_i_regZ0Z_11\ : std_logic;
signal \pid_alt.O_16\ : std_logic;
signal \pid_alt.error_i_regZ0Z_12\ : std_logic;
signal \pid_alt.O_17\ : std_logic;
signal \pid_alt.error_i_regZ0Z_13\ : std_logic;
signal \pid_alt.error_filt_17\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_17\ : std_logic;
signal \pid_alt.error_filt_18\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_18\ : std_logic;
signal \pid_alt.error_filt_22\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_22\ : std_logic;
signal \pid_alt.error_filt_20\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_20\ : std_logic;
signal \pid_alt.error_filt_8\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_8\ : std_logic;
signal \pid_alt.O_8\ : std_logic;
signal \pid_alt.error_d_regZ0Z_4\ : std_logic;
signal \pid_alt.error_filt_1\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_1\ : std_logic;
signal \pid_alt.error_filt_2\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_2\ : std_logic;
signal \pid_alt.error_filt_10\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_10\ : std_logic;
signal \pid_alt.error_filt_11\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_11\ : std_logic;
signal \pid_alt.error_filt_12\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_12\ : std_logic;
signal \pid_alt.error_filt_13\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_13\ : std_logic;
signal \pid_alt.error_filt_15\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_15\ : std_logic;
signal \pid_alt.error_filt_16\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_16\ : std_logic;
signal \pid_alt.error_filt_4\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_4\ : std_logic;
signal \pid_alt.error_filt_5\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_5\ : std_logic;
signal \pid_alt.error_filt_6\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_6\ : std_logic;
signal \pid_alt.error_filt_7\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_7\ : std_logic;
signal \pid_alt.error_filt_9\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_9\ : std_logic;
signal \pid_alt.error_filt_3\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_3\ : std_logic;
signal \pid_alt.error_filt_14\ : std_logic;
signal \pid_alt.error_filt_prevZ0Z_14\ : std_logic;
signal \pid_alt.O_0_11\ : std_logic;
signal \pid_alt.error_i_regZ0Z_7\ : std_logic;
signal \pid_alt.O_0_10\ : std_logic;
signal \pid_alt.error_i_regZ0Z_6\ : std_logic;
signal \pid_alt.O_19\ : std_logic;
signal \pid_alt.error_i_regZ0Z_15\ : std_logic;
signal \pid_alt.O_0_13\ : std_logic;
signal \pid_alt.error_i_regZ0Z_9\ : std_logic;
signal \pid_alt.O_18\ : std_logic;
signal \pid_alt.error_i_regZ0Z_14\ : std_logic;
signal \pid_alt.O_24\ : std_logic;
signal \pid_alt.error_i_regZ0Z_20\ : std_logic;
signal \pid_alt.O_21\ : std_logic;
signal \pid_alt.error_i_regZ0Z_17\ : std_logic;
signal \pid_alt.O_22\ : std_logic;
signal \pid_alt.error_i_regZ0Z_18\ : std_logic;
signal \pid_alt.O_20\ : std_logic;
signal \pid_alt.error_i_regZ0Z_16\ : std_logic;
signal \pid_alt.O_23\ : std_logic;
signal \pid_alt.error_i_regZ0Z_19\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal \pid_alt.N_410_0_g\ : std_logic;
signal \N_411_g\ : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_drone_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal \debug_CH2_18A_wire\ : std_logic;
signal \debug_CH0_16A_wire\ : std_logic;
signal \debug_CH1_0A_wire\ : std_logic;
signal \debug_CH5_31B_wire\ : std_logic;
signal \debug_CH4_2A_wire\ : std_logic;
signal ppm_output_wire : std_logic;
signal \debug_CH3_20A_wire\ : std_logic;
signal \debug_CH6_5B_wire\ : std_logic;
signal \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un9_error_filt_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_mulonly_0_21_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_21_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_21_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_21_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_21_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un9_error_filt_2_mulonly_0_11_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_2_mulonly_0_11_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_2_mulonly_0_11_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_2_mulonly_0_11_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    clk_system_wire <= clk_system;
    uart_input_drone_wire <= uart_input_drone;
    uart_input_pc_wire <= uart_input_pc;
    debug_CH2_18A <= \debug_CH2_18A_wire\;
    debug_CH0_16A <= \debug_CH0_16A_wire\;
    debug_CH1_0A <= \debug_CH1_0A_wire\;
    debug_CH5_31B <= \debug_CH5_31B_wire\;
    debug_CH4_2A <= \debug_CH4_2A_wire\;
    ppm_output <= ppm_output_wire;
    debug_CH3_20A <= \debug_CH3_20A_wire\;
    debug_CH6_5B <= \debug_CH6_5B_wire\;
    \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__22139\&\N__22196\&\N__22243\&\N__21569\&\N__21616\&\N__21672\&\N__21716\&\N__21770\&\N__21830\&\N__21889\&\N__21953\&\N__21329\&\N__21379\&\N__21435\&\N__21485\&\N__24458\;
    \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18534\&\N__19032\&\N__19020\&\N__25506\&\N__18561\&\N__18777\&\N__18546\&\N__19047\;
    \pid_alt.O_0_24\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_0_23\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_0_22\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_0_21\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_0_20\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_0_19\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_0_18\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_0_17\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_0_16\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_0_15\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_1_14\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_1_13\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_1_12\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_1_11\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_1_10\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_1_9\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_1_8\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_1_7\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_1_6\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_1_5\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_1_4\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un9_error_filt_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un9_error_filt_1_mulonly_0_19_0_A_wire\ <= '0'&\N__46254\&\N__45996\&\N__46032\&\N__46071\&\N__46113\&\N__46320\&\N__45534\&\N__46365\&\N__46398\&\N__45837\&\N__45870\&\N__46287\&\N__46149\&\N__45429\&\N__17958\;
    \pid_alt.un9_error_filt_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un9_error_filt_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__43087\&\N__43129\&\N__43086\;
    \pid_alt.un9_error_filt_1_19\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(19);
    \pid_alt.un9_error_filt_1_18\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(18);
    \pid_alt.un9_error_filt_1_17\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(17);
    \pid_alt.un9_error_filt_1_16\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(16);
    \pid_alt.un9_error_filt_1_15\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(15);
    \pid_alt.O_3_14\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(14);
    \pid_alt.O_3_13\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(13);
    \pid_alt.O_3_12\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(12);
    \pid_alt.O_3_11\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(11);
    \pid_alt.O_3_10\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(10);
    \pid_alt.O_3_9\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(9);
    \pid_alt.O_3_8\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(8);
    \pid_alt.O_3_7\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(7);
    \pid_alt.O_3_6\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(6);
    \pid_alt.error_filt\ <= \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\(5);
    \pid_alt.un2_error_mulonly_0_21_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_21_0_A_wire\ <= \N__22132\&\N__22189\&\N__22247\&\N__21562\&\N__21620\&\N__21664\&\N__21709\&\N__21763\&\N__21820\&\N__21890\&\N__21946\&\N__21322\&\N__21383\&\N__21430\&\N__21472\&\N__24451\;
    \pid_alt.un2_error_mulonly_0_21_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_21_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__43055\&\N__43052\&'0'&'0'&\N__43054\;
    \pid_alt.O_1_21\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(21);
    \pid_alt.O_1_20\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(20);
    \pid_alt.O_1_19\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(19);
    \pid_alt.O_1_18\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(18);
    \pid_alt.O_1_17\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(17);
    \pid_alt.O_1_16\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(16);
    \pid_alt.O_1_15\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(15);
    \pid_alt.O_2_14\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(14);
    \pid_alt.O_2_13\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(13);
    \pid_alt.O_2_12\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(12);
    \pid_alt.O_2_11\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(11);
    \pid_alt.O_2_10\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(10);
    \pid_alt.O_2_9\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(9);
    \pid_alt.O_2_8\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(8);
    \pid_alt.O_2_7\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(7);
    \pid_alt.O_2_6\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(6);
    \pid_alt.O_2_5\ <= \pid_alt.un2_error_mulonly_0_21_0_O_wire\(5);
    \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_A_wire\ <= '0'&\N__46277\&\N__46019\&\N__46055\&\N__46094\&\N__46136\&\N__46343\&\N__45557\&\N__46388\&\N__46421\&\N__45860\&\N__45893\&\N__46310\&\N__46172\&\N__45452\&\N__17883\;
    \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18392\&\N__18752\&\N__18731\&\N__18992\&\N__18416\&\N__18440\&\N__18368\&\N__18341\;
    \pid_alt.un1_error_d_reg_1_24\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(24);
    \pid_alt.un1_error_d_reg_1_23\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(23);
    \pid_alt.un1_error_d_reg_1_22\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(22);
    \pid_alt.un1_error_d_reg_1_21\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(21);
    \pid_alt.un1_error_d_reg_1_20\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(20);
    \pid_alt.un1_error_d_reg_1_19\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(19);
    \pid_alt.un1_error_d_reg_1_18\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(18);
    \pid_alt.un1_error_d_reg_1_17\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(17);
    \pid_alt.un1_error_d_reg_1_16\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(16);
    \pid_alt.un1_error_d_reg_1_15\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_14\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_13\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_12\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_11\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_10\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_9\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_8\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_7\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_6\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_5\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_4\ <= \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ <= \N__22149\&\N__22206\&\N__22248\&\N__21579\&\N__21627\&\N__21668\&\N__21726\&\N__21780\&\N__21837\&\N__21891\&\N__21963\&\N__21339\&\N__21390\&\N__21434\&\N__21486\&\N__24462\;
    \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__44877\&\N__33300\&\N__44154\&\N__45237\&\N__43230\&\N__36750\&\N__45078\&\N__23391\;
    \pid_alt.O_24\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_23\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_22\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_21\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_20\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_19\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_18\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_17\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_16\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_15\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_0_14\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_0_13\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_0_12\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_0_11\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_0_10\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_0_9\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_0_8\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_0_7\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_0_6\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_0_5\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_0_4\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_A_wire\ <= \N__45692\&\N__45698\&\N__45694\&\N__45695\&\N__45693\&\N__45696\&\N__45691\&\N__45697\&\N__45690\&\N__44330\&\N__45596\&\N__45050\&\N__45734\&\N__45785\&\N__45935\&\N__45983\;
    \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18393\&\N__18753\&\N__18732\&\N__18996\&\N__18417\&\N__18441\&\N__18369\&\N__18345\;
    \pid_alt.un1_error_d_reg_2_16\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(16);
    \pid_alt.un1_error_d_reg_2_15\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(15);
    \pid_alt.un1_error_d_reg_2_14\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(14);
    \pid_alt.un1_error_d_reg_2_13\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(13);
    \pid_alt.un1_error_d_reg_2_12\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(12);
    \pid_alt.un1_error_d_reg_2_11\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(11);
    \pid_alt.un1_error_d_reg_2_10\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(10);
    \pid_alt.un1_error_d_reg_2_9\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(9);
    \pid_alt.un1_error_d_reg_2_8\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(8);
    \pid_alt.un1_error_d_reg_2_7\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(7);
    \pid_alt.un1_error_d_reg_2_6\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(6);
    \pid_alt.un1_error_d_reg_2_5\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(5);
    \pid_alt.un1_error_d_reg_2_4\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(4);
    \pid_alt.un1_error_d_reg_2_3\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(3);
    \pid_alt.un1_error_d_reg_2_2\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(2);
    \pid_alt.un1_error_d_reg_2_1\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(1);
    \pid_alt.un1_error_d_reg_2_0\ <= \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\(0);
    \pid_alt.un9_error_filt_2_mulonly_0_11_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un9_error_filt_2_mulonly_0_11_0_A_wire\ <= \N__45632\&\N__45635\&\N__45631\&\N__45636\&\N__45630\&\N__45633\&\N__45629\&\N__45634\&\N__45628\&\N__44307\&\N__45567\&\N__45027\&\N__45711\&\N__45762\&\N__45906\&\N__45954\;
    \pid_alt.un9_error_filt_2_mulonly_0_11_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un9_error_filt_2_mulonly_0_11_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__43127\&\N__43125\&\N__43126\;
    \pid_alt.un9_error_filt_2_11\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(11);
    \pid_alt.un9_error_filt_2_10\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(10);
    \pid_alt.un9_error_filt_2_9\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(9);
    \pid_alt.un9_error_filt_2_8\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(8);
    \pid_alt.un9_error_filt_2_7\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(7);
    \pid_alt.un9_error_filt_2_6\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(6);
    \pid_alt.un9_error_filt_2_5\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(5);
    \pid_alt.un9_error_filt_2_4\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(4);
    \pid_alt.un9_error_filt_2_3\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(3);
    \pid_alt.un9_error_filt_2_2\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(2);
    \pid_alt.un9_error_filt_2_1\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(1);
    \pid_alt.un9_error_filt_2_0\ <= \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\(0);

    \pid_alt.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43117\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43116\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un9_error_filt_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43130\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43085\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un9_error_filt_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un9_error_filt_1_mulonly_0_19_0_A_wire\,
            C => \pid_alt.un9_error_filt_1_mulonly_0_19_0_C_wire\,
            B => \pid_alt.un9_error_filt_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un9_error_filt_1_mulonly_0_19_0_O_wire\
        );

    \pid_alt.un2_error_mulonly_0_21_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43053\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43051\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_mulonly_0_21_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_mulonly_0_21_0_A_wire\,
            C => \pid_alt.un2_error_mulonly_0_21_0_C_wire\,
            B => \pid_alt.un2_error_mulonly_0_21_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_mulonly_0_21_0_O_wire\
        );

    \pid_alt.un1_error_d_reg_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43122\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43110\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un1_error_d_reg_1_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_2_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43131\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43138\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un1_error_d_reg_2_mulonly_0_16_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43140\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43139\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_A_wire\,
            C => \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_C_wire\,
            B => \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un1_error_d_reg_2_mulonly_0_16_0_O_wire\
        );

    \pid_alt.un9_error_filt_2_mulonly_0_11_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43128\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43124\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un9_error_filt_2_mulonly_0_11_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un9_error_filt_2_mulonly_0_11_0_A_wire\,
            C => \pid_alt.un9_error_filt_2_mulonly_0_11_0_C_wire\,
            B => \pid_alt.un9_error_filt_2_mulonly_0_11_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un9_error_filt_2_mulonly_0_11_0_O_wire\
        );

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__47734\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47736\,
            DIN => \N__47735\,
            DOUT => \N__47734\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47736\,
            PADOUT => \N__47735\,
            PADIN => \N__47734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47725\,
            DIN => \N__47724\,
            DOUT => \N__47723\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47725\,
            PADOUT => \N__47724\,
            PADIN => \N__47723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47716\,
            DIN => \N__47715\,
            DOUT => \N__47714\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47716\,
            PADOUT => \N__47715\,
            PADIN => \N__47714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH2_18A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47707\,
            DIN => \N__47706\,
            DOUT => \N__47705\,
            PACKAGEPIN => \debug_CH2_18A_wire\
        );

    \debug_CH2_18A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47707\,
            PADOUT => \N__47706\,
            PADIN => \N__47705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31229\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH0_16A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47698\,
            DIN => \N__47697\,
            DOUT => \N__47696\,
            PACKAGEPIN => \debug_CH0_16A_wire\
        );

    \debug_CH0_16A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47698\,
            PADOUT => \N__47697\,
            PADIN => \N__47696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH1_0A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47689\,
            DIN => \N__47688\,
            DOUT => \N__47687\,
            PACKAGEPIN => \debug_CH1_0A_wire\
        );

    \debug_CH1_0A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47689\,
            PADOUT => \N__47688\,
            PADIN => \N__47687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH5_31B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47680\,
            DIN => \N__47679\,
            DOUT => \N__47678\,
            PACKAGEPIN => \debug_CH5_31B_wire\
        );

    \debug_CH5_31B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47680\,
            PADOUT => \N__47679\,
            PADIN => \N__47678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH4_2A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47671\,
            DIN => \N__47670\,
            DOUT => \N__47669\,
            PACKAGEPIN => \debug_CH4_2A_wire\
        );

    \debug_CH4_2A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47671\,
            PADOUT => \N__47670\,
            PADIN => \N__47669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47662\,
            DIN => \N__47661\,
            DOUT => \N__47660\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47662\,
            PADOUT => \N__47661\,
            PADIN => \N__47660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29457\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH3_20A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47653\,
            DIN => \N__47652\,
            DOUT => \N__47651\,
            PACKAGEPIN => \debug_CH3_20A_wire\
        );

    \debug_CH3_20A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47653\,
            PADOUT => \N__47652\,
            PADIN => \N__47651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH6_5B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47644\,
            DIN => \N__47643\,
            DOUT => \N__47642\,
            PACKAGEPIN => \debug_CH6_5B_wire\
        );

    \debug_CH6_5B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47644\,
            PADOUT => \N__47643\,
            PADIN => \N__47642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11503\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47622\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__47622\,
            I => \N__47619\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__47619\,
            I => \pid_alt.O_0_13\
        );

    \I__11500\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47613\
        );

    \I__11499\ : LocalMux
    port map (
            O => \N__47613\,
            I => \N__47610\
        );

    \I__11498\ : Span12Mux_h
    port map (
            O => \N__47610\,
            I => \N__47607\
        );

    \I__11497\ : Odrv12
    port map (
            O => \N__47607\,
            I => \pid_alt.error_i_regZ0Z_9\
        );

    \I__11496\ : InMux
    port map (
            O => \N__47604\,
            I => \N__47601\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__47601\,
            I => \N__47598\
        );

    \I__11494\ : Odrv4
    port map (
            O => \N__47598\,
            I => \pid_alt.O_18\
        );

    \I__11493\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47592\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__47592\,
            I => \N__47589\
        );

    \I__11491\ : Odrv12
    port map (
            O => \N__47589\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__11490\ : InMux
    port map (
            O => \N__47586\,
            I => \N__47583\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__47583\,
            I => \N__47580\
        );

    \I__11488\ : Odrv4
    port map (
            O => \N__47580\,
            I => \pid_alt.O_24\
        );

    \I__11487\ : InMux
    port map (
            O => \N__47577\,
            I => \N__47571\
        );

    \I__11486\ : InMux
    port map (
            O => \N__47576\,
            I => \N__47571\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__47571\,
            I => \N__47568\
        );

    \I__11484\ : Span12Mux_h
    port map (
            O => \N__47568\,
            I => \N__47565\
        );

    \I__11483\ : Odrv12
    port map (
            O => \N__47565\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__11482\ : InMux
    port map (
            O => \N__47562\,
            I => \N__47559\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__47559\,
            I => \N__47556\
        );

    \I__11480\ : Odrv4
    port map (
            O => \N__47556\,
            I => \pid_alt.O_21\
        );

    \I__11479\ : InMux
    port map (
            O => \N__47553\,
            I => \N__47550\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__47550\,
            I => \N__47547\
        );

    \I__11477\ : Span12Mux_h
    port map (
            O => \N__47547\,
            I => \N__47544\
        );

    \I__11476\ : Odrv12
    port map (
            O => \N__47544\,
            I => \pid_alt.error_i_regZ0Z_17\
        );

    \I__11475\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47538\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__47538\,
            I => \N__47535\
        );

    \I__11473\ : Odrv4
    port map (
            O => \N__47535\,
            I => \pid_alt.O_22\
        );

    \I__11472\ : InMux
    port map (
            O => \N__47532\,
            I => \N__47529\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__47529\,
            I => \N__47526\
        );

    \I__11470\ : Span12Mux_h
    port map (
            O => \N__47526\,
            I => \N__47523\
        );

    \I__11469\ : Odrv12
    port map (
            O => \N__47523\,
            I => \pid_alt.error_i_regZ0Z_18\
        );

    \I__11468\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47517\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__47517\,
            I => \N__47514\
        );

    \I__11466\ : Odrv4
    port map (
            O => \N__47514\,
            I => \pid_alt.O_20\
        );

    \I__11465\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47508\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__47508\,
            I => \N__47505\
        );

    \I__11463\ : Odrv12
    port map (
            O => \N__47505\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__11462\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47499\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__47499\,
            I => \pid_alt.O_23\
        );

    \I__11460\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47493\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__47493\,
            I => \N__47490\
        );

    \I__11458\ : Span4Mux_h
    port map (
            O => \N__47490\,
            I => \N__47487\
        );

    \I__11457\ : Span4Mux_h
    port map (
            O => \N__47487\,
            I => \N__47484\
        );

    \I__11456\ : Span4Mux_h
    port map (
            O => \N__47484\,
            I => \N__47481\
        );

    \I__11455\ : Odrv4
    port map (
            O => \N__47481\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__11454\ : ClkMux
    port map (
            O => \N__47478\,
            I => \N__46830\
        );

    \I__11453\ : ClkMux
    port map (
            O => \N__47477\,
            I => \N__46830\
        );

    \I__11452\ : ClkMux
    port map (
            O => \N__47476\,
            I => \N__46830\
        );

    \I__11451\ : ClkMux
    port map (
            O => \N__47475\,
            I => \N__46830\
        );

    \I__11450\ : ClkMux
    port map (
            O => \N__47474\,
            I => \N__46830\
        );

    \I__11449\ : ClkMux
    port map (
            O => \N__47473\,
            I => \N__46830\
        );

    \I__11448\ : ClkMux
    port map (
            O => \N__47472\,
            I => \N__46830\
        );

    \I__11447\ : ClkMux
    port map (
            O => \N__47471\,
            I => \N__46830\
        );

    \I__11446\ : ClkMux
    port map (
            O => \N__47470\,
            I => \N__46830\
        );

    \I__11445\ : ClkMux
    port map (
            O => \N__47469\,
            I => \N__46830\
        );

    \I__11444\ : ClkMux
    port map (
            O => \N__47468\,
            I => \N__46830\
        );

    \I__11443\ : ClkMux
    port map (
            O => \N__47467\,
            I => \N__46830\
        );

    \I__11442\ : ClkMux
    port map (
            O => \N__47466\,
            I => \N__46830\
        );

    \I__11441\ : ClkMux
    port map (
            O => \N__47465\,
            I => \N__46830\
        );

    \I__11440\ : ClkMux
    port map (
            O => \N__47464\,
            I => \N__46830\
        );

    \I__11439\ : ClkMux
    port map (
            O => \N__47463\,
            I => \N__46830\
        );

    \I__11438\ : ClkMux
    port map (
            O => \N__47462\,
            I => \N__46830\
        );

    \I__11437\ : ClkMux
    port map (
            O => \N__47461\,
            I => \N__46830\
        );

    \I__11436\ : ClkMux
    port map (
            O => \N__47460\,
            I => \N__46830\
        );

    \I__11435\ : ClkMux
    port map (
            O => \N__47459\,
            I => \N__46830\
        );

    \I__11434\ : ClkMux
    port map (
            O => \N__47458\,
            I => \N__46830\
        );

    \I__11433\ : ClkMux
    port map (
            O => \N__47457\,
            I => \N__46830\
        );

    \I__11432\ : ClkMux
    port map (
            O => \N__47456\,
            I => \N__46830\
        );

    \I__11431\ : ClkMux
    port map (
            O => \N__47455\,
            I => \N__46830\
        );

    \I__11430\ : ClkMux
    port map (
            O => \N__47454\,
            I => \N__46830\
        );

    \I__11429\ : ClkMux
    port map (
            O => \N__47453\,
            I => \N__46830\
        );

    \I__11428\ : ClkMux
    port map (
            O => \N__47452\,
            I => \N__46830\
        );

    \I__11427\ : ClkMux
    port map (
            O => \N__47451\,
            I => \N__46830\
        );

    \I__11426\ : ClkMux
    port map (
            O => \N__47450\,
            I => \N__46830\
        );

    \I__11425\ : ClkMux
    port map (
            O => \N__47449\,
            I => \N__46830\
        );

    \I__11424\ : ClkMux
    port map (
            O => \N__47448\,
            I => \N__46830\
        );

    \I__11423\ : ClkMux
    port map (
            O => \N__47447\,
            I => \N__46830\
        );

    \I__11422\ : ClkMux
    port map (
            O => \N__47446\,
            I => \N__46830\
        );

    \I__11421\ : ClkMux
    port map (
            O => \N__47445\,
            I => \N__46830\
        );

    \I__11420\ : ClkMux
    port map (
            O => \N__47444\,
            I => \N__46830\
        );

    \I__11419\ : ClkMux
    port map (
            O => \N__47443\,
            I => \N__46830\
        );

    \I__11418\ : ClkMux
    port map (
            O => \N__47442\,
            I => \N__46830\
        );

    \I__11417\ : ClkMux
    port map (
            O => \N__47441\,
            I => \N__46830\
        );

    \I__11416\ : ClkMux
    port map (
            O => \N__47440\,
            I => \N__46830\
        );

    \I__11415\ : ClkMux
    port map (
            O => \N__47439\,
            I => \N__46830\
        );

    \I__11414\ : ClkMux
    port map (
            O => \N__47438\,
            I => \N__46830\
        );

    \I__11413\ : ClkMux
    port map (
            O => \N__47437\,
            I => \N__46830\
        );

    \I__11412\ : ClkMux
    port map (
            O => \N__47436\,
            I => \N__46830\
        );

    \I__11411\ : ClkMux
    port map (
            O => \N__47435\,
            I => \N__46830\
        );

    \I__11410\ : ClkMux
    port map (
            O => \N__47434\,
            I => \N__46830\
        );

    \I__11409\ : ClkMux
    port map (
            O => \N__47433\,
            I => \N__46830\
        );

    \I__11408\ : ClkMux
    port map (
            O => \N__47432\,
            I => \N__46830\
        );

    \I__11407\ : ClkMux
    port map (
            O => \N__47431\,
            I => \N__46830\
        );

    \I__11406\ : ClkMux
    port map (
            O => \N__47430\,
            I => \N__46830\
        );

    \I__11405\ : ClkMux
    port map (
            O => \N__47429\,
            I => \N__46830\
        );

    \I__11404\ : ClkMux
    port map (
            O => \N__47428\,
            I => \N__46830\
        );

    \I__11403\ : ClkMux
    port map (
            O => \N__47427\,
            I => \N__46830\
        );

    \I__11402\ : ClkMux
    port map (
            O => \N__47426\,
            I => \N__46830\
        );

    \I__11401\ : ClkMux
    port map (
            O => \N__47425\,
            I => \N__46830\
        );

    \I__11400\ : ClkMux
    port map (
            O => \N__47424\,
            I => \N__46830\
        );

    \I__11399\ : ClkMux
    port map (
            O => \N__47423\,
            I => \N__46830\
        );

    \I__11398\ : ClkMux
    port map (
            O => \N__47422\,
            I => \N__46830\
        );

    \I__11397\ : ClkMux
    port map (
            O => \N__47421\,
            I => \N__46830\
        );

    \I__11396\ : ClkMux
    port map (
            O => \N__47420\,
            I => \N__46830\
        );

    \I__11395\ : ClkMux
    port map (
            O => \N__47419\,
            I => \N__46830\
        );

    \I__11394\ : ClkMux
    port map (
            O => \N__47418\,
            I => \N__46830\
        );

    \I__11393\ : ClkMux
    port map (
            O => \N__47417\,
            I => \N__46830\
        );

    \I__11392\ : ClkMux
    port map (
            O => \N__47416\,
            I => \N__46830\
        );

    \I__11391\ : ClkMux
    port map (
            O => \N__47415\,
            I => \N__46830\
        );

    \I__11390\ : ClkMux
    port map (
            O => \N__47414\,
            I => \N__46830\
        );

    \I__11389\ : ClkMux
    port map (
            O => \N__47413\,
            I => \N__46830\
        );

    \I__11388\ : ClkMux
    port map (
            O => \N__47412\,
            I => \N__46830\
        );

    \I__11387\ : ClkMux
    port map (
            O => \N__47411\,
            I => \N__46830\
        );

    \I__11386\ : ClkMux
    port map (
            O => \N__47410\,
            I => \N__46830\
        );

    \I__11385\ : ClkMux
    port map (
            O => \N__47409\,
            I => \N__46830\
        );

    \I__11384\ : ClkMux
    port map (
            O => \N__47408\,
            I => \N__46830\
        );

    \I__11383\ : ClkMux
    port map (
            O => \N__47407\,
            I => \N__46830\
        );

    \I__11382\ : ClkMux
    port map (
            O => \N__47406\,
            I => \N__46830\
        );

    \I__11381\ : ClkMux
    port map (
            O => \N__47405\,
            I => \N__46830\
        );

    \I__11380\ : ClkMux
    port map (
            O => \N__47404\,
            I => \N__46830\
        );

    \I__11379\ : ClkMux
    port map (
            O => \N__47403\,
            I => \N__46830\
        );

    \I__11378\ : ClkMux
    port map (
            O => \N__47402\,
            I => \N__46830\
        );

    \I__11377\ : ClkMux
    port map (
            O => \N__47401\,
            I => \N__46830\
        );

    \I__11376\ : ClkMux
    port map (
            O => \N__47400\,
            I => \N__46830\
        );

    \I__11375\ : ClkMux
    port map (
            O => \N__47399\,
            I => \N__46830\
        );

    \I__11374\ : ClkMux
    port map (
            O => \N__47398\,
            I => \N__46830\
        );

    \I__11373\ : ClkMux
    port map (
            O => \N__47397\,
            I => \N__46830\
        );

    \I__11372\ : ClkMux
    port map (
            O => \N__47396\,
            I => \N__46830\
        );

    \I__11371\ : ClkMux
    port map (
            O => \N__47395\,
            I => \N__46830\
        );

    \I__11370\ : ClkMux
    port map (
            O => \N__47394\,
            I => \N__46830\
        );

    \I__11369\ : ClkMux
    port map (
            O => \N__47393\,
            I => \N__46830\
        );

    \I__11368\ : ClkMux
    port map (
            O => \N__47392\,
            I => \N__46830\
        );

    \I__11367\ : ClkMux
    port map (
            O => \N__47391\,
            I => \N__46830\
        );

    \I__11366\ : ClkMux
    port map (
            O => \N__47390\,
            I => \N__46830\
        );

    \I__11365\ : ClkMux
    port map (
            O => \N__47389\,
            I => \N__46830\
        );

    \I__11364\ : ClkMux
    port map (
            O => \N__47388\,
            I => \N__46830\
        );

    \I__11363\ : ClkMux
    port map (
            O => \N__47387\,
            I => \N__46830\
        );

    \I__11362\ : ClkMux
    port map (
            O => \N__47386\,
            I => \N__46830\
        );

    \I__11361\ : ClkMux
    port map (
            O => \N__47385\,
            I => \N__46830\
        );

    \I__11360\ : ClkMux
    port map (
            O => \N__47384\,
            I => \N__46830\
        );

    \I__11359\ : ClkMux
    port map (
            O => \N__47383\,
            I => \N__46830\
        );

    \I__11358\ : ClkMux
    port map (
            O => \N__47382\,
            I => \N__46830\
        );

    \I__11357\ : ClkMux
    port map (
            O => \N__47381\,
            I => \N__46830\
        );

    \I__11356\ : ClkMux
    port map (
            O => \N__47380\,
            I => \N__46830\
        );

    \I__11355\ : ClkMux
    port map (
            O => \N__47379\,
            I => \N__46830\
        );

    \I__11354\ : ClkMux
    port map (
            O => \N__47378\,
            I => \N__46830\
        );

    \I__11353\ : ClkMux
    port map (
            O => \N__47377\,
            I => \N__46830\
        );

    \I__11352\ : ClkMux
    port map (
            O => \N__47376\,
            I => \N__46830\
        );

    \I__11351\ : ClkMux
    port map (
            O => \N__47375\,
            I => \N__46830\
        );

    \I__11350\ : ClkMux
    port map (
            O => \N__47374\,
            I => \N__46830\
        );

    \I__11349\ : ClkMux
    port map (
            O => \N__47373\,
            I => \N__46830\
        );

    \I__11348\ : ClkMux
    port map (
            O => \N__47372\,
            I => \N__46830\
        );

    \I__11347\ : ClkMux
    port map (
            O => \N__47371\,
            I => \N__46830\
        );

    \I__11346\ : ClkMux
    port map (
            O => \N__47370\,
            I => \N__46830\
        );

    \I__11345\ : ClkMux
    port map (
            O => \N__47369\,
            I => \N__46830\
        );

    \I__11344\ : ClkMux
    port map (
            O => \N__47368\,
            I => \N__46830\
        );

    \I__11343\ : ClkMux
    port map (
            O => \N__47367\,
            I => \N__46830\
        );

    \I__11342\ : ClkMux
    port map (
            O => \N__47366\,
            I => \N__46830\
        );

    \I__11341\ : ClkMux
    port map (
            O => \N__47365\,
            I => \N__46830\
        );

    \I__11340\ : ClkMux
    port map (
            O => \N__47364\,
            I => \N__46830\
        );

    \I__11339\ : ClkMux
    port map (
            O => \N__47363\,
            I => \N__46830\
        );

    \I__11338\ : ClkMux
    port map (
            O => \N__47362\,
            I => \N__46830\
        );

    \I__11337\ : ClkMux
    port map (
            O => \N__47361\,
            I => \N__46830\
        );

    \I__11336\ : ClkMux
    port map (
            O => \N__47360\,
            I => \N__46830\
        );

    \I__11335\ : ClkMux
    port map (
            O => \N__47359\,
            I => \N__46830\
        );

    \I__11334\ : ClkMux
    port map (
            O => \N__47358\,
            I => \N__46830\
        );

    \I__11333\ : ClkMux
    port map (
            O => \N__47357\,
            I => \N__46830\
        );

    \I__11332\ : ClkMux
    port map (
            O => \N__47356\,
            I => \N__46830\
        );

    \I__11331\ : ClkMux
    port map (
            O => \N__47355\,
            I => \N__46830\
        );

    \I__11330\ : ClkMux
    port map (
            O => \N__47354\,
            I => \N__46830\
        );

    \I__11329\ : ClkMux
    port map (
            O => \N__47353\,
            I => \N__46830\
        );

    \I__11328\ : ClkMux
    port map (
            O => \N__47352\,
            I => \N__46830\
        );

    \I__11327\ : ClkMux
    port map (
            O => \N__47351\,
            I => \N__46830\
        );

    \I__11326\ : ClkMux
    port map (
            O => \N__47350\,
            I => \N__46830\
        );

    \I__11325\ : ClkMux
    port map (
            O => \N__47349\,
            I => \N__46830\
        );

    \I__11324\ : ClkMux
    port map (
            O => \N__47348\,
            I => \N__46830\
        );

    \I__11323\ : ClkMux
    port map (
            O => \N__47347\,
            I => \N__46830\
        );

    \I__11322\ : ClkMux
    port map (
            O => \N__47346\,
            I => \N__46830\
        );

    \I__11321\ : ClkMux
    port map (
            O => \N__47345\,
            I => \N__46830\
        );

    \I__11320\ : ClkMux
    port map (
            O => \N__47344\,
            I => \N__46830\
        );

    \I__11319\ : ClkMux
    port map (
            O => \N__47343\,
            I => \N__46830\
        );

    \I__11318\ : ClkMux
    port map (
            O => \N__47342\,
            I => \N__46830\
        );

    \I__11317\ : ClkMux
    port map (
            O => \N__47341\,
            I => \N__46830\
        );

    \I__11316\ : ClkMux
    port map (
            O => \N__47340\,
            I => \N__46830\
        );

    \I__11315\ : ClkMux
    port map (
            O => \N__47339\,
            I => \N__46830\
        );

    \I__11314\ : ClkMux
    port map (
            O => \N__47338\,
            I => \N__46830\
        );

    \I__11313\ : ClkMux
    port map (
            O => \N__47337\,
            I => \N__46830\
        );

    \I__11312\ : ClkMux
    port map (
            O => \N__47336\,
            I => \N__46830\
        );

    \I__11311\ : ClkMux
    port map (
            O => \N__47335\,
            I => \N__46830\
        );

    \I__11310\ : ClkMux
    port map (
            O => \N__47334\,
            I => \N__46830\
        );

    \I__11309\ : ClkMux
    port map (
            O => \N__47333\,
            I => \N__46830\
        );

    \I__11308\ : ClkMux
    port map (
            O => \N__47332\,
            I => \N__46830\
        );

    \I__11307\ : ClkMux
    port map (
            O => \N__47331\,
            I => \N__46830\
        );

    \I__11306\ : ClkMux
    port map (
            O => \N__47330\,
            I => \N__46830\
        );

    \I__11305\ : ClkMux
    port map (
            O => \N__47329\,
            I => \N__46830\
        );

    \I__11304\ : ClkMux
    port map (
            O => \N__47328\,
            I => \N__46830\
        );

    \I__11303\ : ClkMux
    port map (
            O => \N__47327\,
            I => \N__46830\
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__47326\,
            I => \N__46830\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__47325\,
            I => \N__46830\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__47324\,
            I => \N__46830\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__47323\,
            I => \N__46830\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__47322\,
            I => \N__46830\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__47321\,
            I => \N__46830\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__47320\,
            I => \N__46830\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__47319\,
            I => \N__46830\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__47318\,
            I => \N__46830\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__47317\,
            I => \N__46830\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__47316\,
            I => \N__46830\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__47315\,
            I => \N__46830\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__47314\,
            I => \N__46830\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__47313\,
            I => \N__46830\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__47312\,
            I => \N__46830\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__47311\,
            I => \N__46830\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__47310\,
            I => \N__46830\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__47309\,
            I => \N__46830\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__47308\,
            I => \N__46830\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__47307\,
            I => \N__46830\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__47306\,
            I => \N__46830\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__47305\,
            I => \N__46830\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__47304\,
            I => \N__46830\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__47303\,
            I => \N__46830\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__47302\,
            I => \N__46830\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__47301\,
            I => \N__46830\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__47300\,
            I => \N__46830\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__47299\,
            I => \N__46830\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__47298\,
            I => \N__46830\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__47297\,
            I => \N__46830\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__47296\,
            I => \N__46830\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__47295\,
            I => \N__46830\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__47294\,
            I => \N__46830\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__47293\,
            I => \N__46830\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__47292\,
            I => \N__46830\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__47291\,
            I => \N__46830\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__47290\,
            I => \N__46830\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__47289\,
            I => \N__46830\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__47288\,
            I => \N__46830\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__47287\,
            I => \N__46830\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__47286\,
            I => \N__46830\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__47285\,
            I => \N__46830\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__47284\,
            I => \N__46830\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__47283\,
            I => \N__46830\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__47282\,
            I => \N__46830\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__47281\,
            I => \N__46830\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__47280\,
            I => \N__46830\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47279\,
            I => \N__46830\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47278\,
            I => \N__46830\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47277\,
            I => \N__46830\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47276\,
            I => \N__46830\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47275\,
            I => \N__46830\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47274\,
            I => \N__46830\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47273\,
            I => \N__46830\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47272\,
            I => \N__46830\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47271\,
            I => \N__46830\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47270\,
            I => \N__46830\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47269\,
            I => \N__46830\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47268\,
            I => \N__46830\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47267\,
            I => \N__46830\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47266\,
            I => \N__46830\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47265\,
            I => \N__46830\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47264\,
            I => \N__46830\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47263\,
            I => \N__46830\
        );

    \I__11238\ : GlobalMux
    port map (
            O => \N__46830\,
            I => \N__46827\
        );

    \I__11237\ : gio2CtrlBuf
    port map (
            O => \N__46827\,
            I => clk_system_c_g
        );

    \I__11236\ : CEMux
    port map (
            O => \N__46824\,
            I => \N__46695\
        );

    \I__11235\ : CEMux
    port map (
            O => \N__46823\,
            I => \N__46695\
        );

    \I__11234\ : CEMux
    port map (
            O => \N__46822\,
            I => \N__46695\
        );

    \I__11233\ : CEMux
    port map (
            O => \N__46821\,
            I => \N__46695\
        );

    \I__11232\ : CEMux
    port map (
            O => \N__46820\,
            I => \N__46695\
        );

    \I__11231\ : CEMux
    port map (
            O => \N__46819\,
            I => \N__46695\
        );

    \I__11230\ : CEMux
    port map (
            O => \N__46818\,
            I => \N__46695\
        );

    \I__11229\ : CEMux
    port map (
            O => \N__46817\,
            I => \N__46695\
        );

    \I__11228\ : CEMux
    port map (
            O => \N__46816\,
            I => \N__46695\
        );

    \I__11227\ : CEMux
    port map (
            O => \N__46815\,
            I => \N__46695\
        );

    \I__11226\ : CEMux
    port map (
            O => \N__46814\,
            I => \N__46695\
        );

    \I__11225\ : CEMux
    port map (
            O => \N__46813\,
            I => \N__46695\
        );

    \I__11224\ : CEMux
    port map (
            O => \N__46812\,
            I => \N__46695\
        );

    \I__11223\ : CEMux
    port map (
            O => \N__46811\,
            I => \N__46695\
        );

    \I__11222\ : CEMux
    port map (
            O => \N__46810\,
            I => \N__46695\
        );

    \I__11221\ : CEMux
    port map (
            O => \N__46809\,
            I => \N__46695\
        );

    \I__11220\ : CEMux
    port map (
            O => \N__46808\,
            I => \N__46695\
        );

    \I__11219\ : CEMux
    port map (
            O => \N__46807\,
            I => \N__46695\
        );

    \I__11218\ : CEMux
    port map (
            O => \N__46806\,
            I => \N__46695\
        );

    \I__11217\ : CEMux
    port map (
            O => \N__46805\,
            I => \N__46695\
        );

    \I__11216\ : CEMux
    port map (
            O => \N__46804\,
            I => \N__46695\
        );

    \I__11215\ : CEMux
    port map (
            O => \N__46803\,
            I => \N__46695\
        );

    \I__11214\ : CEMux
    port map (
            O => \N__46802\,
            I => \N__46695\
        );

    \I__11213\ : CEMux
    port map (
            O => \N__46801\,
            I => \N__46695\
        );

    \I__11212\ : CEMux
    port map (
            O => \N__46800\,
            I => \N__46695\
        );

    \I__11211\ : CEMux
    port map (
            O => \N__46799\,
            I => \N__46695\
        );

    \I__11210\ : CEMux
    port map (
            O => \N__46798\,
            I => \N__46695\
        );

    \I__11209\ : CEMux
    port map (
            O => \N__46797\,
            I => \N__46695\
        );

    \I__11208\ : CEMux
    port map (
            O => \N__46796\,
            I => \N__46695\
        );

    \I__11207\ : CEMux
    port map (
            O => \N__46795\,
            I => \N__46695\
        );

    \I__11206\ : CEMux
    port map (
            O => \N__46794\,
            I => \N__46695\
        );

    \I__11205\ : CEMux
    port map (
            O => \N__46793\,
            I => \N__46695\
        );

    \I__11204\ : CEMux
    port map (
            O => \N__46792\,
            I => \N__46695\
        );

    \I__11203\ : CEMux
    port map (
            O => \N__46791\,
            I => \N__46695\
        );

    \I__11202\ : CEMux
    port map (
            O => \N__46790\,
            I => \N__46695\
        );

    \I__11201\ : CEMux
    port map (
            O => \N__46789\,
            I => \N__46695\
        );

    \I__11200\ : CEMux
    port map (
            O => \N__46788\,
            I => \N__46695\
        );

    \I__11199\ : CEMux
    port map (
            O => \N__46787\,
            I => \N__46695\
        );

    \I__11198\ : CEMux
    port map (
            O => \N__46786\,
            I => \N__46695\
        );

    \I__11197\ : CEMux
    port map (
            O => \N__46785\,
            I => \N__46695\
        );

    \I__11196\ : CEMux
    port map (
            O => \N__46784\,
            I => \N__46695\
        );

    \I__11195\ : CEMux
    port map (
            O => \N__46783\,
            I => \N__46695\
        );

    \I__11194\ : CEMux
    port map (
            O => \N__46782\,
            I => \N__46695\
        );

    \I__11193\ : GlobalMux
    port map (
            O => \N__46695\,
            I => \N__46692\
        );

    \I__11192\ : gio2CtrlBuf
    port map (
            O => \N__46692\,
            I => \pid_alt.N_410_0_g\
        );

    \I__11191\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46671\
        );

    \I__11190\ : InMux
    port map (
            O => \N__46688\,
            I => \N__46668\
        );

    \I__11189\ : InMux
    port map (
            O => \N__46687\,
            I => \N__46663\
        );

    \I__11188\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46663\
        );

    \I__11187\ : InMux
    port map (
            O => \N__46685\,
            I => \N__46658\
        );

    \I__11186\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46658\
        );

    \I__11185\ : InMux
    port map (
            O => \N__46683\,
            I => \N__46655\
        );

    \I__11184\ : InMux
    port map (
            O => \N__46682\,
            I => \N__46652\
        );

    \I__11183\ : InMux
    port map (
            O => \N__46681\,
            I => \N__46649\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46646\
        );

    \I__11181\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46643\
        );

    \I__11180\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46640\
        );

    \I__11179\ : InMux
    port map (
            O => \N__46677\,
            I => \N__46635\
        );

    \I__11178\ : InMux
    port map (
            O => \N__46676\,
            I => \N__46635\
        );

    \I__11177\ : InMux
    port map (
            O => \N__46675\,
            I => \N__46632\
        );

    \I__11176\ : InMux
    port map (
            O => \N__46674\,
            I => \N__46629\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__46671\,
            I => \N__46582\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__46668\,
            I => \N__46579\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__46663\,
            I => \N__46576\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__46658\,
            I => \N__46573\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__46655\,
            I => \N__46570\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__46652\,
            I => \N__46567\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__46649\,
            I => \N__46564\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46646\,
            I => \N__46561\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__46643\,
            I => \N__46558\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__46640\,
            I => \N__46555\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__46635\,
            I => \N__46552\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__46632\,
            I => \N__46549\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__46629\,
            I => \N__46546\
        );

    \I__11162\ : SRMux
    port map (
            O => \N__46628\,
            I => \N__46431\
        );

    \I__11161\ : SRMux
    port map (
            O => \N__46627\,
            I => \N__46431\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__46626\,
            I => \N__46431\
        );

    \I__11159\ : SRMux
    port map (
            O => \N__46625\,
            I => \N__46431\
        );

    \I__11158\ : SRMux
    port map (
            O => \N__46624\,
            I => \N__46431\
        );

    \I__11157\ : SRMux
    port map (
            O => \N__46623\,
            I => \N__46431\
        );

    \I__11156\ : SRMux
    port map (
            O => \N__46622\,
            I => \N__46431\
        );

    \I__11155\ : SRMux
    port map (
            O => \N__46621\,
            I => \N__46431\
        );

    \I__11154\ : SRMux
    port map (
            O => \N__46620\,
            I => \N__46431\
        );

    \I__11153\ : SRMux
    port map (
            O => \N__46619\,
            I => \N__46431\
        );

    \I__11152\ : SRMux
    port map (
            O => \N__46618\,
            I => \N__46431\
        );

    \I__11151\ : SRMux
    port map (
            O => \N__46617\,
            I => \N__46431\
        );

    \I__11150\ : SRMux
    port map (
            O => \N__46616\,
            I => \N__46431\
        );

    \I__11149\ : SRMux
    port map (
            O => \N__46615\,
            I => \N__46431\
        );

    \I__11148\ : SRMux
    port map (
            O => \N__46614\,
            I => \N__46431\
        );

    \I__11147\ : SRMux
    port map (
            O => \N__46613\,
            I => \N__46431\
        );

    \I__11146\ : SRMux
    port map (
            O => \N__46612\,
            I => \N__46431\
        );

    \I__11145\ : SRMux
    port map (
            O => \N__46611\,
            I => \N__46431\
        );

    \I__11144\ : SRMux
    port map (
            O => \N__46610\,
            I => \N__46431\
        );

    \I__11143\ : SRMux
    port map (
            O => \N__46609\,
            I => \N__46431\
        );

    \I__11142\ : SRMux
    port map (
            O => \N__46608\,
            I => \N__46431\
        );

    \I__11141\ : SRMux
    port map (
            O => \N__46607\,
            I => \N__46431\
        );

    \I__11140\ : SRMux
    port map (
            O => \N__46606\,
            I => \N__46431\
        );

    \I__11139\ : SRMux
    port map (
            O => \N__46605\,
            I => \N__46431\
        );

    \I__11138\ : SRMux
    port map (
            O => \N__46604\,
            I => \N__46431\
        );

    \I__11137\ : SRMux
    port map (
            O => \N__46603\,
            I => \N__46431\
        );

    \I__11136\ : SRMux
    port map (
            O => \N__46602\,
            I => \N__46431\
        );

    \I__11135\ : SRMux
    port map (
            O => \N__46601\,
            I => \N__46431\
        );

    \I__11134\ : SRMux
    port map (
            O => \N__46600\,
            I => \N__46431\
        );

    \I__11133\ : SRMux
    port map (
            O => \N__46599\,
            I => \N__46431\
        );

    \I__11132\ : SRMux
    port map (
            O => \N__46598\,
            I => \N__46431\
        );

    \I__11131\ : SRMux
    port map (
            O => \N__46597\,
            I => \N__46431\
        );

    \I__11130\ : SRMux
    port map (
            O => \N__46596\,
            I => \N__46431\
        );

    \I__11129\ : SRMux
    port map (
            O => \N__46595\,
            I => \N__46431\
        );

    \I__11128\ : SRMux
    port map (
            O => \N__46594\,
            I => \N__46431\
        );

    \I__11127\ : SRMux
    port map (
            O => \N__46593\,
            I => \N__46431\
        );

    \I__11126\ : SRMux
    port map (
            O => \N__46592\,
            I => \N__46431\
        );

    \I__11125\ : SRMux
    port map (
            O => \N__46591\,
            I => \N__46431\
        );

    \I__11124\ : SRMux
    port map (
            O => \N__46590\,
            I => \N__46431\
        );

    \I__11123\ : SRMux
    port map (
            O => \N__46589\,
            I => \N__46431\
        );

    \I__11122\ : SRMux
    port map (
            O => \N__46588\,
            I => \N__46431\
        );

    \I__11121\ : SRMux
    port map (
            O => \N__46587\,
            I => \N__46431\
        );

    \I__11120\ : SRMux
    port map (
            O => \N__46586\,
            I => \N__46431\
        );

    \I__11119\ : SRMux
    port map (
            O => \N__46585\,
            I => \N__46431\
        );

    \I__11118\ : Glb2LocalMux
    port map (
            O => \N__46582\,
            I => \N__46431\
        );

    \I__11117\ : Glb2LocalMux
    port map (
            O => \N__46579\,
            I => \N__46431\
        );

    \I__11116\ : Glb2LocalMux
    port map (
            O => \N__46576\,
            I => \N__46431\
        );

    \I__11115\ : Glb2LocalMux
    port map (
            O => \N__46573\,
            I => \N__46431\
        );

    \I__11114\ : Glb2LocalMux
    port map (
            O => \N__46570\,
            I => \N__46431\
        );

    \I__11113\ : Glb2LocalMux
    port map (
            O => \N__46567\,
            I => \N__46431\
        );

    \I__11112\ : Glb2LocalMux
    port map (
            O => \N__46564\,
            I => \N__46431\
        );

    \I__11111\ : Glb2LocalMux
    port map (
            O => \N__46561\,
            I => \N__46431\
        );

    \I__11110\ : Glb2LocalMux
    port map (
            O => \N__46558\,
            I => \N__46431\
        );

    \I__11109\ : Glb2LocalMux
    port map (
            O => \N__46555\,
            I => \N__46431\
        );

    \I__11108\ : Glb2LocalMux
    port map (
            O => \N__46552\,
            I => \N__46431\
        );

    \I__11107\ : Glb2LocalMux
    port map (
            O => \N__46549\,
            I => \N__46431\
        );

    \I__11106\ : Glb2LocalMux
    port map (
            O => \N__46546\,
            I => \N__46431\
        );

    \I__11105\ : GlobalMux
    port map (
            O => \N__46431\,
            I => \N__46428\
        );

    \I__11104\ : gio2CtrlBuf
    port map (
            O => \N__46428\,
            I => \N_411_g\
        );

    \I__11103\ : InMux
    port map (
            O => \N__46425\,
            I => \N__46422\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__46422\,
            I => \N__46418\
        );

    \I__11101\ : InMux
    port map (
            O => \N__46421\,
            I => \N__46415\
        );

    \I__11100\ : Span12Mux_s2_h
    port map (
            O => \N__46418\,
            I => \N__46412\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__46415\,
            I => \N__46409\
        );

    \I__11098\ : Span12Mux_h
    port map (
            O => \N__46412\,
            I => \N__46406\
        );

    \I__11097\ : Span4Mux_v
    port map (
            O => \N__46409\,
            I => \N__46403\
        );

    \I__11096\ : Odrv12
    port map (
            O => \N__46406\,
            I => \pid_alt.error_filt_6\
        );

    \I__11095\ : Odrv4
    port map (
            O => \N__46403\,
            I => \pid_alt.error_filt_6\
        );

    \I__11094\ : InMux
    port map (
            O => \N__46398\,
            I => \N__46395\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__46395\,
            I => \pid_alt.error_filt_prevZ0Z_6\
        );

    \I__11092\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46389\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__46389\,
            I => \N__46385\
        );

    \I__11090\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46382\
        );

    \I__11089\ : Span12Mux_s3_h
    port map (
            O => \N__46385\,
            I => \N__46379\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__46382\,
            I => \N__46376\
        );

    \I__11087\ : Span12Mux_h
    port map (
            O => \N__46379\,
            I => \N__46373\
        );

    \I__11086\ : Span4Mux_v
    port map (
            O => \N__46376\,
            I => \N__46370\
        );

    \I__11085\ : Odrv12
    port map (
            O => \N__46373\,
            I => \pid_alt.error_filt_7\
        );

    \I__11084\ : Odrv4
    port map (
            O => \N__46370\,
            I => \pid_alt.error_filt_7\
        );

    \I__11083\ : InMux
    port map (
            O => \N__46365\,
            I => \N__46362\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46362\,
            I => \pid_alt.error_filt_prevZ0Z_7\
        );

    \I__11081\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46356\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46353\
        );

    \I__11079\ : Span4Mux_v
    port map (
            O => \N__46353\,
            I => \N__46350\
        );

    \I__11078\ : Span4Mux_h
    port map (
            O => \N__46350\,
            I => \N__46347\
        );

    \I__11077\ : Span4Mux_h
    port map (
            O => \N__46347\,
            I => \N__46344\
        );

    \I__11076\ : Span4Mux_h
    port map (
            O => \N__46344\,
            I => \N__46340\
        );

    \I__11075\ : InMux
    port map (
            O => \N__46343\,
            I => \N__46337\
        );

    \I__11074\ : Span4Mux_h
    port map (
            O => \N__46340\,
            I => \N__46334\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__46337\,
            I => \N__46331\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__46334\,
            I => \N__46328\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__46331\,
            I => \N__46325\
        );

    \I__11070\ : Odrv4
    port map (
            O => \N__46328\,
            I => \pid_alt.error_filt_9\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__46325\,
            I => \pid_alt.error_filt_9\
        );

    \I__11068\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46317\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__46317\,
            I => \pid_alt.error_filt_prevZ0Z_9\
        );

    \I__11066\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46311\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__46311\,
            I => \N__46307\
        );

    \I__11064\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46304\
        );

    \I__11063\ : Span12Mux_s7_h
    port map (
            O => \N__46307\,
            I => \N__46301\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__46304\,
            I => \N__46298\
        );

    \I__11061\ : Span12Mux_h
    port map (
            O => \N__46301\,
            I => \N__46295\
        );

    \I__11060\ : Span4Mux_s1_h
    port map (
            O => \N__46298\,
            I => \N__46292\
        );

    \I__11059\ : Odrv12
    port map (
            O => \N__46295\,
            I => \pid_alt.error_filt_3\
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__46292\,
            I => \pid_alt.error_filt_3\
        );

    \I__11057\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__46284\,
            I => \pid_alt.error_filt_prevZ0Z_3\
        );

    \I__11055\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46278\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__46278\,
            I => \N__46274\
        );

    \I__11053\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46271\
        );

    \I__11052\ : Span12Mux_s2_h
    port map (
            O => \N__46274\,
            I => \N__46268\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__46271\,
            I => \N__46265\
        );

    \I__11050\ : Span12Mux_h
    port map (
            O => \N__46268\,
            I => \N__46262\
        );

    \I__11049\ : Span4Mux_v
    port map (
            O => \N__46265\,
            I => \N__46259\
        );

    \I__11048\ : Odrv12
    port map (
            O => \N__46262\,
            I => \pid_alt.error_filt_14\
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__46259\,
            I => \pid_alt.error_filt_14\
        );

    \I__11046\ : InMux
    port map (
            O => \N__46254\,
            I => \N__46251\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__46251\,
            I => \pid_alt.error_filt_prevZ0Z_14\
        );

    \I__11044\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46245\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46245\,
            I => \N__46242\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__46242\,
            I => \pid_alt.O_0_11\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__46239\,
            I => \N__46236\
        );

    \I__11040\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46233\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__46233\,
            I => \N__46230\
        );

    \I__11038\ : Span12Mux_h
    port map (
            O => \N__46230\,
            I => \N__46227\
        );

    \I__11037\ : Odrv12
    port map (
            O => \N__46227\,
            I => \pid_alt.error_i_regZ0Z_7\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46218\
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__46218\,
            I => \pid_alt.O_0_10\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46215\,
            I => \N__46212\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__46212\,
            I => \N__46209\
        );

    \I__11031\ : Span12Mux_h
    port map (
            O => \N__46209\,
            I => \N__46206\
        );

    \I__11030\ : Odrv12
    port map (
            O => \N__46206\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__11029\ : InMux
    port map (
            O => \N__46203\,
            I => \N__46200\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__46200\,
            I => \N__46197\
        );

    \I__11027\ : Odrv4
    port map (
            O => \N__46197\,
            I => \pid_alt.O_19\
        );

    \I__11026\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46191\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__46191\,
            I => \N__46188\
        );

    \I__11024\ : Span4Mux_h
    port map (
            O => \N__46188\,
            I => \N__46185\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__46185\,
            I => \N__46182\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__11021\ : Odrv4
    port map (
            O => \N__46179\,
            I => \pid_alt.error_i_regZ0Z_15\
        );

    \I__11020\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46173\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__46173\,
            I => \N__46169\
        );

    \I__11018\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46166\
        );

    \I__11017\ : Span12Mux_h
    port map (
            O => \N__46169\,
            I => \N__46163\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__46166\,
            I => \N__46160\
        );

    \I__11015\ : Span12Mux_h
    port map (
            O => \N__46163\,
            I => \N__46157\
        );

    \I__11014\ : Span4Mux_s1_h
    port map (
            O => \N__46160\,
            I => \N__46154\
        );

    \I__11013\ : Odrv12
    port map (
            O => \N__46157\,
            I => \pid_alt.error_filt_2\
        );

    \I__11012\ : Odrv4
    port map (
            O => \N__46154\,
            I => \pid_alt.error_filt_2\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46149\,
            I => \N__46146\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46143\
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__46143\,
            I => \pid_alt.error_filt_prevZ0Z_2\
        );

    \I__11008\ : InMux
    port map (
            O => \N__46140\,
            I => \N__46137\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__46137\,
            I => \N__46133\
        );

    \I__11006\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46130\
        );

    \I__11005\ : Span12Mux_h
    port map (
            O => \N__46133\,
            I => \N__46127\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__46130\,
            I => \N__46124\
        );

    \I__11003\ : Span12Mux_h
    port map (
            O => \N__46127\,
            I => \N__46121\
        );

    \I__11002\ : Span4Mux_v
    port map (
            O => \N__46124\,
            I => \N__46118\
        );

    \I__11001\ : Odrv12
    port map (
            O => \N__46121\,
            I => \pid_alt.error_filt_10\
        );

    \I__11000\ : Odrv4
    port map (
            O => \N__46118\,
            I => \pid_alt.error_filt_10\
        );

    \I__10999\ : InMux
    port map (
            O => \N__46113\,
            I => \N__46110\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__46110\,
            I => \N__46107\
        );

    \I__10997\ : Odrv4
    port map (
            O => \N__46107\,
            I => \pid_alt.error_filt_prevZ0Z_10\
        );

    \I__10996\ : InMux
    port map (
            O => \N__46104\,
            I => \N__46101\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__46101\,
            I => \N__46098\
        );

    \I__10994\ : Span4Mux_v
    port map (
            O => \N__46098\,
            I => \N__46095\
        );

    \I__10993\ : Span4Mux_h
    port map (
            O => \N__46095\,
            I => \N__46091\
        );

    \I__10992\ : InMux
    port map (
            O => \N__46094\,
            I => \N__46088\
        );

    \I__10991\ : Sp12to4
    port map (
            O => \N__46091\,
            I => \N__46085\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__46088\,
            I => \N__46082\
        );

    \I__10989\ : Span12Mux_h
    port map (
            O => \N__46085\,
            I => \N__46079\
        );

    \I__10988\ : Span4Mux_v
    port map (
            O => \N__46082\,
            I => \N__46076\
        );

    \I__10987\ : Odrv12
    port map (
            O => \N__46079\,
            I => \pid_alt.error_filt_11\
        );

    \I__10986\ : Odrv4
    port map (
            O => \N__46076\,
            I => \pid_alt.error_filt_11\
        );

    \I__10985\ : InMux
    port map (
            O => \N__46071\,
            I => \N__46068\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__46068\,
            I => \N__46065\
        );

    \I__10983\ : Odrv4
    port map (
            O => \N__46065\,
            I => \pid_alt.error_filt_prevZ0Z_11\
        );

    \I__10982\ : InMux
    port map (
            O => \N__46062\,
            I => \N__46059\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__46059\,
            I => \N__46056\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__46056\,
            I => \N__46052\
        );

    \I__10979\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46049\
        );

    \I__10978\ : Sp12to4
    port map (
            O => \N__46052\,
            I => \N__46046\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__46049\,
            I => \N__46043\
        );

    \I__10976\ : Span12Mux_h
    port map (
            O => \N__46046\,
            I => \N__46040\
        );

    \I__10975\ : Span4Mux_v
    port map (
            O => \N__46043\,
            I => \N__46037\
        );

    \I__10974\ : Odrv12
    port map (
            O => \N__46040\,
            I => \pid_alt.error_filt_12\
        );

    \I__10973\ : Odrv4
    port map (
            O => \N__46037\,
            I => \pid_alt.error_filt_12\
        );

    \I__10972\ : InMux
    port map (
            O => \N__46032\,
            I => \N__46029\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__46029\,
            I => \N__46026\
        );

    \I__10970\ : Odrv4
    port map (
            O => \N__46026\,
            I => \pid_alt.error_filt_prevZ0Z_12\
        );

    \I__10969\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__46020\,
            I => \N__46016\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46019\,
            I => \N__46013\
        );

    \I__10966\ : Span12Mux_v
    port map (
            O => \N__46016\,
            I => \N__46010\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__46013\,
            I => \N__46007\
        );

    \I__10964\ : Span12Mux_h
    port map (
            O => \N__46010\,
            I => \N__46004\
        );

    \I__10963\ : Span4Mux_v
    port map (
            O => \N__46007\,
            I => \N__46001\
        );

    \I__10962\ : Odrv12
    port map (
            O => \N__46004\,
            I => \pid_alt.error_filt_13\
        );

    \I__10961\ : Odrv4
    port map (
            O => \N__46001\,
            I => \pid_alt.error_filt_13\
        );

    \I__10960\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45993\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__45993\,
            I => \N__45990\
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__45990\,
            I => \pid_alt.error_filt_prevZ0Z_13\
        );

    \I__10957\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45984\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__45984\,
            I => \N__45980\
        );

    \I__10955\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45977\
        );

    \I__10954\ : Span4Mux_v
    port map (
            O => \N__45980\,
            I => \N__45974\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__45977\,
            I => \N__45971\
        );

    \I__10952\ : Sp12to4
    port map (
            O => \N__45974\,
            I => \N__45968\
        );

    \I__10951\ : Span4Mux_v
    port map (
            O => \N__45971\,
            I => \N__45965\
        );

    \I__10950\ : Span12Mux_h
    port map (
            O => \N__45968\,
            I => \N__45962\
        );

    \I__10949\ : Span4Mux_v
    port map (
            O => \N__45965\,
            I => \N__45959\
        );

    \I__10948\ : Odrv12
    port map (
            O => \N__45962\,
            I => \pid_alt.error_filt_15\
        );

    \I__10947\ : Odrv4
    port map (
            O => \N__45959\,
            I => \pid_alt.error_filt_15\
        );

    \I__10946\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__45951\,
            I => \N__45948\
        );

    \I__10944\ : Span4Mux_s0_h
    port map (
            O => \N__45948\,
            I => \N__45945\
        );

    \I__10943\ : Odrv4
    port map (
            O => \N__45945\,
            I => \pid_alt.error_filt_prevZ0Z_15\
        );

    \I__10942\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45939\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__45939\,
            I => \N__45936\
        );

    \I__10940\ : Span4Mux_v
    port map (
            O => \N__45936\,
            I => \N__45932\
        );

    \I__10939\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45929\
        );

    \I__10938\ : Sp12to4
    port map (
            O => \N__45932\,
            I => \N__45926\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__45929\,
            I => \N__45923\
        );

    \I__10936\ : Span12Mux_s4_h
    port map (
            O => \N__45926\,
            I => \N__45920\
        );

    \I__10935\ : Span4Mux_v
    port map (
            O => \N__45923\,
            I => \N__45917\
        );

    \I__10934\ : Span12Mux_h
    port map (
            O => \N__45920\,
            I => \N__45914\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__45917\,
            I => \N__45911\
        );

    \I__10932\ : Odrv12
    port map (
            O => \N__45914\,
            I => \pid_alt.error_filt_16\
        );

    \I__10931\ : Odrv4
    port map (
            O => \N__45911\,
            I => \pid_alt.error_filt_16\
        );

    \I__10930\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45903\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__45903\,
            I => \N__45900\
        );

    \I__10928\ : Span4Mux_s0_h
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__10927\ : Odrv4
    port map (
            O => \N__45897\,
            I => \pid_alt.error_filt_prevZ0Z_16\
        );

    \I__10926\ : InMux
    port map (
            O => \N__45894\,
            I => \N__45890\
        );

    \I__10925\ : InMux
    port map (
            O => \N__45893\,
            I => \N__45887\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__45890\,
            I => \N__45884\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__45887\,
            I => \N__45881\
        );

    \I__10922\ : Span12Mux_h
    port map (
            O => \N__45884\,
            I => \N__45878\
        );

    \I__10921\ : Span4Mux_s2_h
    port map (
            O => \N__45881\,
            I => \N__45875\
        );

    \I__10920\ : Odrv12
    port map (
            O => \N__45878\,
            I => \pid_alt.error_filt_4\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__45875\,
            I => \pid_alt.error_filt_4\
        );

    \I__10918\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45867\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__45867\,
            I => \pid_alt.error_filt_prevZ0Z_4\
        );

    \I__10916\ : InMux
    port map (
            O => \N__45864\,
            I => \N__45861\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__45861\,
            I => \N__45857\
        );

    \I__10914\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45854\
        );

    \I__10913\ : Span12Mux_s1_h
    port map (
            O => \N__45857\,
            I => \N__45851\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__45854\,
            I => \N__45848\
        );

    \I__10911\ : Span12Mux_h
    port map (
            O => \N__45851\,
            I => \N__45845\
        );

    \I__10910\ : Span4Mux_s1_h
    port map (
            O => \N__45848\,
            I => \N__45842\
        );

    \I__10909\ : Odrv12
    port map (
            O => \N__45845\,
            I => \pid_alt.error_filt_5\
        );

    \I__10908\ : Odrv4
    port map (
            O => \N__45842\,
            I => \pid_alt.error_filt_5\
        );

    \I__10907\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45834\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__45834\,
            I => \pid_alt.error_filt_prevZ0Z_5\
        );

    \I__10905\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45828\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__45828\,
            I => \N__45825\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__45825\,
            I => \N__45822\
        );

    \I__10902\ : Odrv4
    port map (
            O => \N__45822\,
            I => \pid_alt.O_17\
        );

    \I__10901\ : CascadeMux
    port map (
            O => \N__45819\,
            I => \N__45816\
        );

    \I__10900\ : InMux
    port map (
            O => \N__45816\,
            I => \N__45813\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__10898\ : Span4Mux_h
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10897\ : Span4Mux_h
    port map (
            O => \N__45807\,
            I => \N__45804\
        );

    \I__10896\ : Span4Mux_h
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__10895\ : Odrv4
    port map (
            O => \N__45801\,
            I => \pid_alt.error_i_regZ0Z_13\
        );

    \I__10894\ : InMux
    port map (
            O => \N__45798\,
            I => \N__45795\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__45795\,
            I => \N__45792\
        );

    \I__10892\ : Span4Mux_s3_h
    port map (
            O => \N__45792\,
            I => \N__45789\
        );

    \I__10891\ : Span4Mux_v
    port map (
            O => \N__45789\,
            I => \N__45786\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__45786\,
            I => \N__45782\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45779\
        );

    \I__10888\ : Sp12to4
    port map (
            O => \N__45782\,
            I => \N__45776\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__45779\,
            I => \N__45773\
        );

    \I__10886\ : Span12Mux_h
    port map (
            O => \N__45776\,
            I => \N__45770\
        );

    \I__10885\ : Span12Mux_s1_h
    port map (
            O => \N__45773\,
            I => \N__45767\
        );

    \I__10884\ : Odrv12
    port map (
            O => \N__45770\,
            I => \pid_alt.error_filt_17\
        );

    \I__10883\ : Odrv12
    port map (
            O => \N__45767\,
            I => \pid_alt.error_filt_17\
        );

    \I__10882\ : InMux
    port map (
            O => \N__45762\,
            I => \N__45759\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__10880\ : Span4Mux_s1_h
    port map (
            O => \N__45756\,
            I => \N__45753\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__45753\,
            I => \pid_alt.error_filt_prevZ0Z_17\
        );

    \I__10878\ : InMux
    port map (
            O => \N__45750\,
            I => \N__45747\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__45747\,
            I => \N__45744\
        );

    \I__10876\ : Span4Mux_h
    port map (
            O => \N__45744\,
            I => \N__45741\
        );

    \I__10875\ : Span4Mux_h
    port map (
            O => \N__45741\,
            I => \N__45738\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__45738\,
            I => \N__45735\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__45735\,
            I => \N__45731\
        );

    \I__10872\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45728\
        );

    \I__10871\ : Span4Mux_h
    port map (
            O => \N__45731\,
            I => \N__45725\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__45728\,
            I => \N__45722\
        );

    \I__10869\ : Span4Mux_h
    port map (
            O => \N__45725\,
            I => \N__45717\
        );

    \I__10868\ : Span4Mux_v
    port map (
            O => \N__45722\,
            I => \N__45717\
        );

    \I__10867\ : Span4Mux_v
    port map (
            O => \N__45717\,
            I => \N__45714\
        );

    \I__10866\ : Odrv4
    port map (
            O => \N__45714\,
            I => \pid_alt.error_filt_18\
        );

    \I__10865\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__45708\,
            I => \N__45705\
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__45705\,
            I => \pid_alt.error_filt_prevZ0Z_18\
        );

    \I__10862\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45699\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__45699\,
            I => \N__45687\
        );

    \I__10860\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45678\
        );

    \I__10859\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45678\
        );

    \I__10858\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45678\
        );

    \I__10857\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45678\
        );

    \I__10856\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45667\
        );

    \I__10855\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45667\
        );

    \I__10854\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45667\
        );

    \I__10853\ : InMux
    port map (
            O => \N__45691\,
            I => \N__45667\
        );

    \I__10852\ : InMux
    port map (
            O => \N__45690\,
            I => \N__45667\
        );

    \I__10851\ : Span4Mux_s2_h
    port map (
            O => \N__45687\,
            I => \N__45664\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45659\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__45667\,
            I => \N__45659\
        );

    \I__10848\ : Sp12to4
    port map (
            O => \N__45664\,
            I => \N__45656\
        );

    \I__10847\ : Span4Mux_s1_h
    port map (
            O => \N__45659\,
            I => \N__45653\
        );

    \I__10846\ : Span12Mux_v
    port map (
            O => \N__45656\,
            I => \N__45650\
        );

    \I__10845\ : Span4Mux_v
    port map (
            O => \N__45653\,
            I => \N__45647\
        );

    \I__10844\ : Span12Mux_h
    port map (
            O => \N__45650\,
            I => \N__45644\
        );

    \I__10843\ : Span4Mux_v
    port map (
            O => \N__45647\,
            I => \N__45641\
        );

    \I__10842\ : Odrv12
    port map (
            O => \N__45644\,
            I => \pid_alt.error_filt_22\
        );

    \I__10841\ : Odrv4
    port map (
            O => \N__45641\,
            I => \pid_alt.error_filt_22\
        );

    \I__10840\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45619\
        );

    \I__10839\ : InMux
    port map (
            O => \N__45635\,
            I => \N__45619\
        );

    \I__10838\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45619\
        );

    \I__10837\ : InMux
    port map (
            O => \N__45633\,
            I => \N__45619\
        );

    \I__10836\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45608\
        );

    \I__10835\ : InMux
    port map (
            O => \N__45631\,
            I => \N__45608\
        );

    \I__10834\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45608\
        );

    \I__10833\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45608\
        );

    \I__10832\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45608\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__45619\,
            I => \N__45603\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__45608\,
            I => \N__45603\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__45603\,
            I => \pid_alt.error_filt_prevZ0Z_22\
        );

    \I__10828\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45597\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__45597\,
            I => \N__45593\
        );

    \I__10826\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45590\
        );

    \I__10825\ : Sp12to4
    port map (
            O => \N__45593\,
            I => \N__45587\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__45590\,
            I => \N__45584\
        );

    \I__10823\ : Span12Mux_v
    port map (
            O => \N__45587\,
            I => \N__45581\
        );

    \I__10822\ : Span4Mux_v
    port map (
            O => \N__45584\,
            I => \N__45578\
        );

    \I__10821\ : Span12Mux_h
    port map (
            O => \N__45581\,
            I => \N__45575\
        );

    \I__10820\ : Span4Mux_v
    port map (
            O => \N__45578\,
            I => \N__45572\
        );

    \I__10819\ : Odrv12
    port map (
            O => \N__45575\,
            I => \pid_alt.error_filt_20\
        );

    \I__10818\ : Odrv4
    port map (
            O => \N__45572\,
            I => \pid_alt.error_filt_20\
        );

    \I__10817\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45564\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__45564\,
            I => \pid_alt.error_filt_prevZ0Z_20\
        );

    \I__10815\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45558\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__45558\,
            I => \N__45554\
        );

    \I__10813\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45551\
        );

    \I__10812\ : Span12Mux_h
    port map (
            O => \N__45554\,
            I => \N__45548\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45545\
        );

    \I__10810\ : Span12Mux_h
    port map (
            O => \N__45548\,
            I => \N__45542\
        );

    \I__10809\ : Span4Mux_v
    port map (
            O => \N__45545\,
            I => \N__45539\
        );

    \I__10808\ : Odrv12
    port map (
            O => \N__45542\,
            I => \pid_alt.error_filt_8\
        );

    \I__10807\ : Odrv4
    port map (
            O => \N__45539\,
            I => \pid_alt.error_filt_8\
        );

    \I__10806\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45531\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45528\
        );

    \I__10804\ : Span4Mux_v
    port map (
            O => \N__45528\,
            I => \N__45525\
        );

    \I__10803\ : Odrv4
    port map (
            O => \N__45525\,
            I => \pid_alt.error_filt_prevZ0Z_8\
        );

    \I__10802\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45519\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__45519\,
            I => \N__45516\
        );

    \I__10800\ : Span4Mux_v
    port map (
            O => \N__45516\,
            I => \N__45513\
        );

    \I__10799\ : Span4Mux_h
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__10798\ : Span4Mux_h
    port map (
            O => \N__45510\,
            I => \N__45507\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__45507\,
            I => \N__45504\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__45504\,
            I => \N__45501\
        );

    \I__10795\ : Span4Mux_h
    port map (
            O => \N__45501\,
            I => \N__45498\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__45498\,
            I => \pid_alt.O_8\
        );

    \I__10793\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45490\
        );

    \I__10792\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45485\
        );

    \I__10791\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45485\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__45490\,
            I => \N__45482\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__45485\,
            I => \N__45479\
        );

    \I__10788\ : Span4Mux_v
    port map (
            O => \N__45482\,
            I => \N__45476\
        );

    \I__10787\ : Span4Mux_v
    port map (
            O => \N__45479\,
            I => \N__45473\
        );

    \I__10786\ : Sp12to4
    port map (
            O => \N__45476\,
            I => \N__45468\
        );

    \I__10785\ : Sp12to4
    port map (
            O => \N__45473\,
            I => \N__45468\
        );

    \I__10784\ : Span12Mux_h
    port map (
            O => \N__45468\,
            I => \N__45465\
        );

    \I__10783\ : Odrv12
    port map (
            O => \N__45465\,
            I => \pid_alt.error_d_regZ0Z_4\
        );

    \I__10782\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45459\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__45459\,
            I => \N__45456\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__45456\,
            I => \N__45453\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__45453\,
            I => \N__45449\
        );

    \I__10778\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45446\
        );

    \I__10777\ : Sp12to4
    port map (
            O => \N__45449\,
            I => \N__45443\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__45446\,
            I => \N__45440\
        );

    \I__10775\ : Span12Mux_h
    port map (
            O => \N__45443\,
            I => \N__45437\
        );

    \I__10774\ : Span4Mux_s1_h
    port map (
            O => \N__45440\,
            I => \N__45434\
        );

    \I__10773\ : Odrv12
    port map (
            O => \N__45437\,
            I => \pid_alt.error_filt_1\
        );

    \I__10772\ : Odrv4
    port map (
            O => \N__45434\,
            I => \pid_alt.error_filt_1\
        );

    \I__10771\ : InMux
    port map (
            O => \N__45429\,
            I => \N__45426\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__45426\,
            I => \N__45423\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__45423\,
            I => \pid_alt.error_filt_prevZ0Z_1\
        );

    \I__10768\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45417\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__45417\,
            I => \N__45414\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__45411\,
            I => \pid_alt.O_0_9\
        );

    \I__10764\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45405\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__45405\,
            I => \N__45402\
        );

    \I__10762\ : Span12Mux_h
    port map (
            O => \N__45402\,
            I => \N__45399\
        );

    \I__10761\ : Odrv12
    port map (
            O => \N__45399\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__10758\ : Span4Mux_v
    port map (
            O => \N__45390\,
            I => \N__45387\
        );

    \I__10757\ : Odrv4
    port map (
            O => \N__45387\,
            I => \pid_alt.O_0_12\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__45384\,
            I => \N__45381\
        );

    \I__10755\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45378\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__45378\,
            I => \N__45375\
        );

    \I__10753\ : Span4Mux_h
    port map (
            O => \N__45375\,
            I => \N__45372\
        );

    \I__10752\ : Span4Mux_h
    port map (
            O => \N__45372\,
            I => \N__45369\
        );

    \I__10751\ : Odrv4
    port map (
            O => \N__45369\,
            I => \pid_alt.error_i_regZ0Z_8\
        );

    \I__10750\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45363\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__45363\,
            I => \N__45359\
        );

    \I__10748\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45355\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__45359\,
            I => \N__45352\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45358\,
            I => \N__45347\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__45355\,
            I => \N__45344\
        );

    \I__10744\ : Span4Mux_h
    port map (
            O => \N__45352\,
            I => \N__45341\
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__45351\,
            I => \N__45338\
        );

    \I__10742\ : InMux
    port map (
            O => \N__45350\,
            I => \N__45335\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__45347\,
            I => \N__45332\
        );

    \I__10740\ : Span4Mux_v
    port map (
            O => \N__45344\,
            I => \N__45327\
        );

    \I__10739\ : Span4Mux_h
    port map (
            O => \N__45341\,
            I => \N__45324\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45321\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__45335\,
            I => \N__45318\
        );

    \I__10736\ : Span4Mux_v
    port map (
            O => \N__45332\,
            I => \N__45315\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45331\,
            I => \N__45310\
        );

    \I__10734\ : InMux
    port map (
            O => \N__45330\,
            I => \N__45307\
        );

    \I__10733\ : Span4Mux_h
    port map (
            O => \N__45327\,
            I => \N__45302\
        );

    \I__10732\ : Span4Mux_v
    port map (
            O => \N__45324\,
            I => \N__45302\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45321\,
            I => \N__45299\
        );

    \I__10730\ : Span4Mux_v
    port map (
            O => \N__45318\,
            I => \N__45293\
        );

    \I__10729\ : Span4Mux_v
    port map (
            O => \N__45315\,
            I => \N__45290\
        );

    \I__10728\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45287\
        );

    \I__10727\ : InMux
    port map (
            O => \N__45313\,
            I => \N__45284\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45275\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__45307\,
            I => \N__45275\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__45302\,
            I => \N__45275\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__45299\,
            I => \N__45275\
        );

    \I__10722\ : InMux
    port map (
            O => \N__45298\,
            I => \N__45271\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45268\
        );

    \I__10720\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45265\
        );

    \I__10719\ : Span4Mux_h
    port map (
            O => \N__45293\,
            I => \N__45260\
        );

    \I__10718\ : Span4Mux_v
    port map (
            O => \N__45290\,
            I => \N__45260\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__45287\,
            I => \N__45253\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__45284\,
            I => \N__45253\
        );

    \I__10715\ : Span4Mux_v
    port map (
            O => \N__45275\,
            I => \N__45253\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45274\,
            I => \N__45250\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__45271\,
            I => uart_pc_data_4
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45268\,
            I => uart_pc_data_4
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__45265\,
            I => uart_pc_data_4
        );

    \I__10710\ : Odrv4
    port map (
            O => \N__45260\,
            I => uart_pc_data_4
        );

    \I__10709\ : Odrv4
    port map (
            O => \N__45253\,
            I => uart_pc_data_4
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__45250\,
            I => uart_pc_data_4
        );

    \I__10707\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45234\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__45234\,
            I => \N__45231\
        );

    \I__10705\ : Span4Mux_s3_h
    port map (
            O => \N__45231\,
            I => \N__45228\
        );

    \I__10704\ : Odrv4
    port map (
            O => \N__45228\,
            I => alt_ki_4
        );

    \I__10703\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45221\
        );

    \I__10702\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45218\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__45221\,
            I => \N__45215\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__45218\,
            I => \N__45208\
        );

    \I__10699\ : Span4Mux_h
    port map (
            O => \N__45215\,
            I => \N__45205\
        );

    \I__10698\ : InMux
    port map (
            O => \N__45214\,
            I => \N__45201\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45213\,
            I => \N__45197\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45194\
        );

    \I__10695\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45191\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__45208\,
            I => \N__45187\
        );

    \I__10693\ : Span4Mux_h
    port map (
            O => \N__45205\,
            I => \N__45183\
        );

    \I__10692\ : InMux
    port map (
            O => \N__45204\,
            I => \N__45180\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__45201\,
            I => \N__45177\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45200\,
            I => \N__45173\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__45168\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45194\,
            I => \N__45168\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45165\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45162\
        );

    \I__10685\ : Sp12to4
    port map (
            O => \N__45187\,
            I => \N__45158\
        );

    \I__10684\ : InMux
    port map (
            O => \N__45186\,
            I => \N__45155\
        );

    \I__10683\ : Span4Mux_v
    port map (
            O => \N__45183\,
            I => \N__45150\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__45180\,
            I => \N__45150\
        );

    \I__10681\ : Span4Mux_h
    port map (
            O => \N__45177\,
            I => \N__45147\
        );

    \I__10680\ : InMux
    port map (
            O => \N__45176\,
            I => \N__45144\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45173\,
            I => \N__45141\
        );

    \I__10678\ : Span4Mux_v
    port map (
            O => \N__45168\,
            I => \N__45134\
        );

    \I__10677\ : Span4Mux_h
    port map (
            O => \N__45165\,
            I => \N__45134\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45134\
        );

    \I__10675\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45131\
        );

    \I__10674\ : Span12Mux_v
    port map (
            O => \N__45158\,
            I => \N__45127\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45124\
        );

    \I__10672\ : Span4Mux_h
    port map (
            O => \N__45150\,
            I => \N__45121\
        );

    \I__10671\ : Span4Mux_v
    port map (
            O => \N__45147\,
            I => \N__45118\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__45144\,
            I => \N__45115\
        );

    \I__10669\ : Span12Mux_h
    port map (
            O => \N__45141\,
            I => \N__45112\
        );

    \I__10668\ : Span4Mux_v
    port map (
            O => \N__45134\,
            I => \N__45109\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__45131\,
            I => \N__45106\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45103\
        );

    \I__10665\ : Span12Mux_h
    port map (
            O => \N__45127\,
            I => \N__45096\
        );

    \I__10664\ : Span12Mux_h
    port map (
            O => \N__45124\,
            I => \N__45096\
        );

    \I__10663\ : Sp12to4
    port map (
            O => \N__45121\,
            I => \N__45096\
        );

    \I__10662\ : Span4Mux_v
    port map (
            O => \N__45118\,
            I => \N__45091\
        );

    \I__10661\ : Span4Mux_h
    port map (
            O => \N__45115\,
            I => \N__45091\
        );

    \I__10660\ : Odrv12
    port map (
            O => \N__45112\,
            I => uart_pc_data_1
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__45109\,
            I => uart_pc_data_1
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__45106\,
            I => uart_pc_data_1
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__45103\,
            I => uart_pc_data_1
        );

    \I__10656\ : Odrv12
    port map (
            O => \N__45096\,
            I => uart_pc_data_1
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__45091\,
            I => uart_pc_data_1
        );

    \I__10654\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45075\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__10652\ : Span4Mux_v
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__45069\,
            I => alt_ki_1
        );

    \I__10650\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__45063\,
            I => \N__45060\
        );

    \I__10648\ : Span4Mux_h
    port map (
            O => \N__45060\,
            I => \N__45057\
        );

    \I__10647\ : Span4Mux_h
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10645\ : Span4Mux_h
    port map (
            O => \N__45051\,
            I => \N__45047\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45050\,
            I => \N__45044\
        );

    \I__10643\ : Span4Mux_h
    port map (
            O => \N__45047\,
            I => \N__45041\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__45044\,
            I => \N__45038\
        );

    \I__10641\ : Span4Mux_h
    port map (
            O => \N__45041\,
            I => \N__45033\
        );

    \I__10640\ : Span4Mux_v
    port map (
            O => \N__45038\,
            I => \N__45033\
        );

    \I__10639\ : Span4Mux_v
    port map (
            O => \N__45033\,
            I => \N__45030\
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__45030\,
            I => \pid_alt.error_filt_19\
        );

    \I__10637\ : InMux
    port map (
            O => \N__45027\,
            I => \N__45024\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__45024\,
            I => \N__45021\
        );

    \I__10635\ : Span4Mux_s2_h
    port map (
            O => \N__45021\,
            I => \N__45018\
        );

    \I__10634\ : Odrv4
    port map (
            O => \N__45018\,
            I => \pid_alt.error_filt_prevZ0Z_19\
        );

    \I__10633\ : InMux
    port map (
            O => \N__45015\,
            I => \N__45009\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45014\,
            I => \N__45006\
        );

    \I__10631\ : InMux
    port map (
            O => \N__45013\,
            I => \N__45002\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45012\,
            I => \N__44998\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__45009\,
            I => \N__44995\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__45006\,
            I => \N__44992\
        );

    \I__10627\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44989\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__45002\,
            I => \N__44985\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44979\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__44998\,
            I => \N__44976\
        );

    \I__10623\ : Span4Mux_v
    port map (
            O => \N__44995\,
            I => \N__44973\
        );

    \I__10622\ : Span4Mux_h
    port map (
            O => \N__44992\,
            I => \N__44970\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44967\
        );

    \I__10620\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44964\
        );

    \I__10619\ : Span4Mux_v
    port map (
            O => \N__44985\,
            I => \N__44961\
        );

    \I__10618\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44958\
        );

    \I__10617\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44955\
        );

    \I__10616\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44950\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__44979\,
            I => \N__44947\
        );

    \I__10614\ : Sp12to4
    port map (
            O => \N__44976\,
            I => \N__44941\
        );

    \I__10613\ : Sp12to4
    port map (
            O => \N__44973\,
            I => \N__44941\
        );

    \I__10612\ : Sp12to4
    port map (
            O => \N__44970\,
            I => \N__44934\
        );

    \I__10611\ : Sp12to4
    port map (
            O => \N__44967\,
            I => \N__44934\
        );

    \I__10610\ : LocalMux
    port map (
            O => \N__44964\,
            I => \N__44934\
        );

    \I__10609\ : Sp12to4
    port map (
            O => \N__44961\,
            I => \N__44931\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__44958\,
            I => \N__44926\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__44955\,
            I => \N__44926\
        );

    \I__10606\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44923\
        );

    \I__10605\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44920\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__44950\,
            I => \N__44915\
        );

    \I__10603\ : Span4Mux_h
    port map (
            O => \N__44947\,
            I => \N__44915\
        );

    \I__10602\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44911\
        );

    \I__10601\ : Span12Mux_v
    port map (
            O => \N__44941\,
            I => \N__44908\
        );

    \I__10600\ : Span12Mux_v
    port map (
            O => \N__44934\,
            I => \N__44903\
        );

    \I__10599\ : Span12Mux_v
    port map (
            O => \N__44931\,
            I => \N__44903\
        );

    \I__10598\ : Span4Mux_v
    port map (
            O => \N__44926\,
            I => \N__44898\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__44923\,
            I => \N__44898\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__44920\,
            I => \N__44893\
        );

    \I__10595\ : Span4Mux_v
    port map (
            O => \N__44915\,
            I => \N__44893\
        );

    \I__10594\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44890\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__44911\,
            I => uart_pc_data_7
        );

    \I__10592\ : Odrv12
    port map (
            O => \N__44908\,
            I => uart_pc_data_7
        );

    \I__10591\ : Odrv12
    port map (
            O => \N__44903\,
            I => uart_pc_data_7
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__44898\,
            I => uart_pc_data_7
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__44893\,
            I => uart_pc_data_7
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__44890\,
            I => uart_pc_data_7
        );

    \I__10587\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44874\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__44874\,
            I => \N__44871\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__44871\,
            I => \N__44868\
        );

    \I__10584\ : Odrv4
    port map (
            O => \N__44868\,
            I => alt_ki_7
        );

    \I__10583\ : CEMux
    port map (
            O => \N__44865\,
            I => \N__44861\
        );

    \I__10582\ : CEMux
    port map (
            O => \N__44864\,
            I => \N__44857\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__44861\,
            I => \N__44853\
        );

    \I__10580\ : CEMux
    port map (
            O => \N__44860\,
            I => \N__44850\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__44857\,
            I => \N__44846\
        );

    \I__10578\ : CEMux
    port map (
            O => \N__44856\,
            I => \N__44843\
        );

    \I__10577\ : Span4Mux_v
    port map (
            O => \N__44853\,
            I => \N__44838\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__44850\,
            I => \N__44838\
        );

    \I__10575\ : CEMux
    port map (
            O => \N__44849\,
            I => \N__44835\
        );

    \I__10574\ : Span4Mux_v
    port map (
            O => \N__44846\,
            I => \N__44832\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__44843\,
            I => \N__44829\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__44838\,
            I => \N__44825\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__44835\,
            I => \N__44822\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__44832\,
            I => \N__44816\
        );

    \I__10569\ : Span4Mux_h
    port map (
            O => \N__44829\,
            I => \N__44816\
        );

    \I__10568\ : CEMux
    port map (
            O => \N__44828\,
            I => \N__44813\
        );

    \I__10567\ : Span4Mux_h
    port map (
            O => \N__44825\,
            I => \N__44808\
        );

    \I__10566\ : Span4Mux_v
    port map (
            O => \N__44822\,
            I => \N__44808\
        );

    \I__10565\ : CEMux
    port map (
            O => \N__44821\,
            I => \N__44805\
        );

    \I__10564\ : Span4Mux_h
    port map (
            O => \N__44816\,
            I => \N__44800\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__44813\,
            I => \N__44800\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__44808\,
            I => \N__44795\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44795\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__44800\,
            I => \N__44792\
        );

    \I__10559\ : Span4Mux_h
    port map (
            O => \N__44795\,
            I => \N__44789\
        );

    \I__10558\ : Sp12to4
    port map (
            O => \N__44792\,
            I => \N__44786\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__44789\,
            I => \N__44783\
        );

    \I__10556\ : Span12Mux_h
    port map (
            O => \N__44786\,
            I => \N__44780\
        );

    \I__10555\ : Span4Mux_v
    port map (
            O => \N__44783\,
            I => \N__44777\
        );

    \I__10554\ : Odrv12
    port map (
            O => \N__44780\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__44777\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__10552\ : InMux
    port map (
            O => \N__44772\,
            I => \N__44769\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__44769\,
            I => \N__44766\
        );

    \I__10550\ : Span4Mux_h
    port map (
            O => \N__44766\,
            I => \N__44763\
        );

    \I__10549\ : Odrv4
    port map (
            O => \N__44763\,
            I => \pid_alt.O_0_14\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__44760\,
            I => \N__44757\
        );

    \I__10547\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44754\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__44754\,
            I => \N__44751\
        );

    \I__10545\ : Span4Mux_v
    port map (
            O => \N__44751\,
            I => \N__44748\
        );

    \I__10544\ : Span4Mux_h
    port map (
            O => \N__44748\,
            I => \N__44745\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__44745\,
            I => \N__44742\
        );

    \I__10542\ : Odrv4
    port map (
            O => \N__44742\,
            I => \pid_alt.error_i_regZ0Z_10\
        );

    \I__10541\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44736\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__44736\,
            I => \N__44733\
        );

    \I__10539\ : Span4Mux_h
    port map (
            O => \N__44733\,
            I => \N__44730\
        );

    \I__10538\ : Odrv4
    port map (
            O => \N__44730\,
            I => \pid_alt.O_15\
        );

    \I__10537\ : CascadeMux
    port map (
            O => \N__44727\,
            I => \N__44724\
        );

    \I__10536\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44721\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__44721\,
            I => \N__44718\
        );

    \I__10534\ : Span4Mux_v
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__10533\ : Span4Mux_h
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__10532\ : Span4Mux_h
    port map (
            O => \N__44712\,
            I => \N__44709\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__44709\,
            I => \pid_alt.error_i_regZ0Z_11\
        );

    \I__10530\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44703\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__44703\,
            I => \N__44700\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__44700\,
            I => \N__44697\
        );

    \I__10527\ : Odrv4
    port map (
            O => \N__44697\,
            I => \pid_alt.O_16\
        );

    \I__10526\ : CascadeMux
    port map (
            O => \N__44694\,
            I => \N__44691\
        );

    \I__10525\ : InMux
    port map (
            O => \N__44691\,
            I => \N__44688\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__44688\,
            I => \N__44685\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__10522\ : Span4Mux_h
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__10521\ : Span4Mux_h
    port map (
            O => \N__44679\,
            I => \N__44676\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__44676\,
            I => \pid_alt.error_i_regZ0Z_12\
        );

    \I__10519\ : InMux
    port map (
            O => \N__44673\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__10518\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44667\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__44667\,
            I => \N__44662\
        );

    \I__10516\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44656\
        );

    \I__10515\ : InMux
    port map (
            O => \N__44665\,
            I => \N__44656\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__44662\,
            I => \N__44653\
        );

    \I__10513\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44650\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__44656\,
            I => \N__44647\
        );

    \I__10511\ : Span4Mux_v
    port map (
            O => \N__44653\,
            I => \N__44642\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__44650\,
            I => \N__44642\
        );

    \I__10509\ : Span4Mux_v
    port map (
            O => \N__44647\,
            I => \N__44639\
        );

    \I__10508\ : Odrv4
    port map (
            O => \N__44642\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__10507\ : Odrv4
    port map (
            O => \N__44639\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__10506\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44631\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__44631\,
            I => \N__44628\
        );

    \I__10504\ : Odrv4
    port map (
            O => \N__44628\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__10503\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44622\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__44622\,
            I => \N__44617\
        );

    \I__10501\ : InMux
    port map (
            O => \N__44621\,
            I => \N__44614\
        );

    \I__10500\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44611\
        );

    \I__10499\ : Span4Mux_h
    port map (
            O => \N__44617\,
            I => \N__44608\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__44614\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__44611\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__10496\ : Odrv4
    port map (
            O => \N__44608\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__10495\ : CascadeMux
    port map (
            O => \N__44601\,
            I => \N__44598\
        );

    \I__10494\ : InMux
    port map (
            O => \N__44598\,
            I => \N__44595\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__44595\,
            I => \N__44592\
        );

    \I__10492\ : Odrv4
    port map (
            O => \N__44592\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__10491\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44586\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__44586\,
            I => \N__44581\
        );

    \I__10489\ : InMux
    port map (
            O => \N__44585\,
            I => \N__44578\
        );

    \I__10488\ : InMux
    port map (
            O => \N__44584\,
            I => \N__44575\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__44581\,
            I => \N__44572\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__44578\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__44575\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__44572\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__44565\,
            I => \N__44562\
        );

    \I__10482\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44559\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__44559\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__10480\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44553\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__44553\,
            I => \N__44549\
        );

    \I__10478\ : CascadeMux
    port map (
            O => \N__44552\,
            I => \N__44545\
        );

    \I__10477\ : Span4Mux_h
    port map (
            O => \N__44549\,
            I => \N__44542\
        );

    \I__10476\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44532\
        );

    \I__10475\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44532\
        );

    \I__10474\ : Span4Mux_h
    port map (
            O => \N__44542\,
            I => \N__44529\
        );

    \I__10473\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44526\
        );

    \I__10472\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44523\
        );

    \I__10471\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44520\
        );

    \I__10470\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44515\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44515\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__44532\,
            I => \N__44512\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__44529\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__44526\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__44523\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__44520\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__44515\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10462\ : Odrv4
    port map (
            O => \N__44512\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__10461\ : CascadeMux
    port map (
            O => \N__44499\,
            I => \N__44496\
        );

    \I__10460\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44492\
        );

    \I__10459\ : CascadeMux
    port map (
            O => \N__44495\,
            I => \N__44489\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44486\
        );

    \I__10457\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44482\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__44486\,
            I => \N__44479\
        );

    \I__10455\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44476\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__44482\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__10453\ : Odrv4
    port map (
            O => \N__44479\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44476\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44465\
        );

    \I__10450\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44462\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__44465\,
            I => \N__44458\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44455\
        );

    \I__10447\ : InMux
    port map (
            O => \N__44461\,
            I => \N__44452\
        );

    \I__10446\ : Span4Mux_v
    port map (
            O => \N__44458\,
            I => \N__44448\
        );

    \I__10445\ : Span4Mux_v
    port map (
            O => \N__44455\,
            I => \N__44445\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__44452\,
            I => \N__44442\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44451\,
            I => \N__44439\
        );

    \I__10442\ : Span4Mux_h
    port map (
            O => \N__44448\,
            I => \N__44436\
        );

    \I__10441\ : Span4Mux_h
    port map (
            O => \N__44445\,
            I => \N__44429\
        );

    \I__10440\ : Span4Mux_v
    port map (
            O => \N__44442\,
            I => \N__44429\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__44439\,
            I => \N__44429\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__44436\,
            I => \uart_drone.N_152\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__44429\,
            I => \uart_drone.N_152\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44415\
        );

    \I__10435\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44415\
        );

    \I__10434\ : InMux
    port map (
            O => \N__44422\,
            I => \N__44410\
        );

    \I__10433\ : InMux
    port map (
            O => \N__44421\,
            I => \N__44410\
        );

    \I__10432\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44407\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44398\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__44410\,
            I => \N__44398\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__44407\,
            I => \N__44398\
        );

    \I__10428\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44393\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44405\,
            I => \N__44393\
        );

    \I__10426\ : Span4Mux_v
    port map (
            O => \N__44398\,
            I => \N__44386\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__44393\,
            I => \N__44386\
        );

    \I__10424\ : InMux
    port map (
            O => \N__44392\,
            I => \N__44383\
        );

    \I__10423\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44379\
        );

    \I__10422\ : Span4Mux_h
    port map (
            O => \N__44386\,
            I => \N__44375\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__44383\,
            I => \N__44372\
        );

    \I__10420\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44369\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44366\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44363\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__44375\,
            I => \N__44360\
        );

    \I__10416\ : Span4Mux_v
    port map (
            O => \N__44372\,
            I => \N__44355\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44369\,
            I => \N__44355\
        );

    \I__10414\ : Span12Mux_h
    port map (
            O => \N__44366\,
            I => \N__44352\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__44363\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__10412\ : Odrv4
    port map (
            O => \N__44360\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__10411\ : Odrv4
    port map (
            O => \N__44355\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__10410\ : Odrv12
    port map (
            O => \N__44352\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__10409\ : InMux
    port map (
            O => \N__44343\,
            I => \N__44340\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__44337\,
            I => \N__44334\
        );

    \I__10406\ : Span4Mux_h
    port map (
            O => \N__44334\,
            I => \N__44331\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__44331\,
            I => \N__44327\
        );

    \I__10404\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44324\
        );

    \I__10403\ : Span4Mux_h
    port map (
            O => \N__44327\,
            I => \N__44321\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44324\,
            I => \N__44318\
        );

    \I__10401\ : Span4Mux_h
    port map (
            O => \N__44321\,
            I => \N__44313\
        );

    \I__10400\ : Span4Mux_v
    port map (
            O => \N__44318\,
            I => \N__44313\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__44313\,
            I => \N__44310\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__44310\,
            I => \pid_alt.error_filt_21\
        );

    \I__10397\ : InMux
    port map (
            O => \N__44307\,
            I => \N__44304\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__44304\,
            I => \N__44301\
        );

    \I__10395\ : Span4Mux_s0_h
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__10394\ : Span4Mux_h
    port map (
            O => \N__44298\,
            I => \N__44295\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__44295\,
            I => \pid_alt.error_filt_prevZ0Z_21\
        );

    \I__10392\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44287\
        );

    \I__10391\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44284\
        );

    \I__10390\ : InMux
    port map (
            O => \N__44290\,
            I => \N__44280\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44287\,
            I => \N__44275\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__44284\,
            I => \N__44275\
        );

    \I__10387\ : InMux
    port map (
            O => \N__44283\,
            I => \N__44272\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__44280\,
            I => \N__44267\
        );

    \I__10385\ : Span4Mux_v
    port map (
            O => \N__44275\,
            I => \N__44264\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__44272\,
            I => \N__44259\
        );

    \I__10383\ : CascadeMux
    port map (
            O => \N__44271\,
            I => \N__44255\
        );

    \I__10382\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44251\
        );

    \I__10381\ : Span4Mux_v
    port map (
            O => \N__44267\,
            I => \N__44244\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__44264\,
            I => \N__44244\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44263\,
            I => \N__44241\
        );

    \I__10378\ : InMux
    port map (
            O => \N__44262\,
            I => \N__44237\
        );

    \I__10377\ : Span4Mux_v
    port map (
            O => \N__44259\,
            I => \N__44234\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44258\,
            I => \N__44227\
        );

    \I__10375\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44227\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44254\,
            I => \N__44227\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__44251\,
            I => \N__44224\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44221\
        );

    \I__10371\ : InMux
    port map (
            O => \N__44249\,
            I => \N__44218\
        );

    \I__10370\ : Span4Mux_v
    port map (
            O => \N__44244\,
            I => \N__44213\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__44241\,
            I => \N__44213\
        );

    \I__10368\ : InMux
    port map (
            O => \N__44240\,
            I => \N__44210\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__44237\,
            I => \N__44207\
        );

    \I__10366\ : Sp12to4
    port map (
            O => \N__44234\,
            I => \N__44202\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44199\
        );

    \I__10364\ : Span4Mux_v
    port map (
            O => \N__44224\,
            I => \N__44190\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__44221\,
            I => \N__44190\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44218\,
            I => \N__44190\
        );

    \I__10361\ : Span4Mux_h
    port map (
            O => \N__44213\,
            I => \N__44190\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__44210\,
            I => \N__44187\
        );

    \I__10359\ : Span4Mux_h
    port map (
            O => \N__44207\,
            I => \N__44184\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44206\,
            I => \N__44181\
        );

    \I__10357\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44178\
        );

    \I__10356\ : Span12Mux_v
    port map (
            O => \N__44202\,
            I => \N__44175\
        );

    \I__10355\ : Span4Mux_h
    port map (
            O => \N__44199\,
            I => \N__44172\
        );

    \I__10354\ : Span4Mux_v
    port map (
            O => \N__44190\,
            I => \N__44169\
        );

    \I__10353\ : Odrv12
    port map (
            O => \N__44187\,
            I => uart_pc_data_5
        );

    \I__10352\ : Odrv4
    port map (
            O => \N__44184\,
            I => uart_pc_data_5
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__44181\,
            I => uart_pc_data_5
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__44178\,
            I => uart_pc_data_5
        );

    \I__10349\ : Odrv12
    port map (
            O => \N__44175\,
            I => uart_pc_data_5
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__44172\,
            I => uart_pc_data_5
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__44169\,
            I => uart_pc_data_5
        );

    \I__10346\ : InMux
    port map (
            O => \N__44154\,
            I => \N__44151\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__44151\,
            I => \N__44148\
        );

    \I__10344\ : Span4Mux_s0_h
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__10343\ : Span4Mux_h
    port map (
            O => \N__44145\,
            I => \N__44142\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__44142\,
            I => alt_ki_5
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__44139\,
            I => \N__44132\
        );

    \I__10340\ : CascadeMux
    port map (
            O => \N__44138\,
            I => \N__44129\
        );

    \I__10339\ : CascadeMux
    port map (
            O => \N__44137\,
            I => \N__44119\
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__44136\,
            I => \N__44113\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__44135\,
            I => \N__44093\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44132\,
            I => \N__44060\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44129\,
            I => \N__44060\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44057\
        );

    \I__10333\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44052\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44052\
        );

    \I__10331\ : InMux
    port map (
            O => \N__44125\,
            I => \N__44049\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44046\
        );

    \I__10329\ : InMux
    port map (
            O => \N__44123\,
            I => \N__44043\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44122\,
            I => \N__44040\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44037\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44034\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44117\,
            I => \N__44031\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44116\,
            I => \N__44022\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44113\,
            I => \N__44022\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44022\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44022\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44110\,
            I => \N__44019\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44109\,
            I => \N__44014\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44014\
        );

    \I__10317\ : InMux
    port map (
            O => \N__44107\,
            I => \N__44009\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44106\,
            I => \N__44009\
        );

    \I__10315\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44004\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44104\,
            I => \N__44004\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44103\,
            I => \N__43999\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44102\,
            I => \N__43999\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44101\,
            I => \N__43996\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44100\,
            I => \N__43993\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44099\,
            I => \N__43990\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44098\,
            I => \N__43983\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44097\,
            I => \N__43983\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44096\,
            I => \N__43983\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44093\,
            I => \N__43980\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44092\,
            I => \N__43977\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44091\,
            I => \N__43974\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44090\,
            I => \N__43971\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44089\,
            I => \N__43968\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44088\,
            I => \N__43965\
        );

    \I__10299\ : InMux
    port map (
            O => \N__44087\,
            I => \N__43960\
        );

    \I__10298\ : InMux
    port map (
            O => \N__44086\,
            I => \N__43960\
        );

    \I__10297\ : InMux
    port map (
            O => \N__44085\,
            I => \N__43957\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44084\,
            I => \N__43954\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44083\,
            I => \N__43951\
        );

    \I__10294\ : InMux
    port map (
            O => \N__44082\,
            I => \N__43948\
        );

    \I__10293\ : InMux
    port map (
            O => \N__44081\,
            I => \N__43941\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44080\,
            I => \N__43941\
        );

    \I__10291\ : InMux
    port map (
            O => \N__44079\,
            I => \N__43941\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44078\,
            I => \N__43938\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44077\,
            I => \N__43933\
        );

    \I__10288\ : InMux
    port map (
            O => \N__44076\,
            I => \N__43933\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44075\,
            I => \N__43930\
        );

    \I__10286\ : InMux
    port map (
            O => \N__44074\,
            I => \N__43927\
        );

    \I__10285\ : InMux
    port map (
            O => \N__44073\,
            I => \N__43922\
        );

    \I__10284\ : InMux
    port map (
            O => \N__44072\,
            I => \N__43922\
        );

    \I__10283\ : InMux
    port map (
            O => \N__44071\,
            I => \N__43919\
        );

    \I__10282\ : InMux
    port map (
            O => \N__44070\,
            I => \N__43916\
        );

    \I__10281\ : InMux
    port map (
            O => \N__44069\,
            I => \N__43913\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44068\,
            I => \N__43908\
        );

    \I__10279\ : InMux
    port map (
            O => \N__44067\,
            I => \N__43908\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44066\,
            I => \N__43905\
        );

    \I__10277\ : InMux
    port map (
            O => \N__44065\,
            I => \N__43902\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__43796\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__44057\,
            I => \N__43793\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__43790\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__43787\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__44046\,
            I => \N__43784\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__43781\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__44040\,
            I => \N__43778\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__44037\,
            I => \N__43775\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__43772\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__44031\,
            I => \N__43769\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44022\,
            I => \N__43766\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__44019\,
            I => \N__43763\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44014\,
            I => \N__43760\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44009\,
            I => \N__43757\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44004\,
            I => \N__43754\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__43999\,
            I => \N__43751\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__43996\,
            I => \N__43748\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__43993\,
            I => \N__43745\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__43990\,
            I => \N__43742\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43739\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__43980\,
            I => \N__43736\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__43977\,
            I => \N__43733\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43730\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__43971\,
            I => \N__43727\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__43968\,
            I => \N__43724\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__43965\,
            I => \N__43721\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__43960\,
            I => \N__43718\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__43957\,
            I => \N__43715\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__43954\,
            I => \N__43712\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__43951\,
            I => \N__43709\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43706\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__43941\,
            I => \N__43703\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__43938\,
            I => \N__43700\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43697\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__43930\,
            I => \N__43694\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__43927\,
            I => \N__43691\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__43922\,
            I => \N__43688\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__43919\,
            I => \N__43685\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__43916\,
            I => \N__43682\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43679\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__43908\,
            I => \N__43676\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__43905\,
            I => \N__43673\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__43902\,
            I => \N__43670\
        );

    \I__10233\ : SRMux
    port map (
            O => \N__43901\,
            I => \N__43377\
        );

    \I__10232\ : SRMux
    port map (
            O => \N__43900\,
            I => \N__43377\
        );

    \I__10231\ : SRMux
    port map (
            O => \N__43899\,
            I => \N__43377\
        );

    \I__10230\ : SRMux
    port map (
            O => \N__43898\,
            I => \N__43377\
        );

    \I__10229\ : SRMux
    port map (
            O => \N__43897\,
            I => \N__43377\
        );

    \I__10228\ : SRMux
    port map (
            O => \N__43896\,
            I => \N__43377\
        );

    \I__10227\ : SRMux
    port map (
            O => \N__43895\,
            I => \N__43377\
        );

    \I__10226\ : SRMux
    port map (
            O => \N__43894\,
            I => \N__43377\
        );

    \I__10225\ : SRMux
    port map (
            O => \N__43893\,
            I => \N__43377\
        );

    \I__10224\ : SRMux
    port map (
            O => \N__43892\,
            I => \N__43377\
        );

    \I__10223\ : SRMux
    port map (
            O => \N__43891\,
            I => \N__43377\
        );

    \I__10222\ : SRMux
    port map (
            O => \N__43890\,
            I => \N__43377\
        );

    \I__10221\ : SRMux
    port map (
            O => \N__43889\,
            I => \N__43377\
        );

    \I__10220\ : SRMux
    port map (
            O => \N__43888\,
            I => \N__43377\
        );

    \I__10219\ : SRMux
    port map (
            O => \N__43887\,
            I => \N__43377\
        );

    \I__10218\ : SRMux
    port map (
            O => \N__43886\,
            I => \N__43377\
        );

    \I__10217\ : SRMux
    port map (
            O => \N__43885\,
            I => \N__43377\
        );

    \I__10216\ : SRMux
    port map (
            O => \N__43884\,
            I => \N__43377\
        );

    \I__10215\ : SRMux
    port map (
            O => \N__43883\,
            I => \N__43377\
        );

    \I__10214\ : SRMux
    port map (
            O => \N__43882\,
            I => \N__43377\
        );

    \I__10213\ : SRMux
    port map (
            O => \N__43881\,
            I => \N__43377\
        );

    \I__10212\ : SRMux
    port map (
            O => \N__43880\,
            I => \N__43377\
        );

    \I__10211\ : SRMux
    port map (
            O => \N__43879\,
            I => \N__43377\
        );

    \I__10210\ : SRMux
    port map (
            O => \N__43878\,
            I => \N__43377\
        );

    \I__10209\ : SRMux
    port map (
            O => \N__43877\,
            I => \N__43377\
        );

    \I__10208\ : SRMux
    port map (
            O => \N__43876\,
            I => \N__43377\
        );

    \I__10207\ : SRMux
    port map (
            O => \N__43875\,
            I => \N__43377\
        );

    \I__10206\ : SRMux
    port map (
            O => \N__43874\,
            I => \N__43377\
        );

    \I__10205\ : SRMux
    port map (
            O => \N__43873\,
            I => \N__43377\
        );

    \I__10204\ : SRMux
    port map (
            O => \N__43872\,
            I => \N__43377\
        );

    \I__10203\ : SRMux
    port map (
            O => \N__43871\,
            I => \N__43377\
        );

    \I__10202\ : SRMux
    port map (
            O => \N__43870\,
            I => \N__43377\
        );

    \I__10201\ : SRMux
    port map (
            O => \N__43869\,
            I => \N__43377\
        );

    \I__10200\ : SRMux
    port map (
            O => \N__43868\,
            I => \N__43377\
        );

    \I__10199\ : SRMux
    port map (
            O => \N__43867\,
            I => \N__43377\
        );

    \I__10198\ : SRMux
    port map (
            O => \N__43866\,
            I => \N__43377\
        );

    \I__10197\ : SRMux
    port map (
            O => \N__43865\,
            I => \N__43377\
        );

    \I__10196\ : SRMux
    port map (
            O => \N__43864\,
            I => \N__43377\
        );

    \I__10195\ : SRMux
    port map (
            O => \N__43863\,
            I => \N__43377\
        );

    \I__10194\ : SRMux
    port map (
            O => \N__43862\,
            I => \N__43377\
        );

    \I__10193\ : SRMux
    port map (
            O => \N__43861\,
            I => \N__43377\
        );

    \I__10192\ : SRMux
    port map (
            O => \N__43860\,
            I => \N__43377\
        );

    \I__10191\ : SRMux
    port map (
            O => \N__43859\,
            I => \N__43377\
        );

    \I__10190\ : SRMux
    port map (
            O => \N__43858\,
            I => \N__43377\
        );

    \I__10189\ : SRMux
    port map (
            O => \N__43857\,
            I => \N__43377\
        );

    \I__10188\ : SRMux
    port map (
            O => \N__43856\,
            I => \N__43377\
        );

    \I__10187\ : SRMux
    port map (
            O => \N__43855\,
            I => \N__43377\
        );

    \I__10186\ : SRMux
    port map (
            O => \N__43854\,
            I => \N__43377\
        );

    \I__10185\ : SRMux
    port map (
            O => \N__43853\,
            I => \N__43377\
        );

    \I__10184\ : SRMux
    port map (
            O => \N__43852\,
            I => \N__43377\
        );

    \I__10183\ : SRMux
    port map (
            O => \N__43851\,
            I => \N__43377\
        );

    \I__10182\ : SRMux
    port map (
            O => \N__43850\,
            I => \N__43377\
        );

    \I__10181\ : SRMux
    port map (
            O => \N__43849\,
            I => \N__43377\
        );

    \I__10180\ : SRMux
    port map (
            O => \N__43848\,
            I => \N__43377\
        );

    \I__10179\ : SRMux
    port map (
            O => \N__43847\,
            I => \N__43377\
        );

    \I__10178\ : SRMux
    port map (
            O => \N__43846\,
            I => \N__43377\
        );

    \I__10177\ : SRMux
    port map (
            O => \N__43845\,
            I => \N__43377\
        );

    \I__10176\ : SRMux
    port map (
            O => \N__43844\,
            I => \N__43377\
        );

    \I__10175\ : SRMux
    port map (
            O => \N__43843\,
            I => \N__43377\
        );

    \I__10174\ : SRMux
    port map (
            O => \N__43842\,
            I => \N__43377\
        );

    \I__10173\ : SRMux
    port map (
            O => \N__43841\,
            I => \N__43377\
        );

    \I__10172\ : SRMux
    port map (
            O => \N__43840\,
            I => \N__43377\
        );

    \I__10171\ : SRMux
    port map (
            O => \N__43839\,
            I => \N__43377\
        );

    \I__10170\ : SRMux
    port map (
            O => \N__43838\,
            I => \N__43377\
        );

    \I__10169\ : SRMux
    port map (
            O => \N__43837\,
            I => \N__43377\
        );

    \I__10168\ : SRMux
    port map (
            O => \N__43836\,
            I => \N__43377\
        );

    \I__10167\ : SRMux
    port map (
            O => \N__43835\,
            I => \N__43377\
        );

    \I__10166\ : SRMux
    port map (
            O => \N__43834\,
            I => \N__43377\
        );

    \I__10165\ : SRMux
    port map (
            O => \N__43833\,
            I => \N__43377\
        );

    \I__10164\ : SRMux
    port map (
            O => \N__43832\,
            I => \N__43377\
        );

    \I__10163\ : SRMux
    port map (
            O => \N__43831\,
            I => \N__43377\
        );

    \I__10162\ : SRMux
    port map (
            O => \N__43830\,
            I => \N__43377\
        );

    \I__10161\ : SRMux
    port map (
            O => \N__43829\,
            I => \N__43377\
        );

    \I__10160\ : SRMux
    port map (
            O => \N__43828\,
            I => \N__43377\
        );

    \I__10159\ : SRMux
    port map (
            O => \N__43827\,
            I => \N__43377\
        );

    \I__10158\ : SRMux
    port map (
            O => \N__43826\,
            I => \N__43377\
        );

    \I__10157\ : SRMux
    port map (
            O => \N__43825\,
            I => \N__43377\
        );

    \I__10156\ : SRMux
    port map (
            O => \N__43824\,
            I => \N__43377\
        );

    \I__10155\ : SRMux
    port map (
            O => \N__43823\,
            I => \N__43377\
        );

    \I__10154\ : SRMux
    port map (
            O => \N__43822\,
            I => \N__43377\
        );

    \I__10153\ : SRMux
    port map (
            O => \N__43821\,
            I => \N__43377\
        );

    \I__10152\ : SRMux
    port map (
            O => \N__43820\,
            I => \N__43377\
        );

    \I__10151\ : SRMux
    port map (
            O => \N__43819\,
            I => \N__43377\
        );

    \I__10150\ : SRMux
    port map (
            O => \N__43818\,
            I => \N__43377\
        );

    \I__10149\ : SRMux
    port map (
            O => \N__43817\,
            I => \N__43377\
        );

    \I__10148\ : SRMux
    port map (
            O => \N__43816\,
            I => \N__43377\
        );

    \I__10147\ : SRMux
    port map (
            O => \N__43815\,
            I => \N__43377\
        );

    \I__10146\ : SRMux
    port map (
            O => \N__43814\,
            I => \N__43377\
        );

    \I__10145\ : SRMux
    port map (
            O => \N__43813\,
            I => \N__43377\
        );

    \I__10144\ : SRMux
    port map (
            O => \N__43812\,
            I => \N__43377\
        );

    \I__10143\ : SRMux
    port map (
            O => \N__43811\,
            I => \N__43377\
        );

    \I__10142\ : SRMux
    port map (
            O => \N__43810\,
            I => \N__43377\
        );

    \I__10141\ : SRMux
    port map (
            O => \N__43809\,
            I => \N__43377\
        );

    \I__10140\ : SRMux
    port map (
            O => \N__43808\,
            I => \N__43377\
        );

    \I__10139\ : SRMux
    port map (
            O => \N__43807\,
            I => \N__43377\
        );

    \I__10138\ : SRMux
    port map (
            O => \N__43806\,
            I => \N__43377\
        );

    \I__10137\ : SRMux
    port map (
            O => \N__43805\,
            I => \N__43377\
        );

    \I__10136\ : SRMux
    port map (
            O => \N__43804\,
            I => \N__43377\
        );

    \I__10135\ : SRMux
    port map (
            O => \N__43803\,
            I => \N__43377\
        );

    \I__10134\ : SRMux
    port map (
            O => \N__43802\,
            I => \N__43377\
        );

    \I__10133\ : SRMux
    port map (
            O => \N__43801\,
            I => \N__43377\
        );

    \I__10132\ : SRMux
    port map (
            O => \N__43800\,
            I => \N__43377\
        );

    \I__10131\ : SRMux
    port map (
            O => \N__43799\,
            I => \N__43377\
        );

    \I__10130\ : Glb2LocalMux
    port map (
            O => \N__43796\,
            I => \N__43377\
        );

    \I__10129\ : Glb2LocalMux
    port map (
            O => \N__43793\,
            I => \N__43377\
        );

    \I__10128\ : Glb2LocalMux
    port map (
            O => \N__43790\,
            I => \N__43377\
        );

    \I__10127\ : Glb2LocalMux
    port map (
            O => \N__43787\,
            I => \N__43377\
        );

    \I__10126\ : Glb2LocalMux
    port map (
            O => \N__43784\,
            I => \N__43377\
        );

    \I__10125\ : Glb2LocalMux
    port map (
            O => \N__43781\,
            I => \N__43377\
        );

    \I__10124\ : Glb2LocalMux
    port map (
            O => \N__43778\,
            I => \N__43377\
        );

    \I__10123\ : Glb2LocalMux
    port map (
            O => \N__43775\,
            I => \N__43377\
        );

    \I__10122\ : Glb2LocalMux
    port map (
            O => \N__43772\,
            I => \N__43377\
        );

    \I__10121\ : Glb2LocalMux
    port map (
            O => \N__43769\,
            I => \N__43377\
        );

    \I__10120\ : Glb2LocalMux
    port map (
            O => \N__43766\,
            I => \N__43377\
        );

    \I__10119\ : Glb2LocalMux
    port map (
            O => \N__43763\,
            I => \N__43377\
        );

    \I__10118\ : Glb2LocalMux
    port map (
            O => \N__43760\,
            I => \N__43377\
        );

    \I__10117\ : Glb2LocalMux
    port map (
            O => \N__43757\,
            I => \N__43377\
        );

    \I__10116\ : Glb2LocalMux
    port map (
            O => \N__43754\,
            I => \N__43377\
        );

    \I__10115\ : Glb2LocalMux
    port map (
            O => \N__43751\,
            I => \N__43377\
        );

    \I__10114\ : Glb2LocalMux
    port map (
            O => \N__43748\,
            I => \N__43377\
        );

    \I__10113\ : Glb2LocalMux
    port map (
            O => \N__43745\,
            I => \N__43377\
        );

    \I__10112\ : Glb2LocalMux
    port map (
            O => \N__43742\,
            I => \N__43377\
        );

    \I__10111\ : Glb2LocalMux
    port map (
            O => \N__43739\,
            I => \N__43377\
        );

    \I__10110\ : Glb2LocalMux
    port map (
            O => \N__43736\,
            I => \N__43377\
        );

    \I__10109\ : Glb2LocalMux
    port map (
            O => \N__43733\,
            I => \N__43377\
        );

    \I__10108\ : Glb2LocalMux
    port map (
            O => \N__43730\,
            I => \N__43377\
        );

    \I__10107\ : Glb2LocalMux
    port map (
            O => \N__43727\,
            I => \N__43377\
        );

    \I__10106\ : Glb2LocalMux
    port map (
            O => \N__43724\,
            I => \N__43377\
        );

    \I__10105\ : Glb2LocalMux
    port map (
            O => \N__43721\,
            I => \N__43377\
        );

    \I__10104\ : Glb2LocalMux
    port map (
            O => \N__43718\,
            I => \N__43377\
        );

    \I__10103\ : Glb2LocalMux
    port map (
            O => \N__43715\,
            I => \N__43377\
        );

    \I__10102\ : Glb2LocalMux
    port map (
            O => \N__43712\,
            I => \N__43377\
        );

    \I__10101\ : Glb2LocalMux
    port map (
            O => \N__43709\,
            I => \N__43377\
        );

    \I__10100\ : Glb2LocalMux
    port map (
            O => \N__43706\,
            I => \N__43377\
        );

    \I__10099\ : Glb2LocalMux
    port map (
            O => \N__43703\,
            I => \N__43377\
        );

    \I__10098\ : Glb2LocalMux
    port map (
            O => \N__43700\,
            I => \N__43377\
        );

    \I__10097\ : Glb2LocalMux
    port map (
            O => \N__43697\,
            I => \N__43377\
        );

    \I__10096\ : Glb2LocalMux
    port map (
            O => \N__43694\,
            I => \N__43377\
        );

    \I__10095\ : Glb2LocalMux
    port map (
            O => \N__43691\,
            I => \N__43377\
        );

    \I__10094\ : Glb2LocalMux
    port map (
            O => \N__43688\,
            I => \N__43377\
        );

    \I__10093\ : Glb2LocalMux
    port map (
            O => \N__43685\,
            I => \N__43377\
        );

    \I__10092\ : Glb2LocalMux
    port map (
            O => \N__43682\,
            I => \N__43377\
        );

    \I__10091\ : Glb2LocalMux
    port map (
            O => \N__43679\,
            I => \N__43377\
        );

    \I__10090\ : Glb2LocalMux
    port map (
            O => \N__43676\,
            I => \N__43377\
        );

    \I__10089\ : Glb2LocalMux
    port map (
            O => \N__43673\,
            I => \N__43377\
        );

    \I__10088\ : Glb2LocalMux
    port map (
            O => \N__43670\,
            I => \N__43377\
        );

    \I__10087\ : GlobalMux
    port map (
            O => \N__43377\,
            I => \N__43374\
        );

    \I__10086\ : gio2CtrlBuf
    port map (
            O => \N__43374\,
            I => reset_system_g
        );

    \I__10085\ : IoInMux
    port map (
            O => \N__43371\,
            I => \N__43368\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__43368\,
            I => \GB_BUFFER_reset_system_g_THRU_CO\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43361\
        );

    \I__10082\ : InMux
    port map (
            O => \N__43364\,
            I => \N__43358\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__43361\,
            I => \N__43355\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__43358\,
            I => \N__43350\
        );

    \I__10079\ : Span4Mux_v
    port map (
            O => \N__43355\,
            I => \N__43346\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43354\,
            I => \N__43343\
        );

    \I__10077\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43336\
        );

    \I__10076\ : Span4Mux_v
    port map (
            O => \N__43350\,
            I => \N__43333\
        );

    \I__10075\ : InMux
    port map (
            O => \N__43349\,
            I => \N__43330\
        );

    \I__10074\ : Span4Mux_h
    port map (
            O => \N__43346\,
            I => \N__43325\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__43343\,
            I => \N__43325\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43342\,
            I => \N__43322\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43319\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43316\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43313\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__43336\,
            I => \N__43309\
        );

    \I__10067\ : Span4Mux_h
    port map (
            O => \N__43333\,
            I => \N__43305\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43298\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__43325\,
            I => \N__43298\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__43322\,
            I => \N__43298\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43319\,
            I => \N__43293\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43316\,
            I => \N__43293\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43313\,
            I => \N__43290\
        );

    \I__10060\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43287\
        );

    \I__10059\ : Span4Mux_h
    port map (
            O => \N__43309\,
            I => \N__43283\
        );

    \I__10058\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43280\
        );

    \I__10057\ : Span4Mux_h
    port map (
            O => \N__43305\,
            I => \N__43277\
        );

    \I__10056\ : Span4Mux_v
    port map (
            O => \N__43298\,
            I => \N__43274\
        );

    \I__10055\ : Span4Mux_v
    port map (
            O => \N__43293\,
            I => \N__43267\
        );

    \I__10054\ : Span4Mux_h
    port map (
            O => \N__43290\,
            I => \N__43267\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__43287\,
            I => \N__43267\
        );

    \I__10052\ : InMux
    port map (
            O => \N__43286\,
            I => \N__43263\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__43283\,
            I => \N__43258\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43258\
        );

    \I__10049\ : Span4Mux_v
    port map (
            O => \N__43277\,
            I => \N__43253\
        );

    \I__10048\ : Span4Mux_h
    port map (
            O => \N__43274\,
            I => \N__43253\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__43267\,
            I => \N__43250\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43247\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__43263\,
            I => \N__43244\
        );

    \I__10044\ : Span4Mux_h
    port map (
            O => \N__43258\,
            I => \N__43239\
        );

    \I__10043\ : Span4Mux_v
    port map (
            O => \N__43253\,
            I => \N__43239\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__43250\,
            I => uart_pc_data_3
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__43247\,
            I => uart_pc_data_3
        );

    \I__10040\ : Odrv12
    port map (
            O => \N__43244\,
            I => uart_pc_data_3
        );

    \I__10039\ : Odrv4
    port map (
            O => \N__43239\,
            I => uart_pc_data_3
        );

    \I__10038\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43227\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__43227\,
            I => \N__43224\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__43224\,
            I => \N__43221\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__43221\,
            I => alt_ki_3
        );

    \I__10034\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43215\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43212\
        );

    \I__10032\ : Span4Mux_h
    port map (
            O => \N__43212\,
            I => \N__43209\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__43209\,
            I => \pid_alt.O_0_8\
        );

    \I__10030\ : CascadeMux
    port map (
            O => \N__43206\,
            I => \N__43203\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43203\,
            I => \N__43200\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__43200\,
            I => \N__43197\
        );

    \I__10027\ : Span12Mux_h
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__10026\ : Odrv12
    port map (
            O => \N__43194\,
            I => \pid_alt.error_i_regZ0Z_4\
        );

    \I__10025\ : InMux
    port map (
            O => \N__43191\,
            I => \N__43188\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__43188\,
            I => \N__43185\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__10022\ : Odrv4
    port map (
            O => \N__43182\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__10021\ : CascadeMux
    port map (
            O => \N__43179\,
            I => \N__43176\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43173\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__10018\ : Odrv4
    port map (
            O => \N__43170\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__10017\ : InMux
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43164\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__10015\ : InMux
    port map (
            O => \N__43161\,
            I => \N__43158\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43158\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__10013\ : CascadeMux
    port map (
            O => \N__43155\,
            I => \N__43152\
        );

    \I__10012\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43149\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__43149\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__10010\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43143\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43143\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__10008\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43135\
        );

    \I__10007\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43132\
        );

    \I__10006\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43119\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__43135\,
            I => \N__43111\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__43132\,
            I => \N__43111\
        );

    \I__10003\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43107\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43130\,
            I => \N__43104\
        );

    \I__10001\ : InMux
    port map (
            O => \N__43129\,
            I => \N__43101\
        );

    \I__10000\ : InMux
    port map (
            O => \N__43128\,
            I => \N__43098\
        );

    \I__9999\ : InMux
    port map (
            O => \N__43127\,
            I => \N__43093\
        );

    \I__9998\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43093\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43088\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43088\
        );

    \I__9995\ : CascadeMux
    port map (
            O => \N__43123\,
            I => \N__43082\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43122\,
            I => \N__43078\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43075\
        );

    \I__9992\ : CascadeMux
    port map (
            O => \N__43118\,
            I => \N__43071\
        );

    \I__9991\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43065\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43062\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__43111\,
            I => \N__43059\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43056\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__43107\,
            I => \N__43047\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__43104\,
            I => \N__43042\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__43101\,
            I => \N__43042\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43035\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__43093\,
            I => \N__43035\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__43088\,
            I => \N__43035\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43030\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43030\
        );

    \I__9979\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43027\
        );

    \I__9978\ : InMux
    port map (
            O => \N__43082\,
            I => \N__43024\
        );

    \I__9977\ : CascadeMux
    port map (
            O => \N__43081\,
            I => \N__43021\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__43078\,
            I => \N__43017\
        );

    \I__9975\ : Span4Mux_s2_h
    port map (
            O => \N__43075\,
            I => \N__43014\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43074\,
            I => \N__43009\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43071\,
            I => \N__43009\
        );

    \I__9972\ : CascadeMux
    port map (
            O => \N__43070\,
            I => \N__43004\
        );

    \I__9971\ : CascadeMux
    port map (
            O => \N__43069\,
            I => \N__43000\
        );

    \I__9970\ : CascadeMux
    port map (
            O => \N__43068\,
            I => \N__42996\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43065\,
            I => \N__42989\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__42989\
        );

    \I__9967\ : Span4Mux_h
    port map (
            O => \N__43059\,
            I => \N__42984\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__43056\,
            I => \N__42984\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43055\,
            I => \N__42979\
        );

    \I__9964\ : InMux
    port map (
            O => \N__43054\,
            I => \N__42979\
        );

    \I__9963\ : InMux
    port map (
            O => \N__43053\,
            I => \N__42976\
        );

    \I__9962\ : InMux
    port map (
            O => \N__43052\,
            I => \N__42971\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43051\,
            I => \N__42971\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__43050\,
            I => \N__42968\
        );

    \I__9959\ : Span4Mux_v
    port map (
            O => \N__43047\,
            I => \N__42963\
        );

    \I__9958\ : Span4Mux_v
    port map (
            O => \N__43042\,
            I => \N__42963\
        );

    \I__9957\ : Span4Mux_v
    port map (
            O => \N__43035\,
            I => \N__42956\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__43030\,
            I => \N__42956\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__43027\,
            I => \N__42956\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__43024\,
            I => \N__42953\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43021\,
            I => \N__42950\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__43020\,
            I => \N__42947\
        );

    \I__9951\ : Span4Mux_s3_h
    port map (
            O => \N__43017\,
            I => \N__42944\
        );

    \I__9950\ : Span4Mux_h
    port map (
            O => \N__43014\,
            I => \N__42939\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__43009\,
            I => \N__42939\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43008\,
            I => \N__42924\
        );

    \I__9947\ : InMux
    port map (
            O => \N__43007\,
            I => \N__42924\
        );

    \I__9946\ : InMux
    port map (
            O => \N__43004\,
            I => \N__42924\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42924\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42924\
        );

    \I__9943\ : InMux
    port map (
            O => \N__42999\,
            I => \N__42924\
        );

    \I__9942\ : InMux
    port map (
            O => \N__42996\,
            I => \N__42924\
        );

    \I__9941\ : CascadeMux
    port map (
            O => \N__42995\,
            I => \N__42920\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42917\
        );

    \I__9939\ : Span4Mux_v
    port map (
            O => \N__42989\,
            I => \N__42913\
        );

    \I__9938\ : Span4Mux_v
    port map (
            O => \N__42984\,
            I => \N__42908\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__42979\,
            I => \N__42908\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__42976\,
            I => \N__42903\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__42971\,
            I => \N__42903\
        );

    \I__9934\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42900\
        );

    \I__9933\ : Span4Mux_v
    port map (
            O => \N__42963\,
            I => \N__42895\
        );

    \I__9932\ : Span4Mux_v
    port map (
            O => \N__42956\,
            I => \N__42895\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__42953\,
            I => \N__42890\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__42950\,
            I => \N__42890\
        );

    \I__9929\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42887\
        );

    \I__9928\ : Span4Mux_v
    port map (
            O => \N__42944\,
            I => \N__42882\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__42939\,
            I => \N__42877\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__42924\,
            I => \N__42877\
        );

    \I__9925\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42870\
        );

    \I__9924\ : InMux
    port map (
            O => \N__42920\,
            I => \N__42870\
        );

    \I__9923\ : InMux
    port map (
            O => \N__42917\,
            I => \N__42870\
        );

    \I__9922\ : CascadeMux
    port map (
            O => \N__42916\,
            I => \N__42867\
        );

    \I__9921\ : Span4Mux_v
    port map (
            O => \N__42913\,
            I => \N__42862\
        );

    \I__9920\ : Span4Mux_v
    port map (
            O => \N__42908\,
            I => \N__42862\
        );

    \I__9919\ : Span4Mux_v
    port map (
            O => \N__42903\,
            I => \N__42859\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__42900\,
            I => \N__42856\
        );

    \I__9917\ : Span4Mux_h
    port map (
            O => \N__42895\,
            I => \N__42853\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__42890\,
            I => \N__42848\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__42887\,
            I => \N__42848\
        );

    \I__9914\ : InMux
    port map (
            O => \N__42886\,
            I => \N__42845\
        );

    \I__9913\ : CascadeMux
    port map (
            O => \N__42885\,
            I => \N__42842\
        );

    \I__9912\ : Span4Mux_h
    port map (
            O => \N__42882\,
            I => \N__42838\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__42877\,
            I => \N__42835\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__42870\,
            I => \N__42832\
        );

    \I__9909\ : InMux
    port map (
            O => \N__42867\,
            I => \N__42829\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__42862\,
            I => \N__42824\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__42859\,
            I => \N__42824\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__42856\,
            I => \N__42821\
        );

    \I__9905\ : Span4Mux_h
    port map (
            O => \N__42853\,
            I => \N__42816\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__42848\,
            I => \N__42816\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__42845\,
            I => \N__42813\
        );

    \I__9902\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42810\
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__42841\,
            I => \N__42807\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__42838\,
            I => \N__42802\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__42835\,
            I => \N__42802\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__42832\,
            I => \N__42797\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__42829\,
            I => \N__42797\
        );

    \I__9896\ : Span4Mux_h
    port map (
            O => \N__42824\,
            I => \N__42788\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__42821\,
            I => \N__42788\
        );

    \I__9894\ : Span4Mux_h
    port map (
            O => \N__42816\,
            I => \N__42788\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__42813\,
            I => \N__42788\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__42810\,
            I => \N__42785\
        );

    \I__9891\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42782\
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__42802\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9889\ : Odrv4
    port map (
            O => \N__42797\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9888\ : Odrv4
    port map (
            O => \N__42788\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9887\ : Odrv12
    port map (
            O => \N__42785\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__42782\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9885\ : CascadeMux
    port map (
            O => \N__42771\,
            I => \N__42768\
        );

    \I__9884\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42765\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__42765\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__9882\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42759\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42756\
        );

    \I__9880\ : Span12Mux_v
    port map (
            O => \N__42756\,
            I => \N__42753\
        );

    \I__9879\ : Odrv12
    port map (
            O => \N__42753\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__9878\ : InMux
    port map (
            O => \N__42750\,
            I => \N__42747\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__42747\,
            I => \N__42744\
        );

    \I__9876\ : Odrv12
    port map (
            O => \N__42744\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__42741\,
            I => \N__42737\
        );

    \I__9874\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42733\
        );

    \I__9873\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42730\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42736\,
            I => \N__42727\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42720\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42720\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__42727\,
            I => \N__42720\
        );

    \I__9868\ : Odrv4
    port map (
            O => \N__42720\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__9867\ : CascadeMux
    port map (
            O => \N__42717\,
            I => \N__42714\
        );

    \I__9866\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__42711\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__9864\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42703\
        );

    \I__9863\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42700\
        );

    \I__9862\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42697\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__42703\,
            I => \N__42692\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__42700\,
            I => \N__42692\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__42697\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__42692\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__9857\ : InMux
    port map (
            O => \N__42687\,
            I => \N__42684\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__42684\,
            I => \N__42681\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__42675\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__9852\ : InMux
    port map (
            O => \N__42672\,
            I => \N__42669\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__42663\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__9848\ : InMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__42657\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__9846\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__9844\ : Span4Mux_h
    port map (
            O => \N__42648\,
            I => \N__42645\
        );

    \I__9843\ : Odrv4
    port map (
            O => \N__42645\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__9842\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42639\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__42639\,
            I => \N__42636\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__42636\,
            I => \N__42633\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__42633\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__9838\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42627\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42624\
        );

    \I__9836\ : Span4Mux_h
    port map (
            O => \N__42624\,
            I => \N__42621\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__42621\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__42618\,
            I => \N__42613\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__42617\,
            I => \N__42600\
        );

    \I__9832\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42591\
        );

    \I__9831\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42591\
        );

    \I__9830\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42591\
        );

    \I__9829\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42580\
        );

    \I__9828\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42580\
        );

    \I__9827\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42580\
        );

    \I__9826\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42580\
        );

    \I__9825\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42580\
        );

    \I__9824\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42573\
        );

    \I__9823\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42573\
        );

    \I__9822\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42573\
        );

    \I__9821\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42564\
        );

    \I__9820\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42564\
        );

    \I__9819\ : InMux
    port map (
            O => \N__42599\,
            I => \N__42564\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42598\,
            I => \N__42564\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__42591\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9816\ : LocalMux
    port map (
            O => \N__42580\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__42573\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__42564\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__9813\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__42549\,
            I => \N__42546\
        );

    \I__9810\ : Span4Mux_h
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9809\ : Odrv4
    port map (
            O => \N__42543\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__9808\ : CEMux
    port map (
            O => \N__42540\,
            I => \N__42535\
        );

    \I__9807\ : CEMux
    port map (
            O => \N__42539\,
            I => \N__42532\
        );

    \I__9806\ : CEMux
    port map (
            O => \N__42538\,
            I => \N__42528\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__42535\,
            I => \N__42525\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__42532\,
            I => \N__42522\
        );

    \I__9803\ : CEMux
    port map (
            O => \N__42531\,
            I => \N__42519\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42516\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__42525\,
            I => \N__42513\
        );

    \I__9800\ : Span4Mux_v
    port map (
            O => \N__42522\,
            I => \N__42510\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__42519\,
            I => \N__42507\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__42516\,
            I => \N__42504\
        );

    \I__9797\ : Span4Mux_h
    port map (
            O => \N__42513\,
            I => \N__42501\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__42510\,
            I => \N__42496\
        );

    \I__9795\ : Span4Mux_h
    port map (
            O => \N__42507\,
            I => \N__42496\
        );

    \I__9794\ : Odrv4
    port map (
            O => \N__42504\,
            I => \ppm_encoder_1.N_1330_0\
        );

    \I__9793\ : Odrv4
    port map (
            O => \N__42501\,
            I => \ppm_encoder_1.N_1330_0\
        );

    \I__9792\ : Odrv4
    port map (
            O => \N__42496\,
            I => \ppm_encoder_1.N_1330_0\
        );

    \I__9791\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42486\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__42486\,
            I => \N__42481\
        );

    \I__9789\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42478\
        );

    \I__9788\ : InMux
    port map (
            O => \N__42484\,
            I => \N__42475\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__42481\,
            I => \N__42472\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__42478\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__42475\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__9784\ : Odrv4
    port map (
            O => \N__42472\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__42462\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__42459\,
            I => \N__42456\
        );

    \I__9780\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42453\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__9778\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42447\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__42447\,
            I => \N__42442\
        );

    \I__9776\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42439\
        );

    \I__9775\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42436\
        );

    \I__9774\ : Span4Mux_h
    port map (
            O => \N__42442\,
            I => \N__42433\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__42439\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__42436\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__9771\ : Odrv4
    port map (
            O => \N__42433\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__9770\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42423\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__42420\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__9767\ : CascadeMux
    port map (
            O => \N__42417\,
            I => \N__42414\
        );

    \I__9766\ : InMux
    port map (
            O => \N__42414\,
            I => \N__42411\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__42411\,
            I => \N__42408\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__42408\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__42402\,
            I => \N__42399\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__42399\,
            I => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\
        );

    \I__9760\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42393\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42390\
        );

    \I__9758\ : Odrv12
    port map (
            O => \N__42390\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__9757\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42384\,
            I => \N__42381\
        );

    \I__9755\ : Odrv12
    port map (
            O => \N__42381\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__9754\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42375\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__42375\,
            I => \N__42372\
        );

    \I__9752\ : Odrv4
    port map (
            O => \N__42372\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__9751\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42366\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__42366\,
            I => \N__42363\
        );

    \I__9749\ : Span4Mux_h
    port map (
            O => \N__42363\,
            I => \N__42358\
        );

    \I__9748\ : InMux
    port map (
            O => \N__42362\,
            I => \N__42353\
        );

    \I__9747\ : InMux
    port map (
            O => \N__42361\,
            I => \N__42353\
        );

    \I__9746\ : Odrv4
    port map (
            O => \N__42358\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__42353\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42348\,
            I => \N__42343\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42338\
        );

    \I__9742\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42338\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42343\,
            I => \N__42334\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__42338\,
            I => \N__42331\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42337\,
            I => \N__42328\
        );

    \I__9738\ : Span4Mux_v
    port map (
            O => \N__42334\,
            I => \N__42320\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__42331\,
            I => \N__42317\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42314\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42311\
        );

    \I__9734\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42302\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42302\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42302\
        );

    \I__9731\ : InMux
    port map (
            O => \N__42323\,
            I => \N__42302\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__42320\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__42317\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9728\ : Odrv12
    port map (
            O => \N__42314\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__42311\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42302\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__42291\,
            I => \N__42281\
        );

    \I__9724\ : CascadeMux
    port map (
            O => \N__42290\,
            I => \N__42278\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42267\
        );

    \I__9722\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42260\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42287\,
            I => \N__42260\
        );

    \I__9720\ : InMux
    port map (
            O => \N__42286\,
            I => \N__42260\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__42285\,
            I => \N__42255\
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__42284\,
            I => \N__42251\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42281\,
            I => \N__42238\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42238\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42238\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42238\
        );

    \I__9713\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42235\
        );

    \I__9712\ : InMux
    port map (
            O => \N__42274\,
            I => \N__42225\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42273\,
            I => \N__42222\
        );

    \I__9710\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42219\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42271\,
            I => \N__42214\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42214\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__42267\,
            I => \N__42209\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__42260\,
            I => \N__42209\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42204\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42204\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42195\
        );

    \I__9702\ : InMux
    port map (
            O => \N__42254\,
            I => \N__42195\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42195\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42195\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42188\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42188\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42188\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42238\,
            I => \N__42185\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42235\,
            I => \N__42182\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42179\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42176\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__42232\,
            I => \N__42173\
        );

    \I__9691\ : CascadeMux
    port map (
            O => \N__42231\,
            I => \N__42168\
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__42230\,
            I => \N__42159\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42155\
        );

    \I__9688\ : CascadeMux
    port map (
            O => \N__42228\,
            I => \N__42152\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__42225\,
            I => \N__42148\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__42222\,
            I => \N__42133\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__42219\,
            I => \N__42133\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__42214\,
            I => \N__42133\
        );

    \I__9683\ : Span4Mux_v
    port map (
            O => \N__42209\,
            I => \N__42133\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__42204\,
            I => \N__42133\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__42195\,
            I => \N__42133\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__42188\,
            I => \N__42133\
        );

    \I__9679\ : Span4Mux_v
    port map (
            O => \N__42185\,
            I => \N__42130\
        );

    \I__9678\ : Span4Mux_v
    port map (
            O => \N__42182\,
            I => \N__42127\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42122\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__42176\,
            I => \N__42122\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42115\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42115\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42115\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42111\
        );

    \I__9671\ : InMux
    port map (
            O => \N__42167\,
            I => \N__42106\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42166\,
            I => \N__42106\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42097\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42164\,
            I => \N__42097\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42163\,
            I => \N__42097\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42162\,
            I => \N__42097\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42092\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42158\,
            I => \N__42092\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__42155\,
            I => \N__42089\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42084\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42084\
        );

    \I__9660\ : Span4Mux_h
    port map (
            O => \N__42148\,
            I => \N__42077\
        );

    \I__9659\ : Span4Mux_v
    port map (
            O => \N__42133\,
            I => \N__42077\
        );

    \I__9658\ : Span4Mux_v
    port map (
            O => \N__42130\,
            I => \N__42077\
        );

    \I__9657\ : Span4Mux_h
    port map (
            O => \N__42127\,
            I => \N__42070\
        );

    \I__9656\ : Span4Mux_v
    port map (
            O => \N__42122\,
            I => \N__42070\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42115\,
            I => \N__42070\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42067\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__42111\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42106\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__42097\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__42092\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9649\ : Odrv4
    port map (
            O => \N__42089\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__42084\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__42077\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__42070\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42067\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__9644\ : CascadeMux
    port map (
            O => \N__42048\,
            I => \N__42044\
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__42047\,
            I => \N__42031\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42024\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42043\,
            I => \N__42024\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42042\,
            I => \N__42024\
        );

    \I__9639\ : CascadeMux
    port map (
            O => \N__42041\,
            I => \N__42015\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__42040\,
            I => \N__42012\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__42039\,
            I => \N__42004\
        );

    \I__9636\ : InMux
    port map (
            O => \N__42038\,
            I => \N__41999\
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__42037\,
            I => \N__41988\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__42036\,
            I => \N__41985\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42035\,
            I => \N__41979\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42034\,
            I => \N__41979\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42031\,
            I => \N__41972\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__42024\,
            I => \N__41969\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42023\,
            I => \N__41964\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42022\,
            I => \N__41964\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42021\,
            I => \N__41955\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42020\,
            I => \N__41955\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42019\,
            I => \N__41955\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42018\,
            I => \N__41955\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42015\,
            I => \N__41948\
        );

    \I__9622\ : InMux
    port map (
            O => \N__42012\,
            I => \N__41948\
        );

    \I__9621\ : InMux
    port map (
            O => \N__42011\,
            I => \N__41948\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42010\,
            I => \N__41933\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42009\,
            I => \N__41930\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42008\,
            I => \N__41925\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41925\
        );

    \I__9616\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41916\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41916\
        );

    \I__9614\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41913\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__41999\,
            I => \N__41910\
        );

    \I__9612\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41905\
        );

    \I__9611\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41905\
        );

    \I__9610\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41900\
        );

    \I__9609\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41900\
        );

    \I__9608\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41893\
        );

    \I__9607\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41893\
        );

    \I__9606\ : InMux
    port map (
            O => \N__41992\,
            I => \N__41893\
        );

    \I__9605\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41883\
        );

    \I__9604\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41883\
        );

    \I__9603\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41883\
        );

    \I__9602\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41883\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__41979\,
            I => \N__41880\
        );

    \I__9600\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41871\
        );

    \I__9599\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41871\
        );

    \I__9598\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41871\
        );

    \I__9597\ : InMux
    port map (
            O => \N__41975\,
            I => \N__41871\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__41972\,
            I => \N__41864\
        );

    \I__9595\ : Span4Mux_v
    port map (
            O => \N__41969\,
            I => \N__41864\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41864\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41859\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__41948\,
            I => \N__41859\
        );

    \I__9591\ : InMux
    port map (
            O => \N__41947\,
            I => \N__41848\
        );

    \I__9590\ : InMux
    port map (
            O => \N__41946\,
            I => \N__41848\
        );

    \I__9589\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41848\
        );

    \I__9588\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41848\
        );

    \I__9587\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41848\
        );

    \I__9586\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41841\
        );

    \I__9585\ : InMux
    port map (
            O => \N__41941\,
            I => \N__41841\
        );

    \I__9584\ : InMux
    port map (
            O => \N__41940\,
            I => \N__41841\
        );

    \I__9583\ : InMux
    port map (
            O => \N__41939\,
            I => \N__41837\
        );

    \I__9582\ : InMux
    port map (
            O => \N__41938\,
            I => \N__41830\
        );

    \I__9581\ : InMux
    port map (
            O => \N__41937\,
            I => \N__41830\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41830\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__41933\,
            I => \N__41827\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__41930\,
            I => \N__41822\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__41925\,
            I => \N__41822\
        );

    \I__9576\ : InMux
    port map (
            O => \N__41924\,
            I => \N__41817\
        );

    \I__9575\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41817\
        );

    \I__9574\ : InMux
    port map (
            O => \N__41922\,
            I => \N__41811\
        );

    \I__9573\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41808\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41795\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__41913\,
            I => \N__41795\
        );

    \I__9570\ : Span4Mux_v
    port map (
            O => \N__41910\,
            I => \N__41795\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__41905\,
            I => \N__41795\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__41900\,
            I => \N__41795\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__41893\,
            I => \N__41795\
        );

    \I__9566\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41792\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41785\
        );

    \I__9564\ : Span4Mux_v
    port map (
            O => \N__41880\,
            I => \N__41785\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__41871\,
            I => \N__41785\
        );

    \I__9562\ : Span4Mux_v
    port map (
            O => \N__41864\,
            I => \N__41778\
        );

    \I__9561\ : Span4Mux_v
    port map (
            O => \N__41859\,
            I => \N__41778\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__41848\,
            I => \N__41778\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__41841\,
            I => \N__41767\
        );

    \I__9558\ : InMux
    port map (
            O => \N__41840\,
            I => \N__41764\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__41837\,
            I => \N__41759\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__41830\,
            I => \N__41759\
        );

    \I__9555\ : Span4Mux_h
    port map (
            O => \N__41827\,
            I => \N__41752\
        );

    \I__9554\ : Span4Mux_v
    port map (
            O => \N__41822\,
            I => \N__41752\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41752\
        );

    \I__9552\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41747\
        );

    \I__9551\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41747\
        );

    \I__9550\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41744\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__41811\,
            I => \N__41741\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__41808\,
            I => \N__41736\
        );

    \I__9547\ : Span4Mux_v
    port map (
            O => \N__41795\,
            I => \N__41736\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__41792\,
            I => \N__41729\
        );

    \I__9545\ : Span4Mux_h
    port map (
            O => \N__41785\,
            I => \N__41729\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__41778\,
            I => \N__41729\
        );

    \I__9543\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41726\
        );

    \I__9542\ : InMux
    port map (
            O => \N__41776\,
            I => \N__41723\
        );

    \I__9541\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41710\
        );

    \I__9540\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41710\
        );

    \I__9539\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41710\
        );

    \I__9538\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41710\
        );

    \I__9537\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41710\
        );

    \I__9536\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41710\
        );

    \I__9535\ : Span4Mux_h
    port map (
            O => \N__41767\,
            I => \N__41701\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__41764\,
            I => \N__41701\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__41759\,
            I => \N__41701\
        );

    \I__9532\ : Span4Mux_v
    port map (
            O => \N__41752\,
            I => \N__41701\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__41747\,
            I => \N__41698\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41691\
        );

    \I__9529\ : Span4Mux_v
    port map (
            O => \N__41741\,
            I => \N__41691\
        );

    \I__9528\ : Span4Mux_v
    port map (
            O => \N__41736\,
            I => \N__41691\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__41729\,
            I => \N__41688\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__41726\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__41723\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__41710\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9523\ : Odrv4
    port map (
            O => \N__41701\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9522\ : Odrv12
    port map (
            O => \N__41698\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9521\ : Odrv4
    port map (
            O => \N__41691\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__41688\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__9519\ : InMux
    port map (
            O => \N__41673\,
            I => \N__41670\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__41670\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__9517\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41664\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41661\
        );

    \I__9515\ : Odrv12
    port map (
            O => \N__41661\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__9514\ : InMux
    port map (
            O => \N__41658\,
            I => \N__41655\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__41655\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__9512\ : CascadeMux
    port map (
            O => \N__41652\,
            I => \N__41648\
        );

    \I__9511\ : InMux
    port map (
            O => \N__41651\,
            I => \N__41645\
        );

    \I__9510\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41642\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__41645\,
            I => \N__41638\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__41642\,
            I => \N__41635\
        );

    \I__9507\ : CascadeMux
    port map (
            O => \N__41641\,
            I => \N__41632\
        );

    \I__9506\ : Span4Mux_v
    port map (
            O => \N__41638\,
            I => \N__41627\
        );

    \I__9505\ : Span4Mux_h
    port map (
            O => \N__41635\,
            I => \N__41627\
        );

    \I__9504\ : InMux
    port map (
            O => \N__41632\,
            I => \N__41624\
        );

    \I__9503\ : Odrv4
    port map (
            O => \N__41627\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__41624\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__9501\ : CascadeMux
    port map (
            O => \N__41619\,
            I => \N__41603\
        );

    \I__9500\ : CascadeMux
    port map (
            O => \N__41618\,
            I => \N__41596\
        );

    \I__9499\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41590\
        );

    \I__9498\ : InMux
    port map (
            O => \N__41616\,
            I => \N__41590\
        );

    \I__9497\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41587\
        );

    \I__9496\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41584\
        );

    \I__9495\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41579\
        );

    \I__9494\ : InMux
    port map (
            O => \N__41612\,
            I => \N__41579\
        );

    \I__9493\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41576\
        );

    \I__9492\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41573\
        );

    \I__9491\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41566\
        );

    \I__9490\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41566\
        );

    \I__9489\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41566\
        );

    \I__9488\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41557\
        );

    \I__9487\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41557\
        );

    \I__9486\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41557\
        );

    \I__9485\ : InMux
    port map (
            O => \N__41601\,
            I => \N__41557\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41552\
        );

    \I__9483\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41552\
        );

    \I__9482\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41547\
        );

    \I__9481\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41547\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__41590\,
            I => \N__41542\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__41587\,
            I => \N__41542\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__41584\,
            I => \N__41537\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41537\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__41576\,
            I => \N__41534\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41529\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__41566\,
            I => \N__41529\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__41557\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__41552\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__41547\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9470\ : Odrv4
    port map (
            O => \N__41542\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9469\ : Odrv4
    port map (
            O => \N__41537\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9468\ : Odrv4
    port map (
            O => \N__41534\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9467\ : Odrv12
    port map (
            O => \N__41529\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9466\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41511\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__9464\ : Span4Mux_v
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__41505\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__9462\ : CascadeMux
    port map (
            O => \N__41502\,
            I => \N__41493\
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__41501\,
            I => \N__41490\
        );

    \I__9460\ : CascadeMux
    port map (
            O => \N__41500\,
            I => \N__41487\
        );

    \I__9459\ : CascadeMux
    port map (
            O => \N__41499\,
            I => \N__41484\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__41498\,
            I => \N__41481\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__41497\,
            I => \N__41478\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__41496\,
            I => \N__41475\
        );

    \I__9455\ : InMux
    port map (
            O => \N__41493\,
            I => \N__41466\
        );

    \I__9454\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41466\
        );

    \I__9453\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41466\
        );

    \I__9452\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41463\
        );

    \I__9451\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41458\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41478\,
            I => \N__41458\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41455\
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__41474\,
            I => \N__41452\
        );

    \I__9447\ : CascadeMux
    port map (
            O => \N__41473\,
            I => \N__41449\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__41466\,
            I => \N__41435\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__41463\,
            I => \N__41435\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41458\,
            I => \N__41435\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__41455\,
            I => \N__41435\
        );

    \I__9442\ : InMux
    port map (
            O => \N__41452\,
            I => \N__41430\
        );

    \I__9441\ : InMux
    port map (
            O => \N__41449\,
            I => \N__41430\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__41448\,
            I => \N__41427\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__41447\,
            I => \N__41424\
        );

    \I__9438\ : CascadeMux
    port map (
            O => \N__41446\,
            I => \N__41420\
        );

    \I__9437\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41416\
        );

    \I__9436\ : CascadeMux
    port map (
            O => \N__41444\,
            I => \N__41413\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__41435\,
            I => \N__41406\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__41430\,
            I => \N__41406\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41427\,
            I => \N__41403\
        );

    \I__9432\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41400\
        );

    \I__9431\ : InMux
    port map (
            O => \N__41423\,
            I => \N__41393\
        );

    \I__9430\ : InMux
    port map (
            O => \N__41420\,
            I => \N__41393\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41419\,
            I => \N__41393\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__41416\,
            I => \N__41390\
        );

    \I__9427\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41387\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__41412\,
            I => \N__41384\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__41411\,
            I => \N__41381\
        );

    \I__9424\ : Span4Mux_v
    port map (
            O => \N__41406\,
            I => \N__41377\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__41403\,
            I => \N__41370\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__41400\,
            I => \N__41370\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__41393\,
            I => \N__41370\
        );

    \I__9420\ : Span4Mux_h
    port map (
            O => \N__41390\,
            I => \N__41365\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__41387\,
            I => \N__41365\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41360\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41381\,
            I => \N__41360\
        );

    \I__9416\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41357\
        );

    \I__9415\ : Odrv4
    port map (
            O => \N__41377\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__41370\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__41365\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__41360\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41357\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9410\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41343\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__9408\ : Odrv4
    port map (
            O => \N__41340\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__9407\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41333\
        );

    \I__9406\ : CascadeMux
    port map (
            O => \N__41336\,
            I => \N__41329\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41326\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41323\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41329\,
            I => \N__41320\
        );

    \I__9402\ : Span4Mux_v
    port map (
            O => \N__41326\,
            I => \N__41317\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41314\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__41320\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__41317\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__41314\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41307\,
            I => \N__41304\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__41304\,
            I => \N__41301\
        );

    \I__9395\ : Odrv4
    port map (
            O => \N__41301\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41298\,
            I => \N__41295\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__41295\,
            I => \N__41292\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__41292\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__9391\ : InMux
    port map (
            O => \N__41289\,
            I => \N__41286\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__41286\,
            I => \N__41283\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__41283\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__9388\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41277\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__41277\,
            I => \N__41274\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__41274\,
            I => \N__41271\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__41271\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41268\,
            I => \N__41265\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41265\,
            I => \N__41262\
        );

    \I__9382\ : Span4Mux_h
    port map (
            O => \N__41262\,
            I => \N__41259\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__41259\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__9380\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41253\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41250\
        );

    \I__9378\ : Odrv4
    port map (
            O => \N__41250\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41243\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41246\,
            I => \N__41239\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__41243\,
            I => \N__41236\
        );

    \I__9374\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41233\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41239\,
            I => \N__41230\
        );

    \I__9372\ : Span4Mux_v
    port map (
            O => \N__41236\,
            I => \N__41227\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__41233\,
            I => \N__41222\
        );

    \I__9370\ : Span4Mux_v
    port map (
            O => \N__41230\,
            I => \N__41222\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__41227\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__41222\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41217\,
            I => \N__41214\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__41214\,
            I => \N__41211\
        );

    \I__9365\ : Span4Mux_v
    port map (
            O => \N__41211\,
            I => \N__41208\
        );

    \I__9364\ : Odrv4
    port map (
            O => \N__41208\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41205\,
            I => \N__41202\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41202\,
            I => \N__41199\
        );

    \I__9361\ : Odrv12
    port map (
            O => \N__41199\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__9360\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41193\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41193\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__9358\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41187\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41184\
        );

    \I__9356\ : Span4Mux_v
    port map (
            O => \N__41184\,
            I => \N__41180\
        );

    \I__9355\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41177\
        );

    \I__9354\ : Odrv4
    port map (
            O => \N__41180\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41177\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__9352\ : InMux
    port map (
            O => \N__41172\,
            I => \N__41169\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__9350\ : Span4Mux_v
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__9349\ : Odrv4
    port map (
            O => \N__41163\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__9348\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41151\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41151\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41158\,
            I => \N__41151\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__41151\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41148\,
            I => \N__41142\
        );

    \I__9343\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41138\
        );

    \I__9342\ : InMux
    port map (
            O => \N__41146\,
            I => \N__41133\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41133\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__41142\,
            I => \N__41129\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41125\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__41138\,
            I => \N__41118\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__41133\,
            I => \N__41115\
        );

    \I__9336\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41112\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__41129\,
            I => \N__41109\
        );

    \I__9334\ : InMux
    port map (
            O => \N__41128\,
            I => \N__41106\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__41125\,
            I => \N__41103\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41098\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41098\
        );

    \I__9330\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41095\
        );

    \I__9329\ : CascadeMux
    port map (
            O => \N__41121\,
            I => \N__41091\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__41118\,
            I => \N__41084\
        );

    \I__9327\ : Span4Mux_h
    port map (
            O => \N__41115\,
            I => \N__41084\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__41112\,
            I => \N__41084\
        );

    \I__9325\ : Span4Mux_h
    port map (
            O => \N__41109\,
            I => \N__41079\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41079\
        );

    \I__9323\ : Span4Mux_v
    port map (
            O => \N__41103\,
            I => \N__41074\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__41098\,
            I => \N__41074\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41095\,
            I => \N__41071\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41094\,
            I => \N__41068\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41065\
        );

    \I__9318\ : Span4Mux_v
    port map (
            O => \N__41084\,
            I => \N__41059\
        );

    \I__9317\ : Span4Mux_v
    port map (
            O => \N__41079\,
            I => \N__41054\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__41074\,
            I => \N__41054\
        );

    \I__9315\ : Span4Mux_h
    port map (
            O => \N__41071\,
            I => \N__41051\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41068\,
            I => \N__41046\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__41065\,
            I => \N__41046\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41041\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41041\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41062\,
            I => \N__41038\
        );

    \I__9309\ : Odrv4
    port map (
            O => \N__41059\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9308\ : Odrv4
    port map (
            O => \N__41054\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__41051\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9306\ : Odrv12
    port map (
            O => \N__41046\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__41041\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__41038\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41022\,
            I => \N__41018\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41015\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__41012\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41009\
        );

    \I__9298\ : Span4Mux_h
    port map (
            O => \N__41012\,
            I => \N__41006\
        );

    \I__9297\ : Span4Mux_v
    port map (
            O => \N__41009\,
            I => \N__41003\
        );

    \I__9296\ : Span4Mux_h
    port map (
            O => \N__41006\,
            I => \N__41000\
        );

    \I__9295\ : Span4Mux_v
    port map (
            O => \N__41003\,
            I => \N__40997\
        );

    \I__9294\ : Odrv4
    port map (
            O => \N__41000\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__9293\ : Odrv4
    port map (
            O => \N__40997\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__40992\,
            I => \N__40985\
        );

    \I__9291\ : CascadeMux
    port map (
            O => \N__40991\,
            I => \N__40979\
        );

    \I__9290\ : InMux
    port map (
            O => \N__40990\,
            I => \N__40974\
        );

    \I__9289\ : InMux
    port map (
            O => \N__40989\,
            I => \N__40971\
        );

    \I__9288\ : InMux
    port map (
            O => \N__40988\,
            I => \N__40968\
        );

    \I__9287\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40965\
        );

    \I__9286\ : CascadeMux
    port map (
            O => \N__40984\,
            I => \N__40962\
        );

    \I__9285\ : CascadeMux
    port map (
            O => \N__40983\,
            I => \N__40959\
        );

    \I__9284\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40955\
        );

    \I__9283\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40952\
        );

    \I__9282\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40949\
        );

    \I__9281\ : CascadeMux
    port map (
            O => \N__40977\,
            I => \N__40945\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40936\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__40971\,
            I => \N__40936\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__40968\,
            I => \N__40936\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__40965\,
            I => \N__40936\
        );

    \I__9276\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40931\
        );

    \I__9275\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40931\
        );

    \I__9274\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40923\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40918\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__40952\,
            I => \N__40918\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__40949\,
            I => \N__40915\
        );

    \I__9270\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40910\
        );

    \I__9269\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40910\
        );

    \I__9268\ : Span4Mux_v
    port map (
            O => \N__40936\,
            I => \N__40904\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__40931\,
            I => \N__40904\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__40930\,
            I => \N__40901\
        );

    \I__9265\ : CascadeMux
    port map (
            O => \N__40929\,
            I => \N__40898\
        );

    \I__9264\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40895\
        );

    \I__9263\ : InMux
    port map (
            O => \N__40927\,
            I => \N__40892\
        );

    \I__9262\ : CascadeMux
    port map (
            O => \N__40926\,
            I => \N__40889\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__40923\,
            I => \N__40879\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__40918\,
            I => \N__40879\
        );

    \I__9259\ : Span4Mux_h
    port map (
            O => \N__40915\,
            I => \N__40879\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40910\,
            I => \N__40879\
        );

    \I__9257\ : InMux
    port map (
            O => \N__40909\,
            I => \N__40876\
        );

    \I__9256\ : Span4Mux_v
    port map (
            O => \N__40904\,
            I => \N__40873\
        );

    \I__9255\ : InMux
    port map (
            O => \N__40901\,
            I => \N__40870\
        );

    \I__9254\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40867\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__40895\,
            I => \N__40864\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__40892\,
            I => \N__40861\
        );

    \I__9251\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40858\
        );

    \I__9250\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40855\
        );

    \I__9249\ : Span4Mux_v
    port map (
            O => \N__40879\,
            I => \N__40852\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__40876\,
            I => \N__40849\
        );

    \I__9247\ : Sp12to4
    port map (
            O => \N__40873\,
            I => \N__40840\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__40870\,
            I => \N__40840\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__40867\,
            I => \N__40840\
        );

    \I__9244\ : Span12Mux_v
    port map (
            O => \N__40864\,
            I => \N__40840\
        );

    \I__9243\ : Span12Mux_v
    port map (
            O => \N__40861\,
            I => \N__40837\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__40858\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__40855\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9240\ : Odrv4
    port map (
            O => \N__40852\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__40849\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9238\ : Odrv12
    port map (
            O => \N__40840\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9237\ : Odrv12
    port map (
            O => \N__40837\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9236\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40821\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40818\
        );

    \I__9234\ : Odrv12
    port map (
            O => \N__40818\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__9233\ : InMux
    port map (
            O => \N__40815\,
            I => \N__40812\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__40812\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__9231\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40806\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__40806\,
            I => \N__40803\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__40803\,
            I => \N__40800\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__40800\,
            I => \N__40795\
        );

    \I__9227\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40792\
        );

    \I__9226\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40789\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__40795\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__40792\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__40789\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__9222\ : CascadeMux
    port map (
            O => \N__40782\,
            I => \N__40779\
        );

    \I__9221\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40776\,
            I => \N__40773\
        );

    \I__9219\ : Odrv12
    port map (
            O => \N__40773\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__9218\ : InMux
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__40767\,
            I => \N__40764\
        );

    \I__9216\ : Odrv12
    port map (
            O => \N__40764\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__9215\ : InMux
    port map (
            O => \N__40761\,
            I => \N__40758\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__40758\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__9213\ : InMux
    port map (
            O => \N__40755\,
            I => \N__40751\
        );

    \I__9212\ : InMux
    port map (
            O => \N__40754\,
            I => \N__40748\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__40751\,
            I => \N__40745\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__40748\,
            I => \N__40742\
        );

    \I__9209\ : Span4Mux_h
    port map (
            O => \N__40745\,
            I => \N__40738\
        );

    \I__9208\ : Span4Mux_v
    port map (
            O => \N__40742\,
            I => \N__40735\
        );

    \I__9207\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40732\
        );

    \I__9206\ : Span4Mux_h
    port map (
            O => \N__40738\,
            I => \N__40729\
        );

    \I__9205\ : Odrv4
    port map (
            O => \N__40735\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40732\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__40729\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__9202\ : CascadeMux
    port map (
            O => \N__40722\,
            I => \N__40719\
        );

    \I__9201\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40716\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__40713\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__9198\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40701\
        );

    \I__9197\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40701\
        );

    \I__9196\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40701\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__40701\,
            I => \N__40698\
        );

    \I__9194\ : Odrv4
    port map (
            O => \N__40698\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__9193\ : InMux
    port map (
            O => \N__40695\,
            I => \N__40692\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__40692\,
            I => \N__40687\
        );

    \I__9191\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40684\
        );

    \I__9190\ : CascadeMux
    port map (
            O => \N__40690\,
            I => \N__40681\
        );

    \I__9189\ : Span4Mux_v
    port map (
            O => \N__40687\,
            I => \N__40678\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__40684\,
            I => \N__40675\
        );

    \I__9187\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40672\
        );

    \I__9186\ : Span4Mux_h
    port map (
            O => \N__40678\,
            I => \N__40669\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__40675\,
            I => \N__40666\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__40672\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__40669\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__40666\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__9181\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40656\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__40656\,
            I => \N__40653\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__40653\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__9178\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40647\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__40647\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__9176\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40641\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__40641\,
            I => \N__40636\
        );

    \I__9174\ : InMux
    port map (
            O => \N__40640\,
            I => \N__40633\
        );

    \I__9173\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40630\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__40636\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__40633\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__40630\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9169\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40619\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__40622\,
            I => \N__40616\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N__40613\
        );

    \I__9166\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40610\
        );

    \I__9165\ : Span4Mux_v
    port map (
            O => \N__40613\,
            I => \N__40607\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__40610\,
            I => \N__40604\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__40607\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__40604\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__9161\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__40596\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__9159\ : InMux
    port map (
            O => \N__40593\,
            I => \N__40590\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__40590\,
            I => \N__40587\
        );

    \I__9157\ : Odrv12
    port map (
            O => \N__40587\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__9156\ : InMux
    port map (
            O => \N__40584\,
            I => \N__40581\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__9154\ : Odrv4
    port map (
            O => \N__40578\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__9153\ : CascadeMux
    port map (
            O => \N__40575\,
            I => \N__40571\
        );

    \I__9152\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40568\
        );

    \I__9151\ : InMux
    port map (
            O => \N__40571\,
            I => \N__40565\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__40568\,
            I => \N__40562\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__40565\,
            I => \N__40559\
        );

    \I__9148\ : Odrv12
    port map (
            O => \N__40562\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__40559\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__9146\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40545\
        );

    \I__9145\ : InMux
    port map (
            O => \N__40553\,
            I => \N__40545\
        );

    \I__9144\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40545\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__40545\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__40542\,
            I => \N__40539\
        );

    \I__9141\ : InMux
    port map (
            O => \N__40539\,
            I => \N__40536\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__40536\,
            I => \N__40532\
        );

    \I__9139\ : InMux
    port map (
            O => \N__40535\,
            I => \N__40528\
        );

    \I__9138\ : Span12Mux_h
    port map (
            O => \N__40532\,
            I => \N__40525\
        );

    \I__9137\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40522\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__40528\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__9135\ : Odrv12
    port map (
            O => \N__40525\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__40522\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__9133\ : InMux
    port map (
            O => \N__40515\,
            I => \N__40512\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40509\
        );

    \I__9131\ : Span4Mux_v
    port map (
            O => \N__40509\,
            I => \N__40506\
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__40506\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40503\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__9128\ : InMux
    port map (
            O => \N__40500\,
            I => \bfn_18_13_0_\
        );

    \I__9127\ : InMux
    port map (
            O => \N__40497\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__9126\ : InMux
    port map (
            O => \N__40494\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__9125\ : InMux
    port map (
            O => \N__40491\,
            I => \N__40486\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40482\
        );

    \I__9123\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40479\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__40486\,
            I => \N__40476\
        );

    \I__9121\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40473\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__40482\,
            I => \N__40468\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__40479\,
            I => \N__40465\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__40476\,
            I => \N__40460\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__40473\,
            I => \N__40460\
        );

    \I__9116\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40455\
        );

    \I__9115\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40455\
        );

    \I__9114\ : Span4Mux_h
    port map (
            O => \N__40468\,
            I => \N__40451\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__40465\,
            I => \N__40448\
        );

    \I__9112\ : Span4Mux_h
    port map (
            O => \N__40460\,
            I => \N__40443\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__40455\,
            I => \N__40443\
        );

    \I__9110\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40440\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__40451\,
            I => \N__40437\
        );

    \I__9108\ : Span4Mux_h
    port map (
            O => \N__40448\,
            I => \N__40432\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__40443\,
            I => \N__40432\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__40440\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9105\ : Odrv4
    port map (
            O => \N__40437\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__40432\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9103\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40422\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__40422\,
            I => \N__40418\
        );

    \I__9101\ : InMux
    port map (
            O => \N__40421\,
            I => \N__40415\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__40418\,
            I => \N__40412\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__40415\,
            I => \N__40409\
        );

    \I__9098\ : Span4Mux_v
    port map (
            O => \N__40412\,
            I => \N__40403\
        );

    \I__9097\ : Span4Mux_h
    port map (
            O => \N__40409\,
            I => \N__40400\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40397\
        );

    \I__9095\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40392\
        );

    \I__9094\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40392\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__40403\,
            I => \ppm_encoder_1.N_227\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__40400\,
            I => \ppm_encoder_1.N_227\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__40397\,
            I => \ppm_encoder_1.N_227\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__40392\,
            I => \ppm_encoder_1.N_227\
        );

    \I__9089\ : CascadeMux
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__9088\ : InMux
    port map (
            O => \N__40380\,
            I => \N__40374\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__40379\,
            I => \N__40370\
        );

    \I__9086\ : CascadeMux
    port map (
            O => \N__40378\,
            I => \N__40367\
        );

    \I__9085\ : CascadeMux
    port map (
            O => \N__40377\,
            I => \N__40364\
        );

    \I__9084\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40359\
        );

    \I__9083\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40352\
        );

    \I__9082\ : InMux
    port map (
            O => \N__40370\,
            I => \N__40352\
        );

    \I__9081\ : InMux
    port map (
            O => \N__40367\,
            I => \N__40352\
        );

    \I__9080\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40349\
        );

    \I__9079\ : InMux
    port map (
            O => \N__40363\,
            I => \N__40346\
        );

    \I__9078\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40343\
        );

    \I__9077\ : Span4Mux_h
    port map (
            O => \N__40359\,
            I => \N__40340\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__40352\,
            I => \N__40337\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__40349\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__40346\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__40343\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__40340\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__40337\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9070\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40322\
        );

    \I__9069\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40318\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__40322\,
            I => \N__40315\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__40321\,
            I => \N__40312\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40318\,
            I => \N__40309\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__40315\,
            I => \N__40306\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40312\,
            I => \N__40303\
        );

    \I__9063\ : Span4Mux_h
    port map (
            O => \N__40309\,
            I => \N__40296\
        );

    \I__9062\ : Span4Mux_v
    port map (
            O => \N__40306\,
            I => \N__40291\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__40303\,
            I => \N__40291\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40282\
        );

    \I__9059\ : InMux
    port map (
            O => \N__40301\,
            I => \N__40282\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40282\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40282\
        );

    \I__9056\ : Odrv4
    port map (
            O => \N__40296\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9055\ : Odrv4
    port map (
            O => \N__40291\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__40282\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9053\ : CascadeMux
    port map (
            O => \N__40275\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__40269\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40263\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__40263\,
            I => \N__40260\
        );

    \I__9048\ : Odrv4
    port map (
            O => \N__40260\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40254\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40248\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40248\,
            I => \N__40244\
        );

    \I__9043\ : CascadeMux
    port map (
            O => \N__40247\,
            I => \N__40241\
        );

    \I__9042\ : Span4Mux_h
    port map (
            O => \N__40244\,
            I => \N__40238\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40235\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__40238\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__40235\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__9038\ : InMux
    port map (
            O => \N__40230\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__9037\ : InMux
    port map (
            O => \N__40227\,
            I => \bfn_18_12_0_\
        );

    \I__9036\ : InMux
    port map (
            O => \N__40224\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__9035\ : InMux
    port map (
            O => \N__40221\,
            I => \N__40218\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__40218\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__9033\ : InMux
    port map (
            O => \N__40215\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__40209\,
            I => \N__40206\
        );

    \I__9030\ : Span4Mux_h
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__9028\ : Span4Mux_v
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__40197\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40191\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__40191\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40188\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40182\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__40182\,
            I => \N__40179\
        );

    \I__9021\ : Span12Mux_s11_h
    port map (
            O => \N__40179\,
            I => \N__40176\
        );

    \I__9020\ : Odrv12
    port map (
            O => \N__40176\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__9019\ : InMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__40170\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40167\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40161\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40161\,
            I => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\
        );

    \I__9014\ : CascadeMux
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__9013\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40152\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__40152\,
            I => \N__40149\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__40149\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40146\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40143\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__9008\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40137\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__40137\,
            I => \N__40122\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40136\,
            I => \N__40118\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40135\,
            I => \N__40115\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40134\,
            I => \N__40110\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40105\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40132\,
            I => \N__40105\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40102\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40130\,
            I => \N__40099\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40129\,
            I => \N__40096\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40128\,
            I => \N__40093\
        );

    \I__8997\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40088\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40126\,
            I => \N__40083\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40083\
        );

    \I__8994\ : Span4Mux_v
    port map (
            O => \N__40122\,
            I => \N__40080\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40077\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__40118\,
            I => \N__40072\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__40115\,
            I => \N__40072\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40069\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40066\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__40110\,
            I => \N__40059\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40105\,
            I => \N__40059\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40102\,
            I => \N__40059\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__40099\,
            I => \N__40056\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__40096\,
            I => \N__40052\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__40093\,
            I => \N__40049\
        );

    \I__8982\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40044\
        );

    \I__8981\ : InMux
    port map (
            O => \N__40091\,
            I => \N__40044\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__40088\,
            I => \N__40041\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__40083\,
            I => \N__40036\
        );

    \I__8978\ : Span4Mux_v
    port map (
            O => \N__40080\,
            I => \N__40036\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__40077\,
            I => \N__40033\
        );

    \I__8976\ : Span4Mux_h
    port map (
            O => \N__40072\,
            I => \N__40022\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40022\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__40022\
        );

    \I__8973\ : Span4Mux_v
    port map (
            O => \N__40059\,
            I => \N__40022\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__40056\,
            I => \N__40022\
        );

    \I__8971\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40019\
        );

    \I__8970\ : Span4Mux_v
    port map (
            O => \N__40052\,
            I => \N__40014\
        );

    \I__8969\ : Span4Mux_v
    port map (
            O => \N__40049\,
            I => \N__40014\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__40044\,
            I => \N__40007\
        );

    \I__8967\ : Span4Mux_v
    port map (
            O => \N__40041\,
            I => \N__40007\
        );

    \I__8966\ : Span4Mux_h
    port map (
            O => \N__40036\,
            I => \N__40007\
        );

    \I__8965\ : Span4Mux_v
    port map (
            O => \N__40033\,
            I => \N__40002\
        );

    \I__8964\ : Span4Mux_v
    port map (
            O => \N__40022\,
            I => \N__40002\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__40019\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__40014\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__40007\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__40002\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__8959\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39988\
        );

    \I__8958\ : InMux
    port map (
            O => \N__39992\,
            I => \N__39985\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__39991\,
            I => \N__39982\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__39988\,
            I => \N__39976\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__39985\,
            I => \N__39976\
        );

    \I__8954\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39971\
        );

    \I__8953\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39968\
        );

    \I__8952\ : Span4Mux_h
    port map (
            O => \N__39976\,
            I => \N__39965\
        );

    \I__8951\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39960\
        );

    \I__8950\ : InMux
    port map (
            O => \N__39974\,
            I => \N__39960\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__39971\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__39968\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__39965\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__39960\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__8945\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__39948\,
            I => \N__39945\
        );

    \I__8943\ : Odrv12
    port map (
            O => \N__39945\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\
        );

    \I__8942\ : CascadeMux
    port map (
            O => \N__39942\,
            I => \N__39939\
        );

    \I__8941\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39936\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__39936\,
            I => \N__39933\
        );

    \I__8939\ : Odrv4
    port map (
            O => \N__39933\,
            I => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\
        );

    \I__8938\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39927\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__39927\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__8936\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__39921\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__8934\ : InMux
    port map (
            O => \N__39918\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__8933\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39909\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__39909\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__8929\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__39900\,
            I => \N__39897\
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__39897\,
            I => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\
        );

    \I__8926\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__8924\ : Span4Mux_v
    port map (
            O => \N__39888\,
            I => \N__39885\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__39885\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__8922\ : InMux
    port map (
            O => \N__39882\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__8921\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8919\ : Span4Mux_h
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__8918\ : Odrv4
    port map (
            O => \N__39870\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__8917\ : InMux
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__39864\,
            I => \N__39861\
        );

    \I__8915\ : Span4Mux_v
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__8914\ : Odrv4
    port map (
            O => \N__39858\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__8913\ : InMux
    port map (
            O => \N__39855\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__8912\ : InMux
    port map (
            O => \N__39852\,
            I => \N__39849\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__39849\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__8910\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39843\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__39843\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__8908\ : InMux
    port map (
            O => \N__39840\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__8907\ : InMux
    port map (
            O => \N__39837\,
            I => \N__39834\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39834\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__8905\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39828\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__39828\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__8903\ : InMux
    port map (
            O => \N__39825\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__8902\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39819\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__39819\,
            I => \N__39816\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__39816\,
            I => \N__39813\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__39810\,
            I => \N__39807\
        );

    \I__8897\ : Odrv4
    port map (
            O => \N__39807\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\
        );

    \I__8896\ : CascadeMux
    port map (
            O => \N__39804\,
            I => \N__39801\
        );

    \I__8895\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39798\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__39798\,
            I => \N__39795\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__39795\,
            I => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\
        );

    \I__8892\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39789\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__39789\,
            I => \N__39786\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__39786\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__8889\ : InMux
    port map (
            O => \N__39783\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__8888\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39777\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__39777\,
            I => \N__39774\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__39774\,
            I => \N__39770\
        );

    \I__8885\ : InMux
    port map (
            O => \N__39773\,
            I => \N__39767\
        );

    \I__8884\ : Span4Mux_h
    port map (
            O => \N__39770\,
            I => \N__39764\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__39767\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__8882\ : Odrv4
    port map (
            O => \N__39764\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__8881\ : CascadeMux
    port map (
            O => \N__39759\,
            I => \N__39756\
        );

    \I__8880\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39750\
        );

    \I__8879\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39750\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__39750\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__39747\,
            I => \N__39743\
        );

    \I__8876\ : CascadeMux
    port map (
            O => \N__39746\,
            I => \N__39739\
        );

    \I__8875\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39731\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39731\
        );

    \I__8873\ : InMux
    port map (
            O => \N__39739\,
            I => \N__39731\
        );

    \I__8872\ : CascadeMux
    port map (
            O => \N__39738\,
            I => \N__39728\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__39731\,
            I => \N__39725\
        );

    \I__8870\ : InMux
    port map (
            O => \N__39728\,
            I => \N__39722\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__39725\,
            I => \N__39719\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__39722\,
            I => \N__39716\
        );

    \I__8867\ : Span4Mux_v
    port map (
            O => \N__39719\,
            I => \N__39713\
        );

    \I__8866\ : Span4Mux_h
    port map (
            O => \N__39716\,
            I => \N__39710\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__39713\,
            I => \N__39707\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__39710\,
            I => \N__39704\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__39707\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__39704\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\
        );

    \I__8861\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39694\
        );

    \I__8860\ : InMux
    port map (
            O => \N__39698\,
            I => \N__39689\
        );

    \I__8859\ : InMux
    port map (
            O => \N__39697\,
            I => \N__39689\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__39694\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__39689\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__8856\ : InMux
    port map (
            O => \N__39684\,
            I => \N__39679\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \N__39676\
        );

    \I__8854\ : InMux
    port map (
            O => \N__39682\,
            I => \N__39673\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39670\
        );

    \I__8852\ : InMux
    port map (
            O => \N__39676\,
            I => \N__39667\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__39673\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__39670\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__39667\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__8848\ : CascadeMux
    port map (
            O => \N__39660\,
            I => \N__39656\
        );

    \I__8847\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39652\
        );

    \I__8846\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39647\
        );

    \I__8845\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39647\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__39652\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__39647\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__8842\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39638\
        );

    \I__8841\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39635\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__39638\,
            I => \N__39630\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__39635\,
            I => \N__39630\
        );

    \I__8838\ : Span4Mux_h
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__39627\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__8836\ : InMux
    port map (
            O => \N__39624\,
            I => \N__39620\
        );

    \I__8835\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39617\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__39620\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__39617\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__8832\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39607\
        );

    \I__8831\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39604\
        );

    \I__8830\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39601\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__39607\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__39604\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__39601\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__8826\ : InMux
    port map (
            O => \N__39594\,
            I => \N__39591\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__39591\,
            I => \N__39588\
        );

    \I__8824\ : Odrv12
    port map (
            O => \N__39588\,
            I => \pid_alt.O_0_4\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8822\ : InMux
    port map (
            O => \N__39582\,
            I => \N__39578\
        );

    \I__8821\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39575\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__39578\,
            I => \N__39572\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__39575\,
            I => \N__39569\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__39572\,
            I => \N__39566\
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__39569\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__39566\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__8815\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39558\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__8813\ : Odrv12
    port map (
            O => \N__39555\,
            I => \pid_alt.O_0_7\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__39552\,
            I => \N__39549\
        );

    \I__8811\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39546\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__39546\,
            I => \N__39543\
        );

    \I__8809\ : Span4Mux_h
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__39540\,
            I => \pid_alt.error_i_regZ0Z_3\
        );

    \I__8807\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__39534\,
            I => \uart_drone.CO0\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39531\,
            I => \N__39527\
        );

    \I__8804\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39524\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__39527\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__39524\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__39519\,
            I => \N__39513\
        );

    \I__8800\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39509\
        );

    \I__8799\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39504\
        );

    \I__8798\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39504\
        );

    \I__8797\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39497\
        );

    \I__8796\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39497\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__39509\,
            I => \N__39491\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__39504\,
            I => \N__39488\
        );

    \I__8793\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39483\
        );

    \I__8792\ : InMux
    port map (
            O => \N__39502\,
            I => \N__39483\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__39497\,
            I => \N__39480\
        );

    \I__8790\ : InMux
    port map (
            O => \N__39496\,
            I => \N__39477\
        );

    \I__8789\ : InMux
    port map (
            O => \N__39495\,
            I => \N__39474\
        );

    \I__8788\ : InMux
    port map (
            O => \N__39494\,
            I => \N__39471\
        );

    \I__8787\ : Span12Mux_h
    port map (
            O => \N__39491\,
            I => \N__39468\
        );

    \I__8786\ : Span12Mux_v
    port map (
            O => \N__39488\,
            I => \N__39463\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__39483\,
            I => \N__39463\
        );

    \I__8784\ : Span4Mux_v
    port map (
            O => \N__39480\,
            I => \N__39458\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__39477\,
            I => \N__39458\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39474\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__39471\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8780\ : Odrv12
    port map (
            O => \N__39468\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8779\ : Odrv12
    port map (
            O => \N__39463\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__39458\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8777\ : InMux
    port map (
            O => \N__39447\,
            I => \N__39444\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__39441\,
            I => \N__39438\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__39435\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__39429\,
            I => \N__39426\
        );

    \I__8770\ : Span4Mux_v
    port map (
            O => \N__39426\,
            I => \N__39423\
        );

    \I__8769\ : Span4Mux_h
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__39420\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__8767\ : InMux
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__39414\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__8765\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39408\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__39408\,
            I => \N__39405\
        );

    \I__8763\ : Span4Mux_v
    port map (
            O => \N__39405\,
            I => \N__39402\
        );

    \I__8762\ : Odrv4
    port map (
            O => \N__39402\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\
        );

    \I__8761\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39396\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__39396\,
            I => \N__39393\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__39393\,
            I => \N__39390\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__39390\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__39387\,
            I => \N__39382\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39386\,
            I => \N__39378\
        );

    \I__8755\ : InMux
    port map (
            O => \N__39385\,
            I => \N__39373\
        );

    \I__8754\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39373\
        );

    \I__8753\ : InMux
    port map (
            O => \N__39381\,
            I => \N__39370\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__39378\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__39373\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__39370\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39360\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__39360\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__8747\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39351\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39346\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39355\,
            I => \N__39346\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39343\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__39351\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__39346\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__39343\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__39333\,
            I => \N__39330\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8737\ : Span4Mux_v
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__39324\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39318\,
            I => \N__39315\
        );

    \I__8733\ : Span4Mux_v
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__39312\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__39309\,
            I => \N__39306\
        );

    \I__8730\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39303\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__8728\ : InMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__39297\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__8726\ : CascadeMux
    port map (
            O => \N__39294\,
            I => \N__39290\
        );

    \I__8725\ : InMux
    port map (
            O => \N__39293\,
            I => \N__39286\
        );

    \I__8724\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39283\
        );

    \I__8723\ : InMux
    port map (
            O => \N__39289\,
            I => \N__39280\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__39286\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39283\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__39280\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__8719\ : CascadeMux
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39267\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39267\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__8716\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39259\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39256\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39262\,
            I => \N__39253\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__39259\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__39256\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__39253\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__8710\ : InMux
    port map (
            O => \N__39246\,
            I => \N__39241\
        );

    \I__8709\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39238\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39244\,
            I => \N__39235\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__39241\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__39238\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__39235\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__39228\,
            I => \N__39224\
        );

    \I__8703\ : InMux
    port map (
            O => \N__39227\,
            I => \N__39219\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39224\,
            I => \N__39219\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__39219\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__8700\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39213\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__39213\,
            I => \N__39210\
        );

    \I__8698\ : Span4Mux_v
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__39207\,
            I => \N__39204\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__39204\,
            I => \N__39201\
        );

    \I__8695\ : Span4Mux_v
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__8694\ : Odrv4
    port map (
            O => \N__39198\,
            I => \pid_alt.un9_error_filt_2_9\
        );

    \I__8693\ : CascadeMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39192\,
            I => \N__39189\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__8690\ : Span12Mux_h
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__8689\ : Odrv12
    port map (
            O => \N__39183\,
            I => \pid_alt.un9_error_filt_add_1_cry_9_sZ0\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39180\,
            I => \pid_alt.un9_error_filt_add_1_cry_8\
        );

    \I__8687\ : CascadeMux
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39171\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39171\,
            I => \N__39168\
        );

    \I__8684\ : Span4Mux_h
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__8683\ : Span4Mux_h
    port map (
            O => \N__39165\,
            I => \N__39162\
        );

    \I__8682\ : Span4Mux_v
    port map (
            O => \N__39162\,
            I => \N__39159\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__39159\,
            I => \pid_alt.un9_error_filt_2_10\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39153\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39153\,
            I => \N__39150\
        );

    \I__8678\ : Span4Mux_s2_h
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__39147\,
            I => \N__39144\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__39144\,
            I => \N__39141\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__39141\,
            I => \N__39138\
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__39138\,
            I => \pid_alt.un9_error_filt_add_1_cry_10_sZ0\
        );

    \I__8673\ : InMux
    port map (
            O => \N__39135\,
            I => \pid_alt.un9_error_filt_add_1_cry_9\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__39132\,
            I => \N__39127\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39131\,
            I => \N__39115\
        );

    \I__8670\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39115\
        );

    \I__8669\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39115\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39115\
        );

    \I__8667\ : CascadeMux
    port map (
            O => \N__39125\,
            I => \N__39112\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__39124\,
            I => \N__39108\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__39115\,
            I => \N__39104\
        );

    \I__8664\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39095\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39095\
        );

    \I__8662\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39095\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39095\
        );

    \I__8660\ : Span4Mux_v
    port map (
            O => \N__39104\,
            I => \N__39090\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__39095\,
            I => \N__39090\
        );

    \I__8658\ : Span4Mux_h
    port map (
            O => \N__39090\,
            I => \N__39087\
        );

    \I__8657\ : Span4Mux_h
    port map (
            O => \N__39087\,
            I => \N__39084\
        );

    \I__8656\ : Odrv4
    port map (
            O => \N__39084\,
            I => \pid_alt.un9_error_filt_1_19\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39078\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__39078\,
            I => \N__39075\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__39075\,
            I => \N__39072\
        );

    \I__8652\ : Span4Mux_h
    port map (
            O => \N__39072\,
            I => \N__39069\
        );

    \I__8651\ : Span4Mux_v
    port map (
            O => \N__39069\,
            I => \N__39066\
        );

    \I__8650\ : Odrv4
    port map (
            O => \N__39066\,
            I => \pid_alt.un9_error_filt_2_11\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39063\,
            I => \pid_alt.un9_error_filt_add_1_cry_10\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__39060\,
            I => \N__39056\
        );

    \I__8647\ : InMux
    port map (
            O => \N__39059\,
            I => \N__39051\
        );

    \I__8646\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39051\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8644\ : Span12Mux_s10_h
    port map (
            O => \N__39048\,
            I => \N__39045\
        );

    \I__8643\ : Odrv12
    port map (
            O => \N__39045\,
            I => \pid_alt.un9_error_filt_add_1_sZ0Z_11\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39039\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__39039\,
            I => \N__39036\
        );

    \I__8640\ : Span4Mux_h
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8639\ : Odrv4
    port map (
            O => \N__39033\,
            I => \ppm_encoder_1.N_140_0\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39030\,
            I => \N__39026\
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__39029\,
            I => \N__39023\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__8635\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__8634\ : Span4Mux_v
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39017\,
            I => \N__39011\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__39014\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__8631\ : Odrv12
    port map (
            O => \N__39011\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39002\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39005\,
            I => \N__38998\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__39002\,
            I => \N__38995\
        );

    \I__8627\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38992\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__38998\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__38995\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__38992\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__38985\,
            I => \N__38980\
        );

    \I__8622\ : CascadeMux
    port map (
            O => \N__38984\,
            I => \N__38977\
        );

    \I__8621\ : InMux
    port map (
            O => \N__38983\,
            I => \N__38968\
        );

    \I__8620\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38965\
        );

    \I__8619\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38958\
        );

    \I__8618\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38958\
        );

    \I__8617\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38958\
        );

    \I__8616\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38953\
        );

    \I__8615\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38953\
        );

    \I__8614\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38950\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__38971\,
            I => \N__38942\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__38968\,
            I => \N__38939\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__38965\,
            I => \N__38932\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38932\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__38953\,
            I => \N__38932\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__38950\,
            I => \N__38929\
        );

    \I__8607\ : InMux
    port map (
            O => \N__38949\,
            I => \N__38926\
        );

    \I__8606\ : InMux
    port map (
            O => \N__38948\,
            I => \N__38922\
        );

    \I__8605\ : InMux
    port map (
            O => \N__38947\,
            I => \N__38919\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__38946\,
            I => \N__38913\
        );

    \I__8603\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38910\
        );

    \I__8602\ : InMux
    port map (
            O => \N__38942\,
            I => \N__38907\
        );

    \I__8601\ : Span4Mux_h
    port map (
            O => \N__38939\,
            I => \N__38898\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__38932\,
            I => \N__38898\
        );

    \I__8599\ : Span4Mux_h
    port map (
            O => \N__38929\,
            I => \N__38898\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38898\
        );

    \I__8597\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38895\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38892\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__38919\,
            I => \N__38889\
        );

    \I__8594\ : InMux
    port map (
            O => \N__38918\,
            I => \N__38886\
        );

    \I__8593\ : InMux
    port map (
            O => \N__38917\,
            I => \N__38879\
        );

    \I__8592\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38879\
        );

    \I__8591\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38879\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__38910\,
            I => \N__38876\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38869\
        );

    \I__8588\ : Span4Mux_v
    port map (
            O => \N__38898\,
            I => \N__38869\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__38895\,
            I => \N__38869\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__38892\,
            I => \N__38864\
        );

    \I__8585\ : Span4Mux_v
    port map (
            O => \N__38889\,
            I => \N__38864\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__38886\,
            I => \N__38861\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__38879\,
            I => \N__38852\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__38876\,
            I => \N__38852\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__38869\,
            I => \N__38849\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__38864\,
            I => \N__38844\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__38861\,
            I => \N__38844\
        );

    \I__8578\ : InMux
    port map (
            O => \N__38860\,
            I => \N__38841\
        );

    \I__8577\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38834\
        );

    \I__8576\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38834\
        );

    \I__8575\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38834\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__38852\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__38849\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__38844\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__38841\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__38834\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__8569\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__8567\ : Span4Mux_h
    port map (
            O => \N__38817\,
            I => \N__38814\
        );

    \I__8566\ : Span4Mux_v
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__8565\ : Odrv4
    port map (
            O => \N__38811\,
            I => \ppm_encoder_1.N_300\
        );

    \I__8564\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38805\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__8562\ : Span4Mux_v
    port map (
            O => \N__38802\,
            I => \N__38797\
        );

    \I__8561\ : InMux
    port map (
            O => \N__38801\,
            I => \N__38792\
        );

    \I__8560\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38792\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__38797\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__38792\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__38787\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__8556\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38781\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__38781\,
            I => \N__38778\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__38778\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__8553\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38772\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__38772\,
            I => \N__38769\
        );

    \I__8551\ : Span4Mux_h
    port map (
            O => \N__38769\,
            I => \N__38766\
        );

    \I__8550\ : Span4Mux_h
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__38763\,
            I => \pid_alt.un9_error_filt_1_17\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__38760\,
            I => \N__38757\
        );

    \I__8547\ : InMux
    port map (
            O => \N__38757\,
            I => \N__38754\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__38754\,
            I => \N__38751\
        );

    \I__8545\ : Span4Mux_h
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__8544\ : Span4Mux_h
    port map (
            O => \N__38748\,
            I => \N__38745\
        );

    \I__8543\ : Span4Mux_v
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__38742\,
            I => \pid_alt.un9_error_filt_2_2\
        );

    \I__8541\ : InMux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__8539\ : Span4Mux_s2_h
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__8538\ : Span4Mux_h
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__8537\ : Span4Mux_h
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__8536\ : Span4Mux_h
    port map (
            O => \N__38724\,
            I => \N__38721\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__38721\,
            I => \pid_alt.un9_error_filt_add_1_cry_2_sZ0\
        );

    \I__8534\ : InMux
    port map (
            O => \N__38718\,
            I => \pid_alt.un9_error_filt_add_1_cry_1\
        );

    \I__8533\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__38712\,
            I => \N__38709\
        );

    \I__8531\ : Span4Mux_h
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__8530\ : Span4Mux_h
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__38703\,
            I => \pid_alt.un9_error_filt_1_18\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__8527\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__8525\ : Span4Mux_h
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__8524\ : Span4Mux_h
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__8522\ : Odrv4
    port map (
            O => \N__38682\,
            I => \pid_alt.un9_error_filt_2_3\
        );

    \I__8521\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__8519\ : Span4Mux_s2_h
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__8518\ : Span4Mux_h
    port map (
            O => \N__38670\,
            I => \N__38667\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__38667\,
            I => \N__38664\
        );

    \I__8516\ : Span4Mux_h
    port map (
            O => \N__38664\,
            I => \N__38661\
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__38661\,
            I => \pid_alt.un9_error_filt_add_1_cry_3_sZ0\
        );

    \I__8514\ : InMux
    port map (
            O => \N__38658\,
            I => \pid_alt.un9_error_filt_add_1_cry_2\
        );

    \I__8513\ : CascadeMux
    port map (
            O => \N__38655\,
            I => \N__38652\
        );

    \I__8512\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__8510\ : Span12Mux_v
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8509\ : Odrv12
    port map (
            O => \N__38643\,
            I => \pid_alt.un9_error_filt_2_4\
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__8507\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__8505\ : Span12Mux_s9_h
    port map (
            O => \N__38631\,
            I => \N__38628\
        );

    \I__8504\ : Odrv12
    port map (
            O => \N__38628\,
            I => \pid_alt.un9_error_filt_add_1_cry_4_sZ0\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38625\,
            I => \pid_alt.un9_error_filt_add_1_cry_3\
        );

    \I__8502\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__38619\,
            I => \N__38616\
        );

    \I__8500\ : Span4Mux_h
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__8499\ : Span4Mux_h
    port map (
            O => \N__38613\,
            I => \N__38610\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__38607\,
            I => \pid_alt.un9_error_filt_2_5\
        );

    \I__8496\ : InMux
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__38601\,
            I => \N__38598\
        );

    \I__8494\ : Span12Mux_s8_h
    port map (
            O => \N__38598\,
            I => \N__38595\
        );

    \I__8493\ : Odrv12
    port map (
            O => \N__38595\,
            I => \pid_alt.un9_error_filt_add_1_cry_5_sZ0\
        );

    \I__8492\ : InMux
    port map (
            O => \N__38592\,
            I => \pid_alt.un9_error_filt_add_1_cry_4\
        );

    \I__8491\ : CascadeMux
    port map (
            O => \N__38589\,
            I => \N__38586\
        );

    \I__8490\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38583\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__38583\,
            I => \N__38580\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__38580\,
            I => \N__38577\
        );

    \I__8487\ : Span4Mux_h
    port map (
            O => \N__38577\,
            I => \N__38574\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__8485\ : Odrv4
    port map (
            O => \N__38571\,
            I => \pid_alt.un9_error_filt_2_6\
        );

    \I__8484\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38562\
        );

    \I__8482\ : Span4Mux_h
    port map (
            O => \N__38562\,
            I => \N__38559\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__38559\,
            I => \N__38556\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__38556\,
            I => \N__38553\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__38553\,
            I => \N__38550\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__38550\,
            I => \pid_alt.un9_error_filt_add_1_cry_6_sZ0\
        );

    \I__8477\ : InMux
    port map (
            O => \N__38547\,
            I => \pid_alt.un9_error_filt_add_1_cry_5\
        );

    \I__8476\ : InMux
    port map (
            O => \N__38544\,
            I => \N__38541\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__8474\ : Span4Mux_h
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__8473\ : Span4Mux_h
    port map (
            O => \N__38535\,
            I => \N__38532\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__38532\,
            I => \N__38529\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__38529\,
            I => \pid_alt.un9_error_filt_2_7\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__38526\,
            I => \N__38523\
        );

    \I__8469\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38520\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__38520\,
            I => \N__38517\
        );

    \I__8467\ : Span4Mux_h
    port map (
            O => \N__38517\,
            I => \N__38514\
        );

    \I__8466\ : Span4Mux_h
    port map (
            O => \N__38514\,
            I => \N__38511\
        );

    \I__8465\ : Span4Mux_h
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__8464\ : Span4Mux_h
    port map (
            O => \N__38508\,
            I => \N__38505\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__38505\,
            I => \pid_alt.un9_error_filt_add_1_cry_7_sZ0\
        );

    \I__8462\ : InMux
    port map (
            O => \N__38502\,
            I => \pid_alt.un9_error_filt_add_1_cry_6\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__38499\,
            I => \N__38496\
        );

    \I__8460\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__8456\ : Span4Mux_h
    port map (
            O => \N__38484\,
            I => \N__38481\
        );

    \I__8455\ : Span4Mux_v
    port map (
            O => \N__38481\,
            I => \N__38478\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__38478\,
            I => \pid_alt.un9_error_filt_2_8\
        );

    \I__8453\ : InMux
    port map (
            O => \N__38475\,
            I => \N__38472\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__38472\,
            I => \N__38469\
        );

    \I__8451\ : Span4Mux_s3_h
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__8450\ : Span4Mux_h
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__38463\,
            I => \N__38460\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__38460\,
            I => \N__38457\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__38457\,
            I => \pid_alt.un9_error_filt_add_1_cry_8_sZ0\
        );

    \I__8446\ : InMux
    port map (
            O => \N__38454\,
            I => \bfn_17_18_0_\
        );

    \I__8445\ : CascadeMux
    port map (
            O => \N__38451\,
            I => \N__38448\
        );

    \I__8444\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38445\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__38445\,
            I => \N__38442\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__38442\,
            I => \N__38439\
        );

    \I__8441\ : Span4Mux_h
    port map (
            O => \N__38439\,
            I => \N__38436\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__38436\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\
        );

    \I__8439\ : InMux
    port map (
            O => \N__38433\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__8438\ : InMux
    port map (
            O => \N__38430\,
            I => \bfn_17_16_0_\
        );

    \I__8437\ : InMux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__8434\ : Span4Mux_h
    port map (
            O => \N__38418\,
            I => \N__38415\
        );

    \I__8433\ : Odrv4
    port map (
            O => \N__38415\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__8432\ : InMux
    port map (
            O => \N__38412\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__8431\ : InMux
    port map (
            O => \N__38409\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38402\
        );

    \I__8429\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38398\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__38402\,
            I => \N__38395\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38392\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__38398\,
            I => \N__38387\
        );

    \I__8425\ : Span4Mux_v
    port map (
            O => \N__38395\,
            I => \N__38387\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__38392\,
            I => \N__38384\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__38387\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__8422\ : Odrv12
    port map (
            O => \N__38384\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__8421\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__38376\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__8419\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38369\
        );

    \I__8418\ : InMux
    port map (
            O => \N__38372\,
            I => \N__38366\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__38369\,
            I => \N__38363\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__38366\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__8415\ : Odrv4
    port map (
            O => \N__38363\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__8414\ : InMux
    port map (
            O => \N__38358\,
            I => \N__38355\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__38352\,
            I => \ppm_encoder_1.N_306\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38346\,
            I => \N__38343\
        );

    \I__8409\ : Span4Mux_h
    port map (
            O => \N__38343\,
            I => \N__38340\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__38337\,
            I => \pid_alt.un9_error_filt_1_15\
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__38334\,
            I => \N__38331\
        );

    \I__8405\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38328\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__8403\ : Span4Mux_v
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__8402\ : Span4Mux_h
    port map (
            O => \N__38322\,
            I => \N__38319\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__38316\,
            I => \N__38313\
        );

    \I__8399\ : Odrv4
    port map (
            O => \N__38313\,
            I => \pid_alt.un9_error_filt_2_0\
        );

    \I__8398\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38307\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__38307\,
            I => \N__38304\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__38304\,
            I => \N__38301\
        );

    \I__8395\ : Span4Mux_h
    port map (
            O => \N__38301\,
            I => \N__38298\
        );

    \I__8394\ : Span4Mux_h
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__8393\ : Span4Mux_h
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__8392\ : Odrv4
    port map (
            O => \N__38292\,
            I => \pid_alt.un9_error_filt_add_1_axbZ0Z_0\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__8389\ : Span4Mux_h
    port map (
            O => \N__38283\,
            I => \N__38280\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__8387\ : Odrv4
    port map (
            O => \N__38277\,
            I => \pid_alt.un9_error_filt_1_16\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__8383\ : Span4Mux_v
    port map (
            O => \N__38265\,
            I => \N__38262\
        );

    \I__8382\ : Span4Mux_h
    port map (
            O => \N__38262\,
            I => \N__38259\
        );

    \I__8381\ : Span4Mux_h
    port map (
            O => \N__38259\,
            I => \N__38256\
        );

    \I__8380\ : Span4Mux_v
    port map (
            O => \N__38256\,
            I => \N__38253\
        );

    \I__8379\ : Odrv4
    port map (
            O => \N__38253\,
            I => \pid_alt.un9_error_filt_2_1\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38247\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__38247\,
            I => \N__38244\
        );

    \I__8376\ : Span4Mux_s3_h
    port map (
            O => \N__38244\,
            I => \N__38241\
        );

    \I__8375\ : Span4Mux_h
    port map (
            O => \N__38241\,
            I => \N__38238\
        );

    \I__8374\ : Span4Mux_h
    port map (
            O => \N__38238\,
            I => \N__38235\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__38235\,
            I => \N__38232\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__38232\,
            I => \pid_alt.un9_error_filt_add_1_cry_1_sZ0\
        );

    \I__8371\ : InMux
    port map (
            O => \N__38229\,
            I => \pid_alt.un9_error_filt_add_1_cry_0\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__38223\,
            I => \N__38220\
        );

    \I__8368\ : Span4Mux_h
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__38217\,
            I => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38214\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__8365\ : InMux
    port map (
            O => \N__38211\,
            I => \N__38208\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__38208\,
            I => \N__38205\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__38205\,
            I => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38202\,
            I => \bfn_17_15_0_\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38196\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__38193\,
            I => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38190\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__38184\,
            I => \N__38181\
        );

    \I__8355\ : Span4Mux_h
    port map (
            O => \N__38181\,
            I => \N__38178\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__38178\,
            I => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38172\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38172\,
            I => \N__38169\
        );

    \I__8351\ : Odrv4
    port map (
            O => \N__38169\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38166\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__8349\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38160\,
            I => \N__38157\
        );

    \I__8347\ : Span4Mux_h
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__38154\,
            I => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__38151\,
            I => \N__38148\
        );

    \I__8344\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38145\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38141\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38138\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__38141\,
            I => \N__38135\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38138\,
            I => \N__38132\
        );

    \I__8339\ : Span4Mux_v
    port map (
            O => \N__38135\,
            I => \N__38129\
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__38132\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__8337\ : Odrv4
    port map (
            O => \N__38129\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__8336\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38121\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__38121\,
            I => \N__38118\
        );

    \I__8334\ : Odrv4
    port map (
            O => \N__38118\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__8333\ : InMux
    port map (
            O => \N__38115\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__8332\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38109\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38106\
        );

    \I__8330\ : Span4Mux_v
    port map (
            O => \N__38106\,
            I => \N__38103\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__38103\,
            I => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__38100\,
            I => \N__38097\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38093\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38090\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38093\,
            I => \N__38087\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38090\,
            I => \N__38084\
        );

    \I__8323\ : Span12Mux_v
    port map (
            O => \N__38087\,
            I => \N__38081\
        );

    \I__8322\ : Odrv12
    port map (
            O => \N__38084\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__8321\ : Odrv12
    port map (
            O => \N__38081\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__8320\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38073\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__38073\,
            I => \N__38070\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__38070\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38067\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__8316\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38061\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__8314\ : Span4Mux_v
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__8313\ : Odrv4
    port map (
            O => \N__38055\,
            I => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__38052\,
            I => \N__38049\
        );

    \I__8311\ : InMux
    port map (
            O => \N__38049\,
            I => \N__38046\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__38046\,
            I => \N__38042\
        );

    \I__8309\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38039\
        );

    \I__8308\ : Span4Mux_h
    port map (
            O => \N__38042\,
            I => \N__38036\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38039\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__8306\ : Odrv4
    port map (
            O => \N__38036\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__8305\ : InMux
    port map (
            O => \N__38031\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__38022\,
            I => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38019\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__8300\ : InMux
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__8298\ : Span4Mux_v
    port map (
            O => \N__38010\,
            I => \N__38007\
        );

    \I__8297\ : Odrv4
    port map (
            O => \N__38007\,
            I => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__8295\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37997\
        );

    \I__8294\ : InMux
    port map (
            O => \N__38000\,
            I => \N__37994\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__37997\,
            I => \N__37991\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__37994\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__8291\ : Odrv12
    port map (
            O => \N__37991\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__8290\ : InMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__8288\ : Span4Mux_h
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__8287\ : Odrv4
    port map (
            O => \N__37977\,
            I => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__37974\,
            I => \N__37970\
        );

    \I__8285\ : InMux
    port map (
            O => \N__37973\,
            I => \N__37967\
        );

    \I__8284\ : InMux
    port map (
            O => \N__37970\,
            I => \N__37964\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__37967\,
            I => \N__37961\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37958\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__37961\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__8280\ : Odrv4
    port map (
            O => \N__37958\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__8279\ : CascadeMux
    port map (
            O => \N__37953\,
            I => \N__37950\
        );

    \I__8278\ : InMux
    port map (
            O => \N__37950\,
            I => \N__37947\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__37947\,
            I => \N__37944\
        );

    \I__8276\ : Odrv4
    port map (
            O => \N__37944\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__8275\ : InMux
    port map (
            O => \N__37941\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__8274\ : InMux
    port map (
            O => \N__37938\,
            I => \N__37935\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__37935\,
            I => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__8271\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37925\
        );

    \I__8270\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37922\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__37925\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__37922\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__8267\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37914\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__37914\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__8265\ : InMux
    port map (
            O => \N__37911\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__8264\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__37905\,
            I => \ppm_encoder_1.throttle_RNI82223Z0Z_3\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__37902\,
            I => \N__37899\
        );

    \I__8261\ : InMux
    port map (
            O => \N__37899\,
            I => \N__37895\
        );

    \I__8260\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37892\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__37895\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__37892\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__8257\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__37884\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__8255\ : InMux
    port map (
            O => \N__37881\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__8254\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__37875\,
            I => \N__37872\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__37872\,
            I => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__37869\,
            I => \N__37866\
        );

    \I__8250\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37862\
        );

    \I__8249\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37859\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37856\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__37859\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__8246\ : Odrv12
    port map (
            O => \N__37856\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__8245\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37845\
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__37845\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__8242\ : InMux
    port map (
            O => \N__37842\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__8241\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__37836\,
            I => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\
        );

    \I__8239\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37829\
        );

    \I__8238\ : CascadeMux
    port map (
            O => \N__37832\,
            I => \N__37826\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__37829\,
            I => \N__37823\
        );

    \I__8236\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37820\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__37823\,
            I => \N__37817\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__37820\,
            I => \N__37814\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__37817\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__8232\ : Odrv12
    port map (
            O => \N__37814\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__8231\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37806\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__37806\,
            I => \N__37803\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__37803\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__8228\ : InMux
    port map (
            O => \N__37800\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__8227\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37794\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__8225\ : Odrv4
    port map (
            O => \N__37791\,
            I => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__37788\,
            I => \N__37784\
        );

    \I__8223\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37781\
        );

    \I__8222\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37778\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37781\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__37778\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__8219\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__37770\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__8217\ : InMux
    port map (
            O => \N__37767\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__8216\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37757\
        );

    \I__8215\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37757\
        );

    \I__8214\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37754\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37751\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__37754\,
            I => \N__37746\
        );

    \I__8211\ : Sp12to4
    port map (
            O => \N__37751\,
            I => \N__37746\
        );

    \I__8210\ : Span12Mux_v
    port map (
            O => \N__37746\,
            I => \N__37743\
        );

    \I__8209\ : Odrv12
    port map (
            O => \N__37743\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__8208\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37735\
        );

    \I__8207\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37730\
        );

    \I__8206\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37730\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__37735\,
            I => \N__37725\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__37730\,
            I => \N__37725\
        );

    \I__8203\ : Span12Mux_v
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__8202\ : Odrv12
    port map (
            O => \N__37722\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__37719\,
            I => \N__37714\
        );

    \I__8200\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37705\
        );

    \I__8199\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37705\
        );

    \I__8198\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37705\
        );

    \I__8197\ : InMux
    port map (
            O => \N__37713\,
            I => \N__37700\
        );

    \I__8196\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37697\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37694\
        );

    \I__8194\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37691\
        );

    \I__8193\ : CascadeMux
    port map (
            O => \N__37703\,
            I => \N__37688\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__37700\,
            I => \N__37683\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__37697\,
            I => \N__37680\
        );

    \I__8190\ : Span4Mux_h
    port map (
            O => \N__37694\,
            I => \N__37675\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37675\
        );

    \I__8188\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37670\
        );

    \I__8187\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37670\
        );

    \I__8186\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37667\
        );

    \I__8185\ : Span12Mux_s10_h
    port map (
            O => \N__37683\,
            I => \N__37662\
        );

    \I__8184\ : Sp12to4
    port map (
            O => \N__37680\,
            I => \N__37662\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__37675\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__37670\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__37667\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__8180\ : Odrv12
    port map (
            O => \N__37662\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__8179\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37647\
        );

    \I__8178\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37642\
        );

    \I__8177\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37642\
        );

    \I__8176\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37639\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__37647\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__37642\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__37639\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8172\ : CascadeMux
    port map (
            O => \N__37632\,
            I => \N__37627\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__37631\,
            I => \N__37624\
        );

    \I__8170\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37621\
        );

    \I__8169\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37618\
        );

    \I__8168\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37615\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__37621\,
            I => \N__37612\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__37618\,
            I => \N__37609\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__37615\,
            I => \N__37604\
        );

    \I__8164\ : Span4Mux_v
    port map (
            O => \N__37612\,
            I => \N__37604\
        );

    \I__8163\ : Span4Mux_h
    port map (
            O => \N__37609\,
            I => \N__37601\
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__37604\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__8161\ : Odrv4
    port map (
            O => \N__37601\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__8160\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__37593\,
            I => \N__37587\
        );

    \I__8158\ : InMux
    port map (
            O => \N__37592\,
            I => \N__37584\
        );

    \I__8157\ : InMux
    port map (
            O => \N__37591\,
            I => \N__37578\
        );

    \I__8156\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37575\
        );

    \I__8155\ : Span4Mux_h
    port map (
            O => \N__37587\,
            I => \N__37569\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37569\
        );

    \I__8153\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37565\
        );

    \I__8152\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37562\
        );

    \I__8151\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37559\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__37578\,
            I => \N__37554\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__37575\,
            I => \N__37554\
        );

    \I__8148\ : InMux
    port map (
            O => \N__37574\,
            I => \N__37545\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__37569\,
            I => \N__37542\
        );

    \I__8146\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37539\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37530\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__37562\,
            I => \N__37530\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37530\
        );

    \I__8142\ : Span4Mux_v
    port map (
            O => \N__37554\,
            I => \N__37530\
        );

    \I__8141\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37525\
        );

    \I__8140\ : InMux
    port map (
            O => \N__37552\,
            I => \N__37525\
        );

    \I__8139\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37518\
        );

    \I__8138\ : InMux
    port map (
            O => \N__37550\,
            I => \N__37518\
        );

    \I__8137\ : InMux
    port map (
            O => \N__37549\,
            I => \N__37518\
        );

    \I__8136\ : InMux
    port map (
            O => \N__37548\,
            I => \N__37515\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__37545\,
            I => \N__37512\
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__37542\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__37539\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__37530\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__37525\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__37518\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__37515\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8128\ : Odrv4
    port map (
            O => \N__37512\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__8127\ : CascadeMux
    port map (
            O => \N__37497\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\
        );

    \I__8126\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37491\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__8124\ : Span4Mux_v
    port map (
            O => \N__37488\,
            I => \N__37483\
        );

    \I__8123\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37480\
        );

    \I__8122\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37477\
        );

    \I__8121\ : Odrv4
    port map (
            O => \N__37483\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__37480\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__37477\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__8118\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37461\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37461\
        );

    \I__8116\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37461\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37461\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__37455\,
            I => \N__37451\
        );

    \I__8112\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37448\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__37451\,
            I => \N__37443\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37443\
        );

    \I__8109\ : Odrv4
    port map (
            O => \N__37443\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__8108\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37437\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__37431\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__8104\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37419\
        );

    \I__8103\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37419\
        );

    \I__8102\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37419\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__37419\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__8100\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37413\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__37413\,
            I => \N__37409\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37406\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__37409\,
            I => \N__37401\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37401\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__37401\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37395\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__8092\ : Span4Mux_v
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__37389\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37386\,
            I => \N__37381\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37376\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37376\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__37381\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__37376\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__8085\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37367\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37364\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__37367\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__37364\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__8081\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37355\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37352\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37355\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37352\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__8077\ : CascadeMux
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37340\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37337\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37340\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37337\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37328\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37325\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__37328\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__37325\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37314\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37311\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37308\
        );

    \I__8065\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37305\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37314\,
            I => \N__37302\
        );

    \I__8063\ : LocalMux
    port map (
            O => \N__37311\,
            I => \N__37299\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__37308\,
            I => \N__37294\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__37305\,
            I => \N__37294\
        );

    \I__8060\ : Span4Mux_h
    port map (
            O => \N__37302\,
            I => \N__37291\
        );

    \I__8059\ : Span4Mux_h
    port map (
            O => \N__37299\,
            I => \N__37288\
        );

    \I__8058\ : Span4Mux_h
    port map (
            O => \N__37294\,
            I => \N__37285\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__37291\,
            I => \N__37282\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__37288\,
            I => \reset_module_System.reset6_14\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__37285\,
            I => \reset_module_System.reset6_14\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__37282\,
            I => \reset_module_System.reset6_14\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37272\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__37272\,
            I => \ppm_encoder_1.un1_init_pulses_10_0\
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__37269\,
            I => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\
        );

    \I__8050\ : CascadeMux
    port map (
            O => \N__37266\,
            I => \ppm_encoder_1.un1_init_pulses_0_cascade_\
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__37263\,
            I => \N__37251\
        );

    \I__8048\ : CascadeMux
    port map (
            O => \N__37262\,
            I => \N__37247\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__37261\,
            I => \N__37244\
        );

    \I__8046\ : CascadeMux
    port map (
            O => \N__37260\,
            I => \N__37237\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__37259\,
            I => \N__37234\
        );

    \I__8044\ : CascadeMux
    port map (
            O => \N__37258\,
            I => \N__37228\
        );

    \I__8043\ : CascadeMux
    port map (
            O => \N__37257\,
            I => \N__37221\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__37256\,
            I => \N__37218\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \N__37215\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37207\
        );

    \I__8039\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37207\
        );

    \I__8038\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37207\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37204\
        );

    \I__8036\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37200\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__37243\,
            I => \N__37197\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__37242\,
            I => \N__37194\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__37241\,
            I => \N__37188\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37240\,
            I => \N__37181\
        );

    \I__8031\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37181\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37181\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37172\
        );

    \I__8028\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37172\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37172\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37228\,
            I => \N__37172\
        );

    \I__8025\ : CascadeMux
    port map (
            O => \N__37227\,
            I => \N__37169\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__37226\,
            I => \N__37166\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37225\,
            I => \N__37158\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37158\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37158\
        );

    \I__8020\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37151\
        );

    \I__8019\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37151\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37151\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__37207\,
            I => \N__37142\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__37204\,
            I => \N__37142\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37139\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37136\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37197\,
            I => \N__37129\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37129\
        );

    \I__8011\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37129\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37192\,
            I => \N__37122\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37122\
        );

    \I__8008\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37122\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37117\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37117\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37110\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37110\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37110\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__37158\,
            I => \N__37105\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__37151\,
            I => \N__37105\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__37150\,
            I => \N__37099\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__37149\,
            I => \N__37096\
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__37148\,
            I => \N__37093\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__37147\,
            I => \N__37086\
        );

    \I__7996\ : Span4Mux_v
    port map (
            O => \N__37142\,
            I => \N__37083\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__37139\,
            I => \N__37080\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__37136\,
            I => \N__37071\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__37129\,
            I => \N__37071\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37071\
        );

    \I__7991\ : Span4Mux_v
    port map (
            O => \N__37117\,
            I => \N__37071\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__37110\,
            I => \N__37068\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__37105\,
            I => \N__37065\
        );

    \I__7988\ : InMux
    port map (
            O => \N__37104\,
            I => \N__37054\
        );

    \I__7987\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37054\
        );

    \I__7986\ : InMux
    port map (
            O => \N__37102\,
            I => \N__37054\
        );

    \I__7985\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37054\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37054\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37047\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37047\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37047\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37090\,
            I => \N__37040\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37089\,
            I => \N__37040\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37086\,
            I => \N__37040\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__37083\,
            I => \N__37037\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__37080\,
            I => \N__37032\
        );

    \I__7975\ : Span4Mux_v
    port map (
            O => \N__37071\,
            I => \N__37032\
        );

    \I__7974\ : Sp12to4
    port map (
            O => \N__37068\,
            I => \N__37029\
        );

    \I__7973\ : Span4Mux_h
    port map (
            O => \N__37065\,
            I => \N__37026\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__37054\,
            I => \N__37021\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__37047\,
            I => \N__37021\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37040\,
            I => \N__37012\
        );

    \I__7969\ : Sp12to4
    port map (
            O => \N__37037\,
            I => \N__37012\
        );

    \I__7968\ : Sp12to4
    port map (
            O => \N__37032\,
            I => \N__37012\
        );

    \I__7967\ : Span12Mux_v
    port map (
            O => \N__37029\,
            I => \N__37012\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__37026\,
            I => \N__37009\
        );

    \I__7965\ : Span12Mux_v
    port map (
            O => \N__37021\,
            I => \N__37006\
        );

    \I__7964\ : Span12Mux_h
    port map (
            O => \N__37012\,
            I => \N__37003\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__37009\,
            I => pid_altitude_dv
        );

    \I__7962\ : Odrv12
    port map (
            O => \N__37006\,
            I => pid_altitude_dv
        );

    \I__7961\ : Odrv12
    port map (
            O => \N__37003\,
            I => pid_altitude_dv
        );

    \I__7960\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36989\
        );

    \I__7958\ : CascadeMux
    port map (
            O => \N__36992\,
            I => \N__36985\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__36989\,
            I => \N__36982\
        );

    \I__7956\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36979\
        );

    \I__7955\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36976\
        );

    \I__7954\ : Span4Mux_h
    port map (
            O => \N__36982\,
            I => \N__36971\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__36979\,
            I => \N__36971\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__36976\,
            I => throttle_command_0
        );

    \I__7951\ : Odrv4
    port map (
            O => \N__36971\,
            I => throttle_command_0
        );

    \I__7950\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36960\
        );

    \I__7949\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36957\
        );

    \I__7948\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36952\
        );

    \I__7947\ : InMux
    port map (
            O => \N__36963\,
            I => \N__36952\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__36960\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__36957\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__36952\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__7942\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36936\
        );

    \I__7941\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36933\
        );

    \I__7940\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36928\
        );

    \I__7939\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36928\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__36936\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__36933\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__36928\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__7935\ : InMux
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__36915\,
            I => \N__36912\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__36912\,
            I => \N__36909\
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__36909\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\
        );

    \I__7930\ : InMux
    port map (
            O => \N__36906\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__7929\ : SRMux
    port map (
            O => \N__36903\,
            I => \N__36894\
        );

    \I__7928\ : SRMux
    port map (
            O => \N__36902\,
            I => \N__36894\
        );

    \I__7927\ : SRMux
    port map (
            O => \N__36901\,
            I => \N__36894\
        );

    \I__7926\ : GlobalMux
    port map (
            O => \N__36894\,
            I => \N__36891\
        );

    \I__7925\ : gio2CtrlBuf
    port map (
            O => \N__36891\,
            I => \ppm_encoder_1.N_322_g\
        );

    \I__7924\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36884\
        );

    \I__7923\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36881\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36877\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36874\
        );

    \I__7920\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36868\
        );

    \I__7919\ : Span4Mux_h
    port map (
            O => \N__36877\,
            I => \N__36861\
        );

    \I__7918\ : Span4Mux_v
    port map (
            O => \N__36874\,
            I => \N__36858\
        );

    \I__7917\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36852\
        );

    \I__7916\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36849\
        );

    \I__7915\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36846\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36843\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__36867\,
            I => \N__36840\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__36866\,
            I => \N__36835\
        );

    \I__7911\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36832\
        );

    \I__7910\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36829\
        );

    \I__7909\ : Sp12to4
    port map (
            O => \N__36861\,
            I => \N__36826\
        );

    \I__7908\ : Sp12to4
    port map (
            O => \N__36858\,
            I => \N__36823\
        );

    \I__7907\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36820\
        );

    \I__7906\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36816\
        );

    \I__7905\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36813\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__36852\,
            I => \N__36810\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__36849\,
            I => \N__36807\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__36846\,
            I => \N__36802\
        );

    \I__7901\ : Span12Mux_s10_v
    port map (
            O => \N__36843\,
            I => \N__36802\
        );

    \I__7900\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36799\
        );

    \I__7899\ : InMux
    port map (
            O => \N__36839\,
            I => \N__36792\
        );

    \I__7898\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36792\
        );

    \I__7897\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36792\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36781\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__36829\,
            I => \N__36781\
        );

    \I__7894\ : Span12Mux_s10_v
    port map (
            O => \N__36826\,
            I => \N__36781\
        );

    \I__7893\ : Span12Mux_h
    port map (
            O => \N__36823\,
            I => \N__36781\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__36820\,
            I => \N__36781\
        );

    \I__7891\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36778\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__36816\,
            I => \N__36769\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__36813\,
            I => \N__36769\
        );

    \I__7888\ : Span4Mux_v
    port map (
            O => \N__36810\,
            I => \N__36769\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__36807\,
            I => \N__36769\
        );

    \I__7886\ : Span12Mux_v
    port map (
            O => \N__36802\,
            I => \N__36766\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__36799\,
            I => \N__36759\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36759\
        );

    \I__7883\ : Span12Mux_v
    port map (
            O => \N__36781\,
            I => \N__36759\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__36778\,
            I => uart_pc_data_2
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__36769\,
            I => uart_pc_data_2
        );

    \I__7880\ : Odrv12
    port map (
            O => \N__36766\,
            I => uart_pc_data_2
        );

    \I__7879\ : Odrv12
    port map (
            O => \N__36759\,
            I => uart_pc_data_2
        );

    \I__7878\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__36747\,
            I => \N__36744\
        );

    \I__7876\ : Span12Mux_s9_h
    port map (
            O => \N__36744\,
            I => \N__36741\
        );

    \I__7875\ : Odrv12
    port map (
            O => \N__36741\,
            I => alt_ki_2
        );

    \I__7874\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36735\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__7872\ : Odrv12
    port map (
            O => \N__36732\,
            I => \pid_alt.O_0_6\
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__36729\,
            I => \N__36726\
        );

    \I__7870\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36723\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__36723\,
            I => \N__36720\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__36717\,
            I => \pid_alt.error_i_regZ0Z_2\
        );

    \I__7866\ : CascadeMux
    port map (
            O => \N__36714\,
            I => \N__36711\
        );

    \I__7865\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36707\
        );

    \I__7864\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36704\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__36707\,
            I => \N__36699\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__36704\,
            I => \N__36699\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__36699\,
            I => \N__36696\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__36696\,
            I => \uart_drone.N_144_1\
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__36693\,
            I => \N__36688\
        );

    \I__7858\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36683\
        );

    \I__7857\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36680\
        );

    \I__7856\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36672\
        );

    \I__7855\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36672\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__36686\,
            I => \N__36668\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__36683\,
            I => \N__36663\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__36680\,
            I => \N__36663\
        );

    \I__7851\ : InMux
    port map (
            O => \N__36679\,
            I => \N__36660\
        );

    \I__7850\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36655\
        );

    \I__7849\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36655\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36652\
        );

    \I__7847\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36649\
        );

    \I__7846\ : InMux
    port map (
            O => \N__36668\,
            I => \N__36646\
        );

    \I__7845\ : Span4Mux_v
    port map (
            O => \N__36663\,
            I => \N__36641\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__36660\,
            I => \N__36641\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__36655\,
            I => \N__36638\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__36652\,
            I => \N__36633\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__36649\,
            I => \N__36633\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__36646\,
            I => \N__36626\
        );

    \I__7839\ : Span4Mux_h
    port map (
            O => \N__36641\,
            I => \N__36626\
        );

    \I__7838\ : Span4Mux_v
    port map (
            O => \N__36638\,
            I => \N__36626\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__36633\,
            I => \N__36623\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__36626\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__36623\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__7834\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36612\
        );

    \I__7833\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36609\
        );

    \I__7832\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36601\
        );

    \I__7831\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36598\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__36612\,
            I => \N__36595\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36592\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__36608\,
            I => \N__36589\
        );

    \I__7827\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36586\
        );

    \I__7826\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36583\
        );

    \I__7825\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36580\
        );

    \I__7824\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36577\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__36601\,
            I => \N__36572\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__36598\,
            I => \N__36572\
        );

    \I__7821\ : Span4Mux_v
    port map (
            O => \N__36595\,
            I => \N__36567\
        );

    \I__7820\ : Span4Mux_v
    port map (
            O => \N__36592\,
            I => \N__36567\
        );

    \I__7819\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36564\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__36586\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__36583\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__36580\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__36577\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7814\ : Odrv4
    port map (
            O => \N__36572\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__36567\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__36564\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7811\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36546\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__36546\,
            I => \N__36541\
        );

    \I__7809\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36538\
        );

    \I__7808\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36532\
        );

    \I__7807\ : Span4Mux_v
    port map (
            O => \N__36541\,
            I => \N__36526\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__36538\,
            I => \N__36526\
        );

    \I__7805\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36522\
        );

    \I__7804\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36519\
        );

    \I__7803\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36516\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36513\
        );

    \I__7801\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36510\
        );

    \I__7800\ : Span4Mux_h
    port map (
            O => \N__36526\,
            I => \N__36507\
        );

    \I__7799\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36504\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__36522\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__36519\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__36516\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7795\ : Odrv4
    port map (
            O => \N__36513\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__36510\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__36507\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__36504\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7791\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36485\
        );

    \I__7790\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36480\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__36485\,
            I => \N__36477\
        );

    \I__7788\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36472\
        );

    \I__7787\ : InMux
    port map (
            O => \N__36483\,
            I => \N__36469\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__36480\,
            I => \N__36464\
        );

    \I__7785\ : Span4Mux_h
    port map (
            O => \N__36477\,
            I => \N__36464\
        );

    \I__7784\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36459\
        );

    \I__7783\ : InMux
    port map (
            O => \N__36475\,
            I => \N__36459\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__36472\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36469\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__36464\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__36459\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__36450\,
            I => \uart_drone.un1_state_4_0_cascade_\
        );

    \I__7777\ : InMux
    port map (
            O => \N__36447\,
            I => \bfn_16_20_0_\
        );

    \I__7776\ : InMux
    port map (
            O => \N__36444\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__7775\ : InMux
    port map (
            O => \N__36441\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__7774\ : InMux
    port map (
            O => \N__36438\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__7773\ : InMux
    port map (
            O => \N__36435\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__7772\ : InMux
    port map (
            O => \N__36432\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__7771\ : InMux
    port map (
            O => \N__36429\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36426\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__7769\ : InMux
    port map (
            O => \N__36423\,
            I => \bfn_16_21_0_\
        );

    \I__7768\ : InMux
    port map (
            O => \N__36420\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__36417\,
            I => \N__36413\
        );

    \I__7766\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36410\
        );

    \I__7765\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36407\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__36404\,
            I => \N__36396\
        );

    \I__7761\ : Span4Mux_v
    port map (
            O => \N__36401\,
            I => \N__36396\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__36396\,
            I => \ppm_encoder_1.N_1330_i\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__36393\,
            I => \N__36388\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36392\,
            I => \N__36385\
        );

    \I__7757\ : InMux
    port map (
            O => \N__36391\,
            I => \N__36382\
        );

    \I__7756\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36379\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__36385\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__36382\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__36379\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36366\
        );

    \I__7751\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36361\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36361\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36358\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36366\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__36361\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__36358\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__7745\ : InMux
    port map (
            O => \N__36351\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__7744\ : InMux
    port map (
            O => \N__36348\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__7743\ : InMux
    port map (
            O => \N__36345\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36337\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36334\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36331\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__36337\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__36334\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36331\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36324\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36316\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36313\
        );

    \I__7733\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36310\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__36316\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__36313\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36310\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36303\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__7728\ : InMux
    port map (
            O => \N__36300\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36297\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36291\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__36291\,
            I => \N__36287\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36290\,
            I => \N__36284\
        );

    \I__7723\ : Odrv12
    port map (
            O => \N__36287\,
            I => scaler_4_data_13
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__36284\,
            I => scaler_4_data_13
        );

    \I__7721\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__36276\,
            I => \N__36273\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__36273\,
            I => \N__36270\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__36270\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__7717\ : CEMux
    port map (
            O => \N__36267\,
            I => \N__36263\
        );

    \I__7716\ : CEMux
    port map (
            O => \N__36266\,
            I => \N__36259\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__36263\,
            I => \N__36256\
        );

    \I__7714\ : CEMux
    port map (
            O => \N__36262\,
            I => \N__36253\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36259\,
            I => \N__36250\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__36256\,
            I => \N__36245\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__36253\,
            I => \N__36245\
        );

    \I__7710\ : Span4Mux_v
    port map (
            O => \N__36250\,
            I => \N__36241\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__36245\,
            I => \N__36238\
        );

    \I__7708\ : CEMux
    port map (
            O => \N__36244\,
            I => \N__36235\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__36241\,
            I => \N__36228\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__36238\,
            I => \N__36228\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__36235\,
            I => \N__36228\
        );

    \I__7704\ : Span4Mux_h
    port map (
            O => \N__36228\,
            I => \N__36224\
        );

    \I__7703\ : CEMux
    port map (
            O => \N__36227\,
            I => \N__36221\
        );

    \I__7702\ : Odrv4
    port map (
            O => \N__36224\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__36221\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__36216\,
            I => \N__36213\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36213\,
            I => \N__36209\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36206\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__36209\,
            I => \N__36202\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N__36199\
        );

    \I__7695\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36196\
        );

    \I__7694\ : Span4Mux_v
    port map (
            O => \N__36202\,
            I => \N__36191\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__36199\,
            I => \N__36191\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__36196\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__36191\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36186\,
            I => \N__36182\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36179\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__36182\,
            I => \N__36176\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__36179\,
            I => \N__36173\
        );

    \I__7686\ : Span4Mux_v
    port map (
            O => \N__36176\,
            I => \N__36170\
        );

    \I__7685\ : Span4Mux_h
    port map (
            O => \N__36173\,
            I => \N__36167\
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__36170\,
            I => scaler_2_data_11
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__36167\,
            I => scaler_2_data_11
        );

    \I__7682\ : InMux
    port map (
            O => \N__36162\,
            I => \N__36159\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__36159\,
            I => \N__36156\
        );

    \I__7680\ : Odrv4
    port map (
            O => \N__36156\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36150\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__36150\,
            I => \N__36145\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36142\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36139\
        );

    \I__7675\ : Span4Mux_h
    port map (
            O => \N__36145\,
            I => \N__36136\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36142\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__36139\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__36136\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36126\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36123\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__36123\,
            I => \N__36120\
        );

    \I__7668\ : Odrv4
    port map (
            O => \N__36120\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36114\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__7665\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36108\,
            I => \N__36105\
        );

    \I__7663\ : Span12Mux_v
    port map (
            O => \N__36105\,
            I => \N__36102\
        );

    \I__7662\ : Odrv12
    port map (
            O => \N__36102\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__7660\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__36093\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__7658\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__7656\ : Odrv12
    port map (
            O => \N__36084\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36078\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__36078\,
            I => \N__36075\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__36075\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36069\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__36069\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36066\,
            I => \N__36063\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__36063\,
            I => \N__36060\
        );

    \I__7648\ : Odrv12
    port map (
            O => \N__36060\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36054\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36054\,
            I => \N__36051\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__36051\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36048\,
            I => \N__36044\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36041\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__36044\,
            I => \N__36038\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36035\
        );

    \I__7640\ : Span4Mux_v
    port map (
            O => \N__36038\,
            I => \N__36032\
        );

    \I__7639\ : Odrv4
    port map (
            O => \N__36035\,
            I => scaler_2_data_8
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__36032\,
            I => scaler_2_data_8
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__36027\,
            I => \N__36024\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36024\,
            I => \N__36021\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__36021\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36018\,
            I => \ppm_encoder_1.un1_aileron_cry_7\
        );

    \I__7633\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36011\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36008\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36011\,
            I => \N__36005\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__36000\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__36005\,
            I => \N__36000\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__36000\,
            I => scaler_2_data_9
        );

    \I__7627\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35994\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__35994\,
            I => \N__35991\
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__35991\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__7624\ : InMux
    port map (
            O => \N__35988\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__7623\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35981\
        );

    \I__7622\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35978\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__35981\,
            I => \N__35975\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__35978\,
            I => \N__35972\
        );

    \I__7619\ : Span4Mux_v
    port map (
            O => \N__35975\,
            I => \N__35967\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__35972\,
            I => \N__35967\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__35967\,
            I => scaler_2_data_10
        );

    \I__7616\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35961\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__35961\,
            I => \N__35958\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__35958\,
            I => \N__35955\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__35955\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__7612\ : InMux
    port map (
            O => \N__35952\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__7611\ : InMux
    port map (
            O => \N__35949\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__7610\ : InMux
    port map (
            O => \N__35946\,
            I => \N__35942\
        );

    \I__7609\ : InMux
    port map (
            O => \N__35945\,
            I => \N__35939\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__35942\,
            I => \N__35936\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__35939\,
            I => \N__35933\
        );

    \I__7606\ : Span4Mux_h
    port map (
            O => \N__35936\,
            I => \N__35930\
        );

    \I__7605\ : Span4Mux_h
    port map (
            O => \N__35933\,
            I => \N__35927\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__35930\,
            I => scaler_2_data_12
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__35927\,
            I => scaler_2_data_12
        );

    \I__7602\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__35919\,
            I => \N__35916\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__35916\,
            I => \N__35913\
        );

    \I__7599\ : Odrv4
    port map (
            O => \N__35913\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__7598\ : InMux
    port map (
            O => \N__35910\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__35907\,
            I => \N__35903\
        );

    \I__7596\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35900\
        );

    \I__7595\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35897\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35894\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__35897\,
            I => \N__35891\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__35894\,
            I => \N__35888\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__35891\,
            I => scaler_2_data_13
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__35888\,
            I => scaler_2_data_13
        );

    \I__7589\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35880\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__35880\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__7587\ : InMux
    port map (
            O => \N__35877\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__7586\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35871\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__35871\,
            I => \N__35868\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__35868\,
            I => \N__35865\
        );

    \I__7583\ : Odrv4
    port map (
            O => \N__35865\,
            I => scaler_2_data_14
        );

    \I__7582\ : InMux
    port map (
            O => \N__35862\,
            I => \bfn_16_16_0_\
        );

    \I__7581\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35855\
        );

    \I__7580\ : CascadeMux
    port map (
            O => \N__35858\,
            I => \N__35852\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35849\
        );

    \I__7578\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35845\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__35849\,
            I => \N__35842\
        );

    \I__7576\ : InMux
    port map (
            O => \N__35848\,
            I => \N__35839\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__35845\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__35842\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__35839\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__35832\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\
        );

    \I__7571\ : InMux
    port map (
            O => \N__35829\,
            I => \N__35826\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__35826\,
            I => \N__35823\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__35823\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5\
        );

    \I__7568\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35815\
        );

    \I__7567\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35811\
        );

    \I__7566\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35808\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__35815\,
            I => \N__35805\
        );

    \I__7564\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35802\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__35811\,
            I => \N__35791\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__35808\,
            I => \N__35791\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__35805\,
            I => \N__35791\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__35802\,
            I => \N__35791\
        );

    \I__7559\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35788\
        );

    \I__7558\ : InMux
    port map (
            O => \N__35800\,
            I => \N__35785\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__35791\,
            I => \N__35772\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N__35772\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__35785\,
            I => \N__35772\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35769\
        );

    \I__7553\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35766\
        );

    \I__7552\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35761\
        );

    \I__7551\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35761\
        );

    \I__7550\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35756\
        );

    \I__7549\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35756\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__35772\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__35769\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__35766\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__35761\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__35756\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__7543\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35741\
        );

    \I__7542\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35738\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35735\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35723\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__35735\,
            I => \N__35723\
        );

    \I__7538\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35720\
        );

    \I__7537\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35717\
        );

    \I__7536\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35714\
        );

    \I__7535\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35711\
        );

    \I__7534\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35708\
        );

    \I__7533\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35703\
        );

    \I__7532\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35703\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__35723\,
            I => \N__35698\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35698\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35690\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__35714\,
            I => \N__35690\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__35711\,
            I => \N__35690\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__35708\,
            I => \N__35685\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__35703\,
            I => \N__35685\
        );

    \I__7524\ : Span4Mux_v
    port map (
            O => \N__35698\,
            I => \N__35680\
        );

    \I__7523\ : InMux
    port map (
            O => \N__35697\,
            I => \N__35677\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__35690\,
            I => \N__35672\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__35685\,
            I => \N__35672\
        );

    \I__7520\ : InMux
    port map (
            O => \N__35684\,
            I => \N__35667\
        );

    \I__7519\ : InMux
    port map (
            O => \N__35683\,
            I => \N__35667\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__35680\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__35677\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__35672\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__35667\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__35658\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14_cascade_\
        );

    \I__7513\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35652\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__35652\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__35649\,
            I => \N__35646\
        );

    \I__7510\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35642\
        );

    \I__7509\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35639\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35636\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__35639\,
            I => \N__35633\
        );

    \I__7506\ : Span4Mux_h
    port map (
            O => \N__35636\,
            I => \N__35630\
        );

    \I__7505\ : Odrv12
    port map (
            O => \N__35633\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__35630\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__7503\ : CascadeMux
    port map (
            O => \N__35625\,
            I => \N__35621\
        );

    \I__7502\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35616\
        );

    \I__7501\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35616\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__35616\,
            I => \N__35613\
        );

    \I__7499\ : Span4Mux_h
    port map (
            O => \N__35613\,
            I => \N__35610\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__35610\,
            I => \N__35607\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__35607\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__7496\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35601\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__35601\,
            I => \N__35597\
        );

    \I__7494\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35594\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__35597\,
            I => \N__35591\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__35594\,
            I => scaler_2_data_6
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__35591\,
            I => scaler_2_data_6
        );

    \I__7490\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35583\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__35583\,
            I => \N__35579\
        );

    \I__7488\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35576\
        );

    \I__7487\ : Span12Mux_s11_h
    port map (
            O => \N__35579\,
            I => \N__35573\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__35576\,
            I => scaler_2_data_7
        );

    \I__7485\ : Odrv12
    port map (
            O => \N__35573\,
            I => scaler_2_data_7
        );

    \I__7484\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35565\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__35565\,
            I => \N__35562\
        );

    \I__7482\ : Span12Mux_h
    port map (
            O => \N__35562\,
            I => \N__35559\
        );

    \I__7481\ : Odrv12
    port map (
            O => \N__35559\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__7480\ : InMux
    port map (
            O => \N__35556\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__7479\ : CascadeMux
    port map (
            O => \N__35553\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\
        );

    \I__7478\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35544\
        );

    \I__7477\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35537\
        );

    \I__7476\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35537\
        );

    \I__7475\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35537\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__35544\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__35537\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__7472\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35528\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__35531\,
            I => \N__35524\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__35528\,
            I => \N__35520\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35517\
        );

    \I__7468\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35512\
        );

    \I__7467\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35512\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__35520\,
            I => \N__35509\
        );

    \I__7465\ : LocalMux
    port map (
            O => \N__35517\,
            I => \N__35506\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__35512\,
            I => \N__35503\
        );

    \I__7463\ : Span4Mux_v
    port map (
            O => \N__35509\,
            I => \N__35500\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__7461\ : Odrv4
    port map (
            O => \N__35503\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__35500\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__7459\ : Odrv4
    port map (
            O => \N__35497\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__7458\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35487\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__35487\,
            I => \N__35484\
        );

    \I__7456\ : Span4Mux_h
    port map (
            O => \N__35484\,
            I => \N__35481\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__35481\,
            I => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\
        );

    \I__7454\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35474\
        );

    \I__7453\ : CascadeMux
    port map (
            O => \N__35477\,
            I => \N__35470\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__35474\,
            I => \N__35467\
        );

    \I__7451\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35464\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35461\
        );

    \I__7449\ : Span4Mux_h
    port map (
            O => \N__35467\,
            I => \N__35456\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__35464\,
            I => \N__35456\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35461\,
            I => throttle_command_3
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__35456\,
            I => throttle_command_3
        );

    \I__7445\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35447\
        );

    \I__7444\ : CascadeMux
    port map (
            O => \N__35450\,
            I => \N__35443\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35440\
        );

    \I__7442\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35435\
        );

    \I__7441\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35435\
        );

    \I__7440\ : Odrv4
    port map (
            O => \N__35440\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__35435\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__7438\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35426\
        );

    \I__7437\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35423\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35420\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35417\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__35420\,
            I => \N__35412\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__35417\,
            I => \N__35412\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__35412\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__7431\ : CascadeMux
    port map (
            O => \N__35409\,
            I => \N__35405\
        );

    \I__7430\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35402\
        );

    \I__7429\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35399\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__35402\,
            I => \N__35396\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__35399\,
            I => \N__35393\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__35396\,
            I => \N__35388\
        );

    \I__7425\ : Span4Mux_v
    port map (
            O => \N__35393\,
            I => \N__35388\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__35388\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__35385\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__35382\,
            I => \N__35379\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35375\
        );

    \I__7420\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35371\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__35375\,
            I => \N__35368\
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__35374\,
            I => \N__35365\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35371\,
            I => \N__35360\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__35368\,
            I => \N__35360\
        );

    \I__7415\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35357\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__35360\,
            I => \N__35354\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__35357\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__35354\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__35349\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\
        );

    \I__7410\ : InMux
    port map (
            O => \N__35346\,
            I => \N__35343\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__35343\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4\
        );

    \I__7408\ : CascadeMux
    port map (
            O => \N__35340\,
            I => \N__35335\
        );

    \I__7407\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35330\
        );

    \I__7406\ : InMux
    port map (
            O => \N__35338\,
            I => \N__35330\
        );

    \I__7405\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35327\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__35330\,
            I => \N__35322\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__35327\,
            I => \N__35322\
        );

    \I__7402\ : Odrv4
    port map (
            O => \N__35322\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35316\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__35316\,
            I => \N__35313\
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__35313\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35302\
        );

    \I__7397\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35302\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35299\
        );

    \I__7395\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35296\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__35302\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__35299\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__35296\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35282\
        );

    \I__7390\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35279\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35276\
        );

    \I__7388\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35273\
        );

    \I__7387\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35270\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35256\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35256\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35256\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35256\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35256\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35251\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35251\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35245\
        );

    \I__7378\ : Span4Mux_v
    port map (
            O => \N__35256\,
            I => \N__35240\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35240\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35233\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35249\,
            I => \N__35233\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35233\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35245\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__35240\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__35233\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__7370\ : CascadeMux
    port map (
            O => \N__35226\,
            I => \N__35223\
        );

    \I__7369\ : InMux
    port map (
            O => \N__35223\,
            I => \N__35219\
        );

    \I__7368\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35215\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__35219\,
            I => \N__35212\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35209\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35206\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__35212\,
            I => \N__35203\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__35209\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__7362\ : Odrv12
    port map (
            O => \N__35206\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__35203\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__7360\ : CascadeMux
    port map (
            O => \N__35196\,
            I => \N__35193\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35189\
        );

    \I__7358\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__35189\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__35186\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__7355\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35177\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35174\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35177\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35174\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__7351\ : CascadeMux
    port map (
            O => \N__35169\,
            I => \N__35165\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35160\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35160\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__35160\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__7347\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35153\
        );

    \I__7346\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35150\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__35153\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__35150\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__35145\,
            I => \N__35142\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__35139\,
            I => \reset_module_System.reset6_11\
        );

    \I__7340\ : CascadeMux
    port map (
            O => \N__35136\,
            I => \ppm_encoder_1.N_297_cascade_\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__35133\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_\
        );

    \I__7338\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35125\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35122\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35119\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__35125\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35122\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__35119\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35112\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35109\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35102\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35099\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__35102\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__35099\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35094\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35091\,
            I => \bfn_16_9_0_\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35084\
        );

    \I__7323\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35081\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__35084\,
            I => \N__35078\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__35081\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__35078\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35073\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35070\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__7317\ : CascadeMux
    port map (
            O => \N__35067\,
            I => \N__35063\
        );

    \I__7316\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35057\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__35060\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__35057\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__7312\ : InMux
    port map (
            O => \N__35052\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__7311\ : InMux
    port map (
            O => \N__35049\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__35046\,
            I => \N__35043\
        );

    \I__7309\ : InMux
    port map (
            O => \N__35043\,
            I => \N__35037\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35037\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__35037\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35030\
        );

    \I__7305\ : InMux
    port map (
            O => \N__35033\,
            I => \N__35027\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35030\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__35027\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__7302\ : InMux
    port map (
            O => \N__35022\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35019\,
            I => \N__35015\
        );

    \I__7300\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35012\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__35015\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__35012\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35007\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35004\,
            I => \N__35000\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35003\,
            I => \N__34997\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35000\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__34997\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__7292\ : InMux
    port map (
            O => \N__34992\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__7291\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34985\
        );

    \I__7290\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34982\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__34985\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__34982\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__7287\ : InMux
    port map (
            O => \N__34977\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__34974\,
            I => \N__34971\
        );

    \I__7285\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34967\
        );

    \I__7284\ : InMux
    port map (
            O => \N__34970\,
            I => \N__34964\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34961\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__34964\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__34961\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__7280\ : InMux
    port map (
            O => \N__34956\,
            I => \bfn_16_8_0_\
        );

    \I__7279\ : InMux
    port map (
            O => \N__34953\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__7278\ : InMux
    port map (
            O => \N__34950\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__7277\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34943\
        );

    \I__7276\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34940\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__34943\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__34940\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__7273\ : InMux
    port map (
            O => \N__34935\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__7272\ : InMux
    port map (
            O => \N__34932\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__34929\,
            I => \N__34925\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__34928\,
            I => \N__34922\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34918\
        );

    \I__7268\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34915\
        );

    \I__7267\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34912\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34909\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__34915\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__34912\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__34909\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__7262\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__34896\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__7259\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34889\
        );

    \I__7258\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34886\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__34889\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__34886\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__34878\,
            I => \N__34875\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__34875\,
            I => \N__34872\
        );

    \I__7252\ : Sp12to4
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__7251\ : Odrv12
    port map (
            O => \N__34869\,
            I => \pid_alt.O_0_5\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__7249\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__34857\,
            I => \pid_alt.error_i_regZ0Z_1\
        );

    \I__7246\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34850\
        );

    \I__7245\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34846\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__34850\,
            I => \N__34843\
        );

    \I__7243\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34840\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__34846\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7241\ : Odrv12
    port map (
            O => \N__34843\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__34840\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__34833\,
            I => \N__34828\
        );

    \I__7238\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34825\
        );

    \I__7237\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34822\
        );

    \I__7236\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34819\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__34825\,
            I => \N__34815\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__34822\,
            I => \N__34812\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__34819\,
            I => \N__34809\
        );

    \I__7232\ : InMux
    port map (
            O => \N__34818\,
            I => \N__34806\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__34815\,
            I => \N__34803\
        );

    \I__7230\ : Sp12to4
    port map (
            O => \N__34812\,
            I => \N__34798\
        );

    \I__7229\ : Span12Mux_s8_v
    port map (
            O => \N__34809\,
            I => \N__34798\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__34806\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__34803\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__7226\ : Odrv12
    port map (
            O => \N__34798\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__7225\ : InMux
    port map (
            O => \N__34791\,
            I => \N__34787\
        );

    \I__7224\ : InMux
    port map (
            O => \N__34790\,
            I => \N__34784\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__34787\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__34784\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7221\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__34776\,
            I => \reset_module_System.count_1_2\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34773\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__7218\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34766\
        );

    \I__7217\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34763\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__34766\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__34763\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__7214\ : InMux
    port map (
            O => \N__34758\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__7213\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34751\
        );

    \I__7212\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34748\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__34751\,
            I => \N__34745\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__34748\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__34745\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__7208\ : InMux
    port map (
            O => \N__34740\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__7207\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34732\
        );

    \I__7206\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34727\
        );

    \I__7205\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34727\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__34732\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__34727\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__7202\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__34719\,
            I => \ppm_encoder_1.N_145_17\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__34716\,
            I => \ppm_encoder_1.N_145_17_cascade_\
        );

    \I__7199\ : InMux
    port map (
            O => \N__34713\,
            I => \N__34704\
        );

    \I__7198\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34704\
        );

    \I__7197\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34704\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__34704\,
            I => \ppm_encoder_1.N_238\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__34701\,
            I => \N__34698\
        );

    \I__7194\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34695\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__34695\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__7192\ : InMux
    port map (
            O => \N__34692\,
            I => \N__34689\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__34689\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10\
        );

    \I__7190\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34683\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10\
        );

    \I__7188\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34676\
        );

    \I__7187\ : CascadeMux
    port map (
            O => \N__34679\,
            I => \N__34672\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__34676\,
            I => \N__34668\
        );

    \I__7185\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34665\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34660\
        );

    \I__7183\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34660\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__34668\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__34665\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__34660\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__7179\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34650\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__34650\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__34647\,
            I => \N__34644\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34641\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__34641\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\
        );

    \I__7174\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34635\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__34635\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__34632\,
            I => \N__34627\
        );

    \I__7171\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34624\
        );

    \I__7170\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34619\
        );

    \I__7169\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34619\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__34624\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__34619\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__7166\ : CascadeMux
    port map (
            O => \N__34614\,
            I => \ppm_encoder_1.N_303_cascade_\
        );

    \I__7165\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34608\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__34608\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__34605\,
            I => \N__34602\
        );

    \I__7162\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34597\
        );

    \I__7161\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34594\
        );

    \I__7160\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34591\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__34597\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__34594\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__34591\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__34584\,
            I => \ppm_encoder_1.N_319_cascade_\
        );

    \I__7155\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34578\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__34578\,
            I => \N__34574\
        );

    \I__7153\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34571\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__34574\,
            I => \N__34567\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__34571\,
            I => \N__34564\
        );

    \I__7150\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34561\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__34567\,
            I => \N__34558\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__34564\,
            I => \N__34555\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__34561\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__34558\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__34555\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7144\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__34545\,
            I => \ppm_encoder_1.N_302\
        );

    \I__7142\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34539\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__7140\ : Span4Mux_v
    port map (
            O => \N__34536\,
            I => \N__34533\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34530\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__34530\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__7137\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__34524\,
            I => \N__34521\
        );

    \I__7135\ : Span4Mux_h
    port map (
            O => \N__34521\,
            I => \N__34517\
        );

    \I__7134\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34514\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__34517\,
            I => scaler_4_data_8
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__34514\,
            I => scaler_4_data_8
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__34509\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\
        );

    \I__7130\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__34503\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13\
        );

    \I__7128\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34496\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34493\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34490\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__34493\,
            I => \N__34487\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__34490\,
            I => \N__34484\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__34487\,
            I => \N__34481\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__34484\,
            I => scaler_3_data_13
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__34481\,
            I => scaler_3_data_13
        );

    \I__7120\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34473\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34470\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__34470\,
            I => \N__34467\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__34467\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__7116\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34461\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__34461\,
            I => \N__34457\
        );

    \I__7114\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34454\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__34457\,
            I => \N__34449\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34449\
        );

    \I__7111\ : Span4Mux_h
    port map (
            O => \N__34449\,
            I => \N__34446\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__34443\,
            I => throttle_command_13
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__34440\,
            I => \N__34437\
        );

    \I__7107\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34434\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34431\
        );

    \I__7105\ : Span4Mux_h
    port map (
            O => \N__34431\,
            I => \N__34428\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__34428\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__34425\,
            I => \N__34420\
        );

    \I__7102\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34417\
        );

    \I__7101\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34412\
        );

    \I__7100\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34412\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__34417\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__34412\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__34407\,
            I => \N__34402\
        );

    \I__7096\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34399\
        );

    \I__7095\ : InMux
    port map (
            O => \N__34405\,
            I => \N__34394\
        );

    \I__7094\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34394\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__34399\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__34394\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__7091\ : CascadeMux
    port map (
            O => \N__34389\,
            I => \ppm_encoder_1.N_305_cascade_\
        );

    \I__7090\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34381\
        );

    \I__7089\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34376\
        );

    \I__7088\ : InMux
    port map (
            O => \N__34384\,
            I => \N__34376\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__34381\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__34376\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__34371\,
            I => \ppm_encoder_1.N_298_cascade_\
        );

    \I__7084\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34359\
        );

    \I__7083\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34359\
        );

    \I__7082\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34359\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__34359\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__7080\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34352\
        );

    \I__7079\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34349\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34346\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34343\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__34346\,
            I => \N__34340\
        );

    \I__7075\ : Odrv12
    port map (
            O => \N__34343\,
            I => scaler_3_data_6
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__34340\,
            I => scaler_3_data_6
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__34335\,
            I => \N__34330\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34323\
        );

    \I__7071\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34323\
        );

    \I__7070\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34323\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34323\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__7068\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34314\
        );

    \I__7066\ : Span4Mux_h
    port map (
            O => \N__34314\,
            I => \N__34311\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__34311\,
            I => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34304\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__34307\,
            I => \N__34301\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34304\,
            I => \N__34298\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34295\
        );

    \I__7060\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34292\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__34295\,
            I => \N__34289\
        );

    \I__7058\ : Span4Mux_h
    port map (
            O => \N__34292\,
            I => \N__34286\
        );

    \I__7057\ : Span4Mux_h
    port map (
            O => \N__34289\,
            I => \N__34283\
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__34286\,
            I => throttle_command_6
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__34283\,
            I => throttle_command_6
        );

    \I__7054\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34271\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34271\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34268\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__34271\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34268\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__7049\ : CascadeMux
    port map (
            O => \N__34263\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8_cascade_\
        );

    \I__7048\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34257\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__7046\ : Odrv12
    port map (
            O => \N__34254\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8\
        );

    \I__7045\ : CascadeMux
    port map (
            O => \N__34251\,
            I => \N__34247\
        );

    \I__7044\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34242\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34242\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__34242\,
            I => \N__34238\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34235\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__34238\,
            I => \N__34232\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__34235\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7038\ : Odrv4
    port map (
            O => \N__34232\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7037\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34224\,
            I => \N__34220\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34217\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__34220\,
            I => \N__34214\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__34217\,
            I => \N__34211\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__34214\,
            I => \N__34208\
        );

    \I__7031\ : Span4Mux_h
    port map (
            O => \N__34211\,
            I => \N__34205\
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__34208\,
            I => throttle_command_8
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__34205\,
            I => throttle_command_8
        );

    \I__7028\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34197\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__7026\ : Span4Mux_h
    port map (
            O => \N__34194\,
            I => \N__34191\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__34191\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34180\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34175\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34175\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__34180\,
            I => \N__34172\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34175\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__34172\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__7017\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34163\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__34166\,
            I => \N__34160\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34163\,
            I => \N__34157\
        );

    \I__7014\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34154\
        );

    \I__7013\ : Span4Mux_v
    port map (
            O => \N__34157\,
            I => \N__34149\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__34154\,
            I => \N__34149\
        );

    \I__7011\ : Odrv4
    port map (
            O => \N__34149\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__34146\,
            I => \ppm_encoder_1.N_296_cascade_\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34140\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34136\
        );

    \I__7007\ : InMux
    port map (
            O => \N__34139\,
            I => \N__34133\
        );

    \I__7006\ : Span4Mux_v
    port map (
            O => \N__34136\,
            I => \N__34128\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34128\
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__34128\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__34125\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__34122\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6_cascade_\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34116\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__34116\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__34113\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__34110\,
            I => \ppm_encoder_1.N_227_cascade_\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__34107\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34101\,
            I => \N__34095\
        );

    \I__6994\ : InMux
    port map (
            O => \N__34100\,
            I => \N__34095\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__34095\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__34092\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__6991\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34086\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__34086\,
            I => \N__34083\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__34083\,
            I => \N__34080\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__34080\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34077\,
            I => \N__34074\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__34071\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34068\,
            I => \N__34065\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__34065\,
            I => \N__34061\
        );

    \I__6982\ : CascadeMux
    port map (
            O => \N__34064\,
            I => \N__34057\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__34061\,
            I => \N__34054\
        );

    \I__6980\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34049\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34057\,
            I => \N__34049\
        );

    \I__6978\ : Odrv4
    port map (
            O => \N__34054\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34049\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__6976\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34041\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__34037\
        );

    \I__6974\ : CascadeMux
    port map (
            O => \N__34040\,
            I => \N__34033\
        );

    \I__6973\ : Span4Mux_v
    port map (
            O => \N__34037\,
            I => \N__34030\
        );

    \I__6972\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34025\
        );

    \I__6971\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34025\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__34030\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__34025\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__6968\ : InMux
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__6966\ : Span4Mux_v
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__34011\,
            I => \ppm_encoder_1.N_304\
        );

    \I__6964\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__34005\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__6962\ : CascadeMux
    port map (
            O => \N__34002\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\
        );

    \I__6961\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33994\
        );

    \I__6960\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33991\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33988\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__33994\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__33991\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__33988\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__6955\ : CascadeMux
    port map (
            O => \N__33981\,
            I => \N__33976\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__33980\,
            I => \N__33973\
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__33979\,
            I => \N__33970\
        );

    \I__6952\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33967\
        );

    \I__6951\ : InMux
    port map (
            O => \N__33973\,
            I => \N__33962\
        );

    \I__6950\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33962\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__33967\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__33962\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__6947\ : CascadeMux
    port map (
            O => \N__33957\,
            I => \N__33951\
        );

    \I__6946\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33948\
        );

    \I__6945\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33945\
        );

    \I__6944\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33940\
        );

    \I__6943\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33940\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__33948\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__33945\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__33940\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__33933\,
            I => \uart_drone.timer_Count_RNO_0_0_1_cascade_\
        );

    \I__6938\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33926\
        );

    \I__6937\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33923\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__33926\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__33923\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__6934\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33908\
        );

    \I__6933\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33908\
        );

    \I__6932\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33905\
        );

    \I__6931\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33902\
        );

    \I__6930\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33899\
        );

    \I__6929\ : InMux
    port map (
            O => \N__33913\,
            I => \N__33896\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__33908\,
            I => \uart_drone.N_143\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__33905\,
            I => \uart_drone.N_143\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33902\,
            I => \uart_drone.N_143\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__33899\,
            I => \uart_drone.N_143\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__33896\,
            I => \uart_drone.N_143\
        );

    \I__6923\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33881\
        );

    \I__6922\ : CascadeMux
    port map (
            O => \N__33884\,
            I => \N__33878\
        );

    \I__6921\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__6920\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33872\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33864\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__33872\,
            I => \N__33864\
        );

    \I__6917\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33859\
        );

    \I__6916\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33859\
        );

    \I__6915\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33856\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__33864\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__33859\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__33856\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__6910\ : InMux
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__33843\,
            I => \N__33837\
        );

    \I__6908\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33834\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__33841\,
            I => \N__33831\
        );

    \I__6906\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33828\
        );

    \I__6905\ : Span4Mux_v
    port map (
            O => \N__33837\,
            I => \N__33823\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__33834\,
            I => \N__33823\
        );

    \I__6903\ : InMux
    port map (
            O => \N__33831\,
            I => \N__33820\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__33828\,
            I => \N__33817\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__33823\,
            I => \N__33814\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__33820\,
            I => \N__33811\
        );

    \I__6899\ : Span4Mux_h
    port map (
            O => \N__33817\,
            I => \N__33808\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__33814\,
            I => \reset_module_System.reset6_15\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__33811\,
            I => \reset_module_System.reset6_15\
        );

    \I__6896\ : Odrv4
    port map (
            O => \N__33808\,
            I => \reset_module_System.reset6_15\
        );

    \I__6895\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33798\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__33795\,
            I => \reset_module_System.reset6_17\
        );

    \I__6892\ : InMux
    port map (
            O => \N__33792\,
            I => \N__33788\
        );

    \I__6891\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33783\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33780\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33777\
        );

    \I__6888\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33774\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__33783\,
            I => \N__33771\
        );

    \I__6886\ : Span4Mux_h
    port map (
            O => \N__33780\,
            I => \N__33768\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33765\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33760\
        );

    \I__6883\ : Span12Mux_s8_v
    port map (
            O => \N__33771\,
            I => \N__33760\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__33768\,
            I => \reset_module_System.reset6_19\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__33765\,
            I => \reset_module_System.reset6_19\
        );

    \I__6880\ : Odrv12
    port map (
            O => \N__33760\,
            I => \reset_module_System.reset6_19\
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__33753\,
            I => \N__33747\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__33752\,
            I => \N__33744\
        );

    \I__6877\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33741\
        );

    \I__6876\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33738\
        );

    \I__6875\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33735\
        );

    \I__6874\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33732\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__33741\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__33738\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__33735\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__33732\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__33723\,
            I => \uart_drone.N_145_cascade_\
        );

    \I__6868\ : SRMux
    port map (
            O => \N__33720\,
            I => \N__33715\
        );

    \I__6867\ : SRMux
    port map (
            O => \N__33719\,
            I => \N__33712\
        );

    \I__6866\ : SRMux
    port map (
            O => \N__33718\,
            I => \N__33709\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__33715\,
            I => \N__33704\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__33712\,
            I => \N__33704\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33700\
        );

    \I__6862\ : Span4Mux_v
    port map (
            O => \N__33704\,
            I => \N__33697\
        );

    \I__6861\ : SRMux
    port map (
            O => \N__33703\,
            I => \N__33694\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__33700\,
            I => \N__33690\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__33697\,
            I => \N__33687\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33684\
        );

    \I__6857\ : SRMux
    port map (
            O => \N__33693\,
            I => \N__33681\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__33690\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__33687\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__6854\ : Odrv12
    port map (
            O => \N__33684\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__33681\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__6852\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33669\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__33666\,
            I => \N__33662\
        );

    \I__6849\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33659\
        );

    \I__6848\ : Odrv4
    port map (
            O => \N__33662\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__33659\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__6846\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33650\
        );

    \I__6845\ : InMux
    port map (
            O => \N__33653\,
            I => \N__33647\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33644\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__33647\,
            I => \N__33641\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__33644\,
            I => \N__33638\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__33641\,
            I => \N__33635\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__33638\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__33635\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__6838\ : CEMux
    port map (
            O => \N__33630\,
            I => \N__33531\
        );

    \I__6837\ : CEMux
    port map (
            O => \N__33629\,
            I => \N__33531\
        );

    \I__6836\ : CEMux
    port map (
            O => \N__33628\,
            I => \N__33531\
        );

    \I__6835\ : CEMux
    port map (
            O => \N__33627\,
            I => \N__33531\
        );

    \I__6834\ : CEMux
    port map (
            O => \N__33626\,
            I => \N__33531\
        );

    \I__6833\ : CEMux
    port map (
            O => \N__33625\,
            I => \N__33531\
        );

    \I__6832\ : CEMux
    port map (
            O => \N__33624\,
            I => \N__33531\
        );

    \I__6831\ : CEMux
    port map (
            O => \N__33623\,
            I => \N__33531\
        );

    \I__6830\ : CEMux
    port map (
            O => \N__33622\,
            I => \N__33531\
        );

    \I__6829\ : CEMux
    port map (
            O => \N__33621\,
            I => \N__33531\
        );

    \I__6828\ : CEMux
    port map (
            O => \N__33620\,
            I => \N__33531\
        );

    \I__6827\ : CEMux
    port map (
            O => \N__33619\,
            I => \N__33531\
        );

    \I__6826\ : CEMux
    port map (
            O => \N__33618\,
            I => \N__33531\
        );

    \I__6825\ : CEMux
    port map (
            O => \N__33617\,
            I => \N__33531\
        );

    \I__6824\ : CEMux
    port map (
            O => \N__33616\,
            I => \N__33531\
        );

    \I__6823\ : CEMux
    port map (
            O => \N__33615\,
            I => \N__33531\
        );

    \I__6822\ : CEMux
    port map (
            O => \N__33614\,
            I => \N__33531\
        );

    \I__6821\ : CEMux
    port map (
            O => \N__33613\,
            I => \N__33531\
        );

    \I__6820\ : CEMux
    port map (
            O => \N__33612\,
            I => \N__33531\
        );

    \I__6819\ : CEMux
    port map (
            O => \N__33611\,
            I => \N__33531\
        );

    \I__6818\ : CEMux
    port map (
            O => \N__33610\,
            I => \N__33531\
        );

    \I__6817\ : CEMux
    port map (
            O => \N__33609\,
            I => \N__33531\
        );

    \I__6816\ : CEMux
    port map (
            O => \N__33608\,
            I => \N__33531\
        );

    \I__6815\ : CEMux
    port map (
            O => \N__33607\,
            I => \N__33531\
        );

    \I__6814\ : CEMux
    port map (
            O => \N__33606\,
            I => \N__33531\
        );

    \I__6813\ : CEMux
    port map (
            O => \N__33605\,
            I => \N__33531\
        );

    \I__6812\ : CEMux
    port map (
            O => \N__33604\,
            I => \N__33531\
        );

    \I__6811\ : CEMux
    port map (
            O => \N__33603\,
            I => \N__33531\
        );

    \I__6810\ : CEMux
    port map (
            O => \N__33602\,
            I => \N__33531\
        );

    \I__6809\ : CEMux
    port map (
            O => \N__33601\,
            I => \N__33531\
        );

    \I__6808\ : CEMux
    port map (
            O => \N__33600\,
            I => \N__33531\
        );

    \I__6807\ : CEMux
    port map (
            O => \N__33599\,
            I => \N__33531\
        );

    \I__6806\ : CEMux
    port map (
            O => \N__33598\,
            I => \N__33531\
        );

    \I__6805\ : GlobalMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6804\ : gio2CtrlBuf
    port map (
            O => \N__33528\,
            I => \pid_alt.state_0_g_0\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6802\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__33519\,
            I => \N__33516\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__33513\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__6798\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33505\
        );

    \I__6797\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33502\
        );

    \I__6796\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33499\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33496\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__33502\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__33499\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__33496\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6791\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33486\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__33486\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33483\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__6788\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__6786\ : Span4Mux_v
    port map (
            O => \N__33474\,
            I => \N__33471\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__33471\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__6784\ : InMux
    port map (
            O => \N__33468\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__6783\ : InMux
    port map (
            O => \N__33465\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__6782\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33459\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__33459\,
            I => \N__33456\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__33456\,
            I => \N__33453\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__33453\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__6778\ : CascadeMux
    port map (
            O => \N__33450\,
            I => \reset_module_System.reset6_13_cascade_\
        );

    \I__6777\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__33444\,
            I => \reset_module_System.reset6_3\
        );

    \I__6775\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33436\
        );

    \I__6774\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33432\
        );

    \I__6773\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33429\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33426\
        );

    \I__6771\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33423\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__33432\,
            I => \N__33420\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33417\
        );

    \I__6768\ : Span4Mux_v
    port map (
            O => \N__33426\,
            I => \N__33414\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33423\,
            I => \N__33410\
        );

    \I__6766\ : Span4Mux_v
    port map (
            O => \N__33420\,
            I => \N__33406\
        );

    \I__6765\ : Span4Mux_v
    port map (
            O => \N__33417\,
            I => \N__33401\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__33414\,
            I => \N__33398\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33395\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__33410\,
            I => \N__33390\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33386\
        );

    \I__6760\ : Span4Mux_h
    port map (
            O => \N__33406\,
            I => \N__33383\
        );

    \I__6759\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33380\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__33404\,
            I => \N__33377\
        );

    \I__6757\ : Span4Mux_h
    port map (
            O => \N__33401\,
            I => \N__33374\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__33398\,
            I => \N__33369\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__33395\,
            I => \N__33369\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33366\
        );

    \I__6753\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33363\
        );

    \I__6752\ : Span4Mux_v
    port map (
            O => \N__33390\,
            I => \N__33359\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33356\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__33386\,
            I => \N__33349\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__33383\,
            I => \N__33349\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__33380\,
            I => \N__33349\
        );

    \I__6747\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33346\
        );

    \I__6746\ : Span4Mux_h
    port map (
            O => \N__33374\,
            I => \N__33336\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__33369\,
            I => \N__33336\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33336\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__33363\,
            I => \N__33336\
        );

    \I__6742\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33333\
        );

    \I__6741\ : Sp12to4
    port map (
            O => \N__33359\,
            I => \N__33330\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33325\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__33349\,
            I => \N__33325\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33322\
        );

    \I__6737\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33319\
        );

    \I__6736\ : Sp12to4
    port map (
            O => \N__33336\,
            I => \N__33312\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33312\
        );

    \I__6734\ : Span12Mux_h
    port map (
            O => \N__33330\,
            I => \N__33312\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__33325\,
            I => \N__33307\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__33322\,
            I => \N__33307\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__33319\,
            I => uart_pc_data_6
        );

    \I__6730\ : Odrv12
    port map (
            O => \N__33312\,
            I => uart_pc_data_6
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__33307\,
            I => uart_pc_data_6
        );

    \I__6728\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6726\ : Span4Mux_s2_h
    port map (
            O => \N__33294\,
            I => \N__33291\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__33288\,
            I => \N__33285\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__33285\,
            I => alt_ki_6
        );

    \I__6722\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__33276\,
            I => \N__33271\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33266\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33266\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__33271\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__33266\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33257\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33254\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__33254\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33251\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__33246\,
            I => \N__33241\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__33245\,
            I => \N__33237\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__33244\,
            I => \N__33232\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33241\,
            I => \N__33224\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33224\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33219\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33219\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33210\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33210\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33210\
        );

    \I__6700\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33210\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33205\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33201\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33196\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__33210\,
            I => \N__33196\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33191\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33191\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__33205\,
            I => \N__33188\
        );

    \I__6692\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33185\
        );

    \I__6691\ : Span4Mux_v
    port map (
            O => \N__33201\,
            I => \N__33182\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__33196\,
            I => \N__33178\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33175\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__33188\,
            I => \N__33167\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__33185\,
            I => \N__33167\
        );

    \I__6686\ : Span4Mux_h
    port map (
            O => \N__33182\,
            I => \N__33160\
        );

    \I__6685\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33157\
        );

    \I__6684\ : Span4Mux_v
    port map (
            O => \N__33178\,
            I => \N__33152\
        );

    \I__6683\ : Span4Mux_v
    port map (
            O => \N__33175\,
            I => \N__33152\
        );

    \I__6682\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33147\
        );

    \I__6681\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33147\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__33172\,
            I => \N__33143\
        );

    \I__6679\ : Span4Mux_h
    port map (
            O => \N__33167\,
            I => \N__33140\
        );

    \I__6678\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33131\
        );

    \I__6677\ : InMux
    port map (
            O => \N__33165\,
            I => \N__33131\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33131\
        );

    \I__6675\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33131\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__33160\,
            I => \N__33126\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__33157\,
            I => \N__33126\
        );

    \I__6672\ : Span4Mux_h
    port map (
            O => \N__33152\,
            I => \N__33121\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33147\,
            I => \N__33121\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33116\
        );

    \I__6669\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33116\
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__33140\,
            I => \pid_alt.N_96_i\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__33131\,
            I => \pid_alt.N_96_i\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__33126\,
            I => \pid_alt.N_96_i\
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__33121\,
            I => \pid_alt.N_96_i\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__33116\,
            I => \pid_alt.N_96_i\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33094\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33091\
        );

    \I__6659\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33088\
        );

    \I__6658\ : Span4Mux_h
    port map (
            O => \N__33094\,
            I => \N__33081\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__33091\,
            I => \N__33081\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__33088\,
            I => \N__33081\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__33081\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__6654\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33071\
        );

    \I__6653\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33071\
        );

    \I__6652\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33064\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__33071\,
            I => \N__33061\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33058\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33069\,
            I => \N__33051\
        );

    \I__6648\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33051\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33051\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__33064\,
            I => \N__33044\
        );

    \I__6645\ : Span4Mux_v
    port map (
            O => \N__33061\,
            I => \N__33044\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__33058\,
            I => \N__33039\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33039\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33034\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33049\,
            I => \N__33034\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__33044\,
            I => \pid_alt.N_128\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__33039\,
            I => \pid_alt.N_128\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__33034\,
            I => \pid_alt.N_128\
        );

    \I__6637\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33023\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33020\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__33023\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__33020\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__6633\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__33008\
        );

    \I__6631\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33005\
        );

    \I__6630\ : Span4Mux_h
    port map (
            O => \N__33008\,
            I => \N__33002\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__33005\,
            I => \N__32999\
        );

    \I__6628\ : Span4Mux_v
    port map (
            O => \N__33002\,
            I => \N__32996\
        );

    \I__6627\ : Span4Mux_v
    port map (
            O => \N__32999\,
            I => \N__32993\
        );

    \I__6626\ : Odrv4
    port map (
            O => \N__32996\,
            I => scaler_3_data_10
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__32993\,
            I => scaler_3_data_10
        );

    \I__6624\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32985\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__32985\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__32982\,
            I => \N__32977\
        );

    \I__6621\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32970\
        );

    \I__6620\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32970\
        );

    \I__6619\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32970\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__32970\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__6617\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32964\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__6615\ : Span4Mux_h
    port map (
            O => \N__32961\,
            I => \N__32957\
        );

    \I__6614\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32954\
        );

    \I__6613\ : Odrv4
    port map (
            O => \N__32957\,
            I => scaler_4_data_10
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__32954\,
            I => scaler_4_data_10
        );

    \I__6611\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__32946\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__6609\ : CascadeMux
    port map (
            O => \N__32943\,
            I => \N__32939\
        );

    \I__6608\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32935\
        );

    \I__6607\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32932\
        );

    \I__6606\ : IoInMux
    port map (
            O => \N__32938\,
            I => \N__32929\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32923\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32923\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__32929\,
            I => \N__32920\
        );

    \I__6602\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32917\
        );

    \I__6601\ : Span4Mux_h
    port map (
            O => \N__32923\,
            I => \N__32914\
        );

    \I__6600\ : IoSpan4Mux
    port map (
            O => \N__32920\,
            I => \N__32911\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32908\
        );

    \I__6598\ : Span4Mux_v
    port map (
            O => \N__32914\,
            I => \N__32905\
        );

    \I__6597\ : Span4Mux_s3_v
    port map (
            O => \N__32911\,
            I => \N__32902\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__32908\,
            I => \N__32899\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__32905\,
            I => \N__32896\
        );

    \I__6594\ : Span4Mux_v
    port map (
            O => \N__32902\,
            I => \N__32893\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__32899\,
            I => reset_system
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__32896\,
            I => reset_system
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__32893\,
            I => reset_system
        );

    \I__6590\ : IoInMux
    port map (
            O => \N__32886\,
            I => \N__32883\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__6588\ : Span4Mux_s3_v
    port map (
            O => \N__32880\,
            I => \N__32877\
        );

    \I__6587\ : Span4Mux_v
    port map (
            O => \N__32877\,
            I => \N__32874\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__32874\,
            I => \N__32871\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__32871\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__6584\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32865\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32862\
        );

    \I__6582\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__32859\,
            I => \ppm_encoder_1.N_145\
        );

    \I__6580\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32849\
        );

    \I__6578\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32846\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__32849\,
            I => \N__32839\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__32846\,
            I => \N__32839\
        );

    \I__6575\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32836\
        );

    \I__6574\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32833\
        );

    \I__6573\ : Odrv4
    port map (
            O => \N__32839\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__32836\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__32833\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6570\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32823\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32818\
        );

    \I__6568\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32815\
        );

    \I__6567\ : InMux
    port map (
            O => \N__32821\,
            I => \N__32812\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__32818\,
            I => \N__32805\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32805\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32805\
        );

    \I__6563\ : Span4Mux_h
    port map (
            O => \N__32805\,
            I => \N__32802\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__32802\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__6561\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32796\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__32796\,
            I => \N__32792\
        );

    \I__6559\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32789\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__32792\,
            I => \pid_alt.N_238\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__32789\,
            I => \pid_alt.N_238\
        );

    \I__6556\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32778\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__32778\,
            I => \pid_alt.error_i_acummZ0Z_13\
        );

    \I__6553\ : CEMux
    port map (
            O => \N__32775\,
            I => \N__32772\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32768\
        );

    \I__6551\ : CEMux
    port map (
            O => \N__32771\,
            I => \N__32765\
        );

    \I__6550\ : Span4Mux_h
    port map (
            O => \N__32768\,
            I => \N__32762\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32759\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__32762\,
            I => \pid_alt.N_96_i_0\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__32759\,
            I => \pid_alt.N_96_i_0\
        );

    \I__6546\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__32751\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__6544\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32745\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32745\,
            I => \N__32742\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__32742\,
            I => \N__32738\
        );

    \I__6541\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32735\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__32738\,
            I => scaler_4_data_11
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__32735\,
            I => scaler_4_data_11
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__32730\,
            I => \N__32727\
        );

    \I__6537\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32724\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32720\
        );

    \I__6535\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__6534\ : Span4Mux_h
    port map (
            O => \N__32720\,
            I => \N__32712\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32712\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__32712\,
            I => \N__32709\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__32709\,
            I => throttle_command_11
        );

    \I__6530\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32703\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32700\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__32700\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__6527\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32693\
        );

    \I__6526\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32690\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__32693\,
            I => \N__32687\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__32690\,
            I => \N__32684\
        );

    \I__6523\ : Span4Mux_v
    port map (
            O => \N__32687\,
            I => \N__32681\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__32684\,
            I => \N__32678\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__32681\,
            I => scaler_3_data_11
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__32678\,
            I => scaler_3_data_11
        );

    \I__6519\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__6517\ : Span4Mux_h
    port map (
            O => \N__32667\,
            I => \N__32664\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__32664\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__6515\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__6513\ : Span4Mux_v
    port map (
            O => \N__32655\,
            I => \N__32651\
        );

    \I__6512\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32648\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__32651\,
            I => scaler_4_data_12
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__32648\,
            I => scaler_4_data_12
        );

    \I__6509\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32640\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__32640\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__6507\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32630\
        );

    \I__6506\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32630\
        );

    \I__6505\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32627\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__32630\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__32627\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__32622\,
            I => \ppm_encoder_1.N_320_cascade_\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \N__32614\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__32618\,
            I => \N__32611\
        );

    \I__6499\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32606\
        );

    \I__6498\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32606\
        );

    \I__6497\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32603\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__32606\,
            I => \N__32600\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__32603\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__32600\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__6493\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32592\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32589\
        );

    \I__6491\ : Span4Mux_h
    port map (
            O => \N__32589\,
            I => \N__32585\
        );

    \I__6490\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32582\
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__32585\,
            I => throttle_command_9
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__32582\,
            I => throttle_command_9
        );

    \I__6487\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32574\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__32574\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__32571\,
            I => \N__32566\
        );

    \I__6484\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32559\
        );

    \I__6483\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32559\
        );

    \I__6482\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32559\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__32559\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__32556\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\
        );

    \I__6479\ : InMux
    port map (
            O => \N__32553\,
            I => \N__32550\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__32550\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__32547\,
            I => \N__32544\
        );

    \I__6476\ : InMux
    port map (
            O => \N__32544\,
            I => \N__32539\
        );

    \I__6475\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32534\
        );

    \I__6474\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32534\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__32539\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__32534\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__6471\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32525\
        );

    \I__6470\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32522\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32519\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__32522\,
            I => \N__32516\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__32519\,
            I => \N__32513\
        );

    \I__6466\ : Span4Mux_v
    port map (
            O => \N__32516\,
            I => \N__32510\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__32513\,
            I => scaler_3_data_12
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__32510\,
            I => scaler_3_data_12
        );

    \I__6463\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32502\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__32502\,
            I => \N__32499\
        );

    \I__6461\ : Span4Mux_h
    port map (
            O => \N__32499\,
            I => \N__32496\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__32496\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__6459\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32489\
        );

    \I__6458\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32486\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__32489\,
            I => \N__32483\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__32486\,
            I => \N__32480\
        );

    \I__6455\ : Span4Mux_h
    port map (
            O => \N__32483\,
            I => \N__32477\
        );

    \I__6454\ : Span4Mux_h
    port map (
            O => \N__32480\,
            I => \N__32474\
        );

    \I__6453\ : Span4Mux_h
    port map (
            O => \N__32477\,
            I => \N__32471\
        );

    \I__6452\ : Span4Mux_h
    port map (
            O => \N__32474\,
            I => \N__32468\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__32471\,
            I => throttle_command_12
        );

    \I__6450\ : Odrv4
    port map (
            O => \N__32468\,
            I => throttle_command_12
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__32463\,
            I => \N__32460\
        );

    \I__6448\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__32454\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__6445\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32447\
        );

    \I__6444\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32444\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32441\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32444\,
            I => \N__32438\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__32441\,
            I => \N__32435\
        );

    \I__6440\ : Span4Mux_h
    port map (
            O => \N__32438\,
            I => \N__32432\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__32435\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__32432\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__6436\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__32415\,
            I => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\
        );

    \I__6432\ : InMux
    port map (
            O => \N__32412\,
            I => \bfn_14_14_0_\
        );

    \I__6431\ : InMux
    port map (
            O => \N__32409\,
            I => \scaler_2.un2_source_data_0_cry_9\
        );

    \I__6430\ : CEMux
    port map (
            O => \N__32406\,
            I => \N__32385\
        );

    \I__6429\ : CEMux
    port map (
            O => \N__32405\,
            I => \N__32385\
        );

    \I__6428\ : CEMux
    port map (
            O => \N__32404\,
            I => \N__32385\
        );

    \I__6427\ : CEMux
    port map (
            O => \N__32403\,
            I => \N__32385\
        );

    \I__6426\ : CEMux
    port map (
            O => \N__32402\,
            I => \N__32385\
        );

    \I__6425\ : CEMux
    port map (
            O => \N__32401\,
            I => \N__32385\
        );

    \I__6424\ : CEMux
    port map (
            O => \N__32400\,
            I => \N__32385\
        );

    \I__6423\ : GlobalMux
    port map (
            O => \N__32385\,
            I => \N__32382\
        );

    \I__6422\ : gio2CtrlBuf
    port map (
            O => \N__32382\,
            I => \debug_CH3_20A_c_0_g\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__32379\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\
        );

    \I__6420\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__32373\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \ppm_encoder_1.N_301_cascade_\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32358\
        );

    \I__6416\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32358\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32365\,
            I => \N__32358\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__32358\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__6413\ : CascadeMux
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__6412\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32348\
        );

    \I__6411\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32345\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__32348\,
            I => \N__32342\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32339\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__32342\,
            I => \N__32336\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32333\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__32336\,
            I => scaler_3_data_9
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__32333\,
            I => scaler_3_data_9
        );

    \I__6404\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32325\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32325\,
            I => \N__32322\
        );

    \I__6402\ : Span4Mux_v
    port map (
            O => \N__32322\,
            I => \N__32319\
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__32319\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__32316\,
            I => \N__32311\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32304\
        );

    \I__6398\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32304\
        );

    \I__6397\ : InMux
    port map (
            O => \N__32311\,
            I => \N__32304\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__32304\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__6394\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32295\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__32295\,
            I => \N__32292\
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__32292\,
            I => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__32289\,
            I => \N__32286\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32279\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32279\
        );

    \I__6388\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32275\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32272\
        );

    \I__6386\ : InMux
    port map (
            O => \N__32278\,
            I => \N__32269\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__32275\,
            I => \N__32264\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__32272\,
            I => \N__32264\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__32269\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__32264\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32259\,
            I => \scaler_2.un2_source_data_0_cry_1\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32247\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32247\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__6376\ : Span4Mux_v
    port map (
            O => \N__32244\,
            I => \N__32241\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__32241\,
            I => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32238\,
            I => \scaler_2.un2_source_data_0_cry_2\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32226\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32226\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__6369\ : Span4Mux_v
    port map (
            O => \N__32223\,
            I => \N__32220\
        );

    \I__6368\ : Odrv4
    port map (
            O => \N__32220\,
            I => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\
        );

    \I__6367\ : InMux
    port map (
            O => \N__32217\,
            I => \scaler_2.un2_source_data_0_cry_3\
        );

    \I__6366\ : CascadeMux
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32205\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32205\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32202\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__32202\,
            I => \N__32199\
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__32199\,
            I => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32196\,
            I => \scaler_2.un2_source_data_0_cry_4\
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__32193\,
            I => \N__32190\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32184\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32184\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__32184\,
            I => \N__32181\
        );

    \I__6355\ : Span4Mux_h
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__6354\ : Odrv4
    port map (
            O => \N__32178\,
            I => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32175\,
            I => \scaler_2.un2_source_data_0_cry_5\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32163\
        );

    \I__6350\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32163\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__6348\ : Span4Mux_h
    port map (
            O => \N__32160\,
            I => \N__32157\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__32157\,
            I => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32154\,
            I => \scaler_2.un2_source_data_0_cry_6\
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32142\
        );

    \I__6343\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32142\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__6341\ : Span4Mux_h
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__32136\,
            I => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\
        );

    \I__6339\ : InMux
    port map (
            O => \N__32133\,
            I => \scaler_2.un2_source_data_0_cry_7\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__32130\,
            I => \N__32126\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32110\
        );

    \I__6336\ : InMux
    port map (
            O => \N__32126\,
            I => \N__32110\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32110\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32103\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32103\
        );

    \I__6332\ : InMux
    port map (
            O => \N__32122\,
            I => \N__32103\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32096\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32096\
        );

    \I__6329\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32096\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32091\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32091\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__32110\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__32103\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__32096\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__32091\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__32082\,
            I => \N__32077\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__32081\,
            I => \N__32068\
        );

    \I__6320\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32062\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32062\
        );

    \I__6318\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32055\
        );

    \I__6317\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32055\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32055\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32048\
        );

    \I__6314\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32048\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32048\
        );

    \I__6312\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32043\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32043\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__32062\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__32055\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__32048\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__32043\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__32034\,
            I => \N__32026\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32020\
        );

    \I__6304\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32013\
        );

    \I__6303\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32013\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32013\
        );

    \I__6301\ : InMux
    port map (
            O => \N__32029\,
            I => \N__32006\
        );

    \I__6300\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32006\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32006\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32001\
        );

    \I__6297\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32001\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__32020\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__32013\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__32006\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__32001\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__6292\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31989\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__6290\ : Span4Mux_h
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__31983\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__31980\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7_cascade_\
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__31977\,
            I => \ppm_encoder_1.N_299_cascade_\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__31974\,
            I => \N__31971\
        );

    \I__6285\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31966\
        );

    \I__6284\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31961\
        );

    \I__6283\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31961\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__31966\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__31961\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__6280\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31953\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31950\
        );

    \I__6278\ : Span4Mux_v
    port map (
            O => \N__31950\,
            I => \N__31947\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__31947\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__6276\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31940\
        );

    \I__6275\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31937\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31934\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31931\
        );

    \I__6272\ : Span4Mux_v
    port map (
            O => \N__31934\,
            I => \N__31928\
        );

    \I__6271\ : Span4Mux_v
    port map (
            O => \N__31931\,
            I => \N__31925\
        );

    \I__6270\ : Odrv4
    port map (
            O => \N__31928\,
            I => scaler_3_data_7
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__31925\,
            I => scaler_3_data_7
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__31920\,
            I => \N__31915\
        );

    \I__6267\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31908\
        );

    \I__6266\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31908\
        );

    \I__6265\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31908\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__31908\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__6263\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31902\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__31902\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__6260\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31893\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31889\
        );

    \I__6258\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31886\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__31889\,
            I => \N__31883\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31880\
        );

    \I__6255\ : Span4Mux_h
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__6254\ : Sp12to4
    port map (
            O => \N__31880\,
            I => \N__31874\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__31877\,
            I => throttle_command_7
        );

    \I__6252\ : Odrv12
    port map (
            O => \N__31874\,
            I => throttle_command_7
        );

    \I__6251\ : SRMux
    port map (
            O => \N__31869\,
            I => \N__31866\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__31863\,
            I => \N__31860\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__31860\,
            I => \N__31857\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__31857\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__31854\,
            I => \uart_pc.CO0_cascade_\
        );

    \I__6245\ : CascadeMux
    port map (
            O => \N__31851\,
            I => \N__31846\
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__31850\,
            I => \N__31843\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__31849\,
            I => \N__31839\
        );

    \I__6242\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31836\
        );

    \I__6241\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31829\
        );

    \I__6240\ : InMux
    port map (
            O => \N__31842\,
            I => \N__31829\
        );

    \I__6239\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31829\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31825\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31822\
        );

    \I__6236\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31819\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__31825\,
            I => \N__31814\
        );

    \I__6234\ : Span4Mux_h
    port map (
            O => \N__31822\,
            I => \N__31814\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__31819\,
            I => \N__31811\
        );

    \I__6232\ : Span4Mux_v
    port map (
            O => \N__31814\,
            I => \N__31807\
        );

    \I__6231\ : Span4Mux_h
    port map (
            O => \N__31811\,
            I => \N__31804\
        );

    \I__6230\ : InMux
    port map (
            O => \N__31810\,
            I => \N__31801\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__31807\,
            I => \N__31796\
        );

    \I__6228\ : Span4Mux_h
    port map (
            O => \N__31804\,
            I => \N__31796\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__31801\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__31796\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__6225\ : CEMux
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__31788\,
            I => \N__31785\
        );

    \I__6223\ : Span4Mux_h
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__6222\ : Sp12to4
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__6221\ : Span12Mux_v
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__6220\ : Odrv12
    port map (
            O => \N__31776\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\
        );

    \I__6219\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31769\
        );

    \I__6218\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31765\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31762\
        );

    \I__6216\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31759\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__31765\,
            I => \N__31754\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__31762\,
            I => \N__31754\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__31759\,
            I => \uart_pc.N_152\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__31754\,
            I => \uart_pc.N_152\
        );

    \I__6211\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31739\
        );

    \I__6210\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31739\
        );

    \I__6209\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31739\
        );

    \I__6208\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31736\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__31739\,
            I => \N__31731\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__31736\,
            I => \N__31731\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__31731\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \uart_pc.N_152_cascade_\
        );

    \I__6203\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31718\
        );

    \I__6202\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31715\
        );

    \I__6201\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31712\
        );

    \I__6200\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31704\
        );

    \I__6199\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31704\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__31718\,
            I => \N__31699\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31699\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__31712\,
            I => \N__31696\
        );

    \I__6195\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31693\
        );

    \I__6194\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31688\
        );

    \I__6193\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31688\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31683\
        );

    \I__6191\ : Span4Mux_v
    port map (
            O => \N__31699\,
            I => \N__31683\
        );

    \I__6190\ : Span4Mux_h
    port map (
            O => \N__31696\,
            I => \N__31680\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__31693\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__31688\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__31683\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__31680\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__6185\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31665\
        );

    \I__6184\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31665\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__31662\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__6181\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31655\
        );

    \I__6180\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31652\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__31655\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__31652\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__6177\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31644\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__31644\,
            I => \N__31639\
        );

    \I__6175\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31634\
        );

    \I__6174\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31634\
        );

    \I__6173\ : Span4Mux_v
    port map (
            O => \N__31639\,
            I => \N__31631\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__31634\,
            I => \N__31628\
        );

    \I__6171\ : Span4Mux_h
    port map (
            O => \N__31631\,
            I => \N__31623\
        );

    \I__6170\ : Span4Mux_v
    port map (
            O => \N__31628\,
            I => \N__31623\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__31623\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__6168\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31616\
        );

    \I__6167\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31612\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__31616\,
            I => \N__31608\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__31615\,
            I => \N__31602\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__31612\,
            I => \N__31598\
        );

    \I__6163\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31595\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__31608\,
            I => \N__31592\
        );

    \I__6161\ : InMux
    port map (
            O => \N__31607\,
            I => \N__31589\
        );

    \I__6160\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31584\
        );

    \I__6159\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31584\
        );

    \I__6158\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31579\
        );

    \I__6157\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31579\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__31598\,
            I => \N__31576\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__31595\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__31592\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__31589\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__31584\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__31579\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__31576\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__6149\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31559\
        );

    \I__6148\ : InMux
    port map (
            O => \N__31562\,
            I => \N__31556\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__31559\,
            I => \N__31551\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__31556\,
            I => \N__31548\
        );

    \I__6145\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31543\
        );

    \I__6144\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31540\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__31551\,
            I => \N__31535\
        );

    \I__6142\ : Span4Mux_h
    port map (
            O => \N__31548\,
            I => \N__31535\
        );

    \I__6141\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31530\
        );

    \I__6140\ : InMux
    port map (
            O => \N__31546\,
            I => \N__31530\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__31543\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__31540\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__31535\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__31530\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__31521\,
            I => \N__31516\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31513\
        );

    \I__6133\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31510\
        );

    \I__6132\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31506\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31500\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31497\
        );

    \I__6129\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31494\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__31506\,
            I => \N__31491\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__31505\,
            I => \N__31486\
        );

    \I__6126\ : InMux
    port map (
            O => \N__31504\,
            I => \N__31483\
        );

    \I__6125\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31480\
        );

    \I__6124\ : Span4Mux_v
    port map (
            O => \N__31500\,
            I => \N__31473\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__31497\,
            I => \N__31473\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__31494\,
            I => \N__31473\
        );

    \I__6121\ : Span4Mux_h
    port map (
            O => \N__31491\,
            I => \N__31470\
        );

    \I__6120\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31463\
        );

    \I__6119\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31463\
        );

    \I__6118\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31463\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__31483\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__31480\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__31473\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__31470\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__31463\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__6111\ : InMux
    port map (
            O => \N__31449\,
            I => \N__31445\
        );

    \I__6110\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31442\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31445\,
            I => \uart_drone.N_126_li\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__31442\,
            I => \uart_drone.N_126_li\
        );

    \I__6107\ : InMux
    port map (
            O => \N__31437\,
            I => \N__31413\
        );

    \I__6106\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31413\
        );

    \I__6105\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31413\
        );

    \I__6104\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31413\
        );

    \I__6103\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31413\
        );

    \I__6102\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31413\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31413\
        );

    \I__6100\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31413\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__31407\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__6096\ : IoInMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__6094\ : IoSpan4Mux
    port map (
            O => \N__31398\,
            I => \N__31394\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__31397\,
            I => \N__31385\
        );

    \I__6092\ : Span4Mux_s1_v
    port map (
            O => \N__31394\,
            I => \N__31379\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31376\
        );

    \I__6090\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31373\
        );

    \I__6089\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31359\
        );

    \I__6088\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31359\
        );

    \I__6087\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31359\
        );

    \I__6086\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31359\
        );

    \I__6085\ : InMux
    port map (
            O => \N__31385\,
            I => \N__31359\
        );

    \I__6084\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31352\
        );

    \I__6083\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31352\
        );

    \I__6082\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31352\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__31379\,
            I => \N__31345\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__31376\,
            I => \N__31345\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31345\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31342\
        );

    \I__6077\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31339\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31336\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31331\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31331\
        );

    \I__6073\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31326\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31326\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31323\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__31336\,
            I => \N__31320\
        );

    \I__6069\ : Span4Mux_v
    port map (
            O => \N__31331\,
            I => \N__31315\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__31326\,
            I => \N__31315\
        );

    \I__6067\ : Span4Mux_v
    port map (
            O => \N__31323\,
            I => \N__31310\
        );

    \I__6066\ : Span4Mux_h
    port map (
            O => \N__31320\,
            I => \N__31310\
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__31315\,
            I => \debug_CH0_16A_c\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__31310\,
            I => \debug_CH0_16A_c\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__31305\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31297\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__31301\,
            I => \N__31294\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31289\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31289\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31286\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__31289\,
            I => \N__31283\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__31286\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__31283\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__31272\,
            I => \N__31268\
        );

    \I__6051\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31265\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__31268\,
            I => \uart_pc.N_126_li\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__31265\,
            I => \uart_pc.N_126_li\
        );

    \I__6048\ : CascadeMux
    port map (
            O => \N__31260\,
            I => \uart_pc.state_srsts_0_0_0_cascade_\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__31254\,
            I => \uart_drone.state_srsts_0_0_0\
        );

    \I__6045\ : CascadeMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31241\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31238\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__31241\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__31238\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__31233\,
            I => \uart_drone.N_126_li_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31217\
        );

    \I__6037\ : IoInMux
    port map (
            O => \N__31229\,
            I => \N__31213\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31209\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31200\
        );

    \I__6034\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31200\
        );

    \I__6033\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31200\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31200\
        );

    \I__6031\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31191\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31191\
        );

    \I__6029\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31191\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31191\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31188\
        );

    \I__6026\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31185\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__31213\,
            I => \N__31182\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31179\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31175\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31170\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31170\
        );

    \I__6020\ : Span4Mux_v
    port map (
            O => \N__31188\,
            I => \N__31165\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31185\,
            I => \N__31165\
        );

    \I__6018\ : Span4Mux_s2_v
    port map (
            O => \N__31182\,
            I => \N__31162\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31159\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31156\
        );

    \I__6015\ : Span4Mux_v
    port map (
            O => \N__31175\,
            I => \N__31149\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__31170\,
            I => \N__31149\
        );

    \I__6013\ : Span4Mux_h
    port map (
            O => \N__31165\,
            I => \N__31149\
        );

    \I__6012\ : Span4Mux_h
    port map (
            O => \N__31162\,
            I => \N__31144\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__31159\,
            I => \N__31144\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__31156\,
            I => \N__31141\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__31149\,
            I => \debug_CH2_18A_c\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__31144\,
            I => \debug_CH2_18A_c\
        );

    \I__6007\ : Odrv12
    port map (
            O => \N__31141\,
            I => \debug_CH2_18A_c\
        );

    \I__6006\ : CascadeMux
    port map (
            O => \N__31134\,
            I => \uart_pc.state_srsts_i_0_2_cascade_\
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__31131\,
            I => \N__31126\
        );

    \I__6004\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31123\
        );

    \I__6003\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31118\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31118\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__31123\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__31118\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__31113\,
            I => \N__31109\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__31112\,
            I => \N__31105\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31102\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31098\
        );

    \I__5995\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31095\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31102\,
            I => \N__31092\
        );

    \I__5993\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31089\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31084\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31084\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__31092\,
            I => \N__31081\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__31089\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__31084\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__31081\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__31074\,
            I => \N__31069\
        );

    \I__5985\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31064\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31061\
        );

    \I__5983\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31053\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31053\
        );

    \I__5981\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31053\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__31064\,
            I => \N__31047\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__31061\,
            I => \N__31047\
        );

    \I__5978\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31044\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__31053\,
            I => \N__31040\
        );

    \I__5976\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31037\
        );

    \I__5975\ : Span4Mux_h
    port map (
            O => \N__31047\,
            I => \N__31032\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31032\
        );

    \I__5973\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31029\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__31040\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__31037\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__31032\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__31029\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__31020\,
            I => \N__31016\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__31019\,
            I => \N__31013\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31010\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31007\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__31010\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__31007\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30996\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__31001\,
            I => \N__30993\
        );

    \I__5960\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30987\
        );

    \I__5959\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30984\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30981\
        );

    \I__5957\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30978\
        );

    \I__5956\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30975\
        );

    \I__5955\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30970\
        );

    \I__5954\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30970\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30967\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30962\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__30981\,
            I => \N__30962\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__30978\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__30975\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__30970\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__30967\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__30962\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__5945\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30945\
        );

    \I__5944\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30945\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30941\
        );

    \I__5942\ : InMux
    port map (
            O => \N__30944\,
            I => \N__30938\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__30941\,
            I => \N__30935\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__30938\,
            I => \N__30932\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__30935\,
            I => \N__30929\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__30932\,
            I => \N__30926\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__30929\,
            I => \N__30923\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__30926\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__30923\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__5934\ : InMux
    port map (
            O => \N__30918\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_14\
        );

    \I__5933\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30908\
        );

    \I__5932\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30908\
        );

    \I__5931\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30905\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__30908\,
            I => \N__30902\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__30905\,
            I => \N__30899\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__30902\,
            I => \N__30896\
        );

    \I__5927\ : Span4Mux_h
    port map (
            O => \N__30899\,
            I => \N__30891\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__30896\,
            I => \N__30891\
        );

    \I__5925\ : Sp12to4
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__5924\ : Odrv12
    port map (
            O => \N__30888\,
            I => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\
        );

    \I__5923\ : InMux
    port map (
            O => \N__30885\,
            I => \bfn_13_23_0_\
        );

    \I__5922\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30876\
        );

    \I__5921\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30876\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30872\
        );

    \I__5919\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30869\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__30872\,
            I => \N__30866\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__30869\,
            I => \N__30863\
        );

    \I__5916\ : Span4Mux_v
    port map (
            O => \N__30866\,
            I => \N__30860\
        );

    \I__5915\ : Span4Mux_h
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__5914\ : Span4Mux_h
    port map (
            O => \N__30860\,
            I => \N__30854\
        );

    \I__5913\ : Odrv4
    port map (
            O => \N__30857\,
            I => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\
        );

    \I__5912\ : Odrv4
    port map (
            O => \N__30854\,
            I => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\
        );

    \I__5911\ : InMux
    port map (
            O => \N__30849\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_16\
        );

    \I__5910\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30840\
        );

    \I__5909\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30840\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__30840\,
            I => \N__30836\
        );

    \I__5907\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30833\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__30836\,
            I => \N__30830\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__30833\,
            I => \N__30827\
        );

    \I__5904\ : Sp12to4
    port map (
            O => \N__30830\,
            I => \N__30824\
        );

    \I__5903\ : Span4Mux_h
    port map (
            O => \N__30827\,
            I => \N__30821\
        );

    \I__5902\ : Span12Mux_v
    port map (
            O => \N__30824\,
            I => \N__30818\
        );

    \I__5901\ : Odrv4
    port map (
            O => \N__30821\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__5900\ : Odrv12
    port map (
            O => \N__30818\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__5899\ : InMux
    port map (
            O => \N__30813\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_17\
        );

    \I__5898\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30804\
        );

    \I__5897\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30804\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__5895\ : Span4Mux_h
    port map (
            O => \N__30801\,
            I => \N__30797\
        );

    \I__5894\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30794\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__30797\,
            I => \N__30791\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30788\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__30791\,
            I => \N__30785\
        );

    \I__5890\ : Span4Mux_h
    port map (
            O => \N__30788\,
            I => \N__30782\
        );

    \I__5889\ : Span4Mux_h
    port map (
            O => \N__30785\,
            I => \N__30779\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__30782\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__30779\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__5886\ : InMux
    port map (
            O => \N__30774\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_18\
        );

    \I__5885\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30767\
        );

    \I__5884\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30763\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30760\
        );

    \I__5882\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30757\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30754\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__30760\,
            I => \N__30751\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__30757\,
            I => \N__30748\
        );

    \I__5878\ : Span4Mux_v
    port map (
            O => \N__30754\,
            I => \N__30745\
        );

    \I__5877\ : Sp12to4
    port map (
            O => \N__30751\,
            I => \N__30742\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__30748\,
            I => \N__30739\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__30745\,
            I => \N__30736\
        );

    \I__5874\ : Span12Mux_v
    port map (
            O => \N__30742\,
            I => \N__30733\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__30739\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__30736\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__5871\ : Odrv12
    port map (
            O => \N__30733\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__5870\ : InMux
    port map (
            O => \N__30726\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19\
        );

    \I__5869\ : InMux
    port map (
            O => \N__30723\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20\
        );

    \I__5868\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30714\
        );

    \I__5867\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30707\
        );

    \I__5866\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30707\
        );

    \I__5865\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30707\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__30714\,
            I => \N__30691\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__30707\,
            I => \N__30687\
        );

    \I__5862\ : InMux
    port map (
            O => \N__30706\,
            I => \N__30684\
        );

    \I__5861\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30681\
        );

    \I__5860\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30676\
        );

    \I__5859\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30676\
        );

    \I__5858\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30667\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30667\
        );

    \I__5856\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30667\
        );

    \I__5855\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30667\
        );

    \I__5854\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30664\
        );

    \I__5853\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30655\
        );

    \I__5852\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30655\
        );

    \I__5851\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30655\
        );

    \I__5850\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30655\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__30691\,
            I => \N__30652\
        );

    \I__5848\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30648\
        );

    \I__5847\ : Span4Mux_h
    port map (
            O => \N__30687\,
            I => \N__30645\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__30684\,
            I => \N__30642\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__30681\,
            I => \N__30639\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30636\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__30667\,
            I => \N__30629\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30629\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30629\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__30652\,
            I => \N__30626\
        );

    \I__5839\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30623\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30618\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__30645\,
            I => \N__30618\
        );

    \I__5836\ : Span4Mux_h
    port map (
            O => \N__30642\,
            I => \N__30615\
        );

    \I__5835\ : Span4Mux_h
    port map (
            O => \N__30639\,
            I => \N__30612\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__30636\,
            I => \N__30607\
        );

    \I__5833\ : Span4Mux_v
    port map (
            O => \N__30629\,
            I => \N__30607\
        );

    \I__5832\ : Span4Mux_h
    port map (
            O => \N__30626\,
            I => \N__30604\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__30623\,
            I => \N__30601\
        );

    \I__5830\ : Span4Mux_h
    port map (
            O => \N__30618\,
            I => \N__30598\
        );

    \I__5829\ : Span4Mux_h
    port map (
            O => \N__30615\,
            I => \N__30593\
        );

    \I__5828\ : Span4Mux_v
    port map (
            O => \N__30612\,
            I => \N__30593\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__30607\,
            I => \N__30590\
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__30604\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__5825\ : Odrv12
    port map (
            O => \N__30601\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__5824\ : Odrv4
    port map (
            O => \N__30598\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__30593\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__30590\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__5821\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30574\
        );

    \I__5820\ : IoInMux
    port map (
            O => \N__30578\,
            I => \N__30571\
        );

    \I__5819\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30568\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30563\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30560\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30557\
        );

    \I__5815\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30552\
        );

    \I__5814\ : InMux
    port map (
            O => \N__30566\,
            I => \N__30552\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__30563\,
            I => \N__30549\
        );

    \I__5812\ : Span4Mux_s1_v
    port map (
            O => \N__30560\,
            I => \N__30546\
        );

    \I__5811\ : Span4Mux_v
    port map (
            O => \N__30557\,
            I => \N__30543\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30540\
        );

    \I__5809\ : Span4Mux_h
    port map (
            O => \N__30549\,
            I => \N__30537\
        );

    \I__5808\ : Span4Mux_v
    port map (
            O => \N__30546\,
            I => \N__30534\
        );

    \I__5807\ : Span4Mux_v
    port map (
            O => \N__30543\,
            I => \N__30529\
        );

    \I__5806\ : Span4Mux_h
    port map (
            O => \N__30540\,
            I => \N__30529\
        );

    \I__5805\ : Sp12to4
    port map (
            O => \N__30537\,
            I => \N__30525\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__30534\,
            I => \N__30520\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__30529\,
            I => \N__30520\
        );

    \I__5802\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30517\
        );

    \I__5801\ : Span12Mux_v
    port map (
            O => \N__30525\,
            I => \N__30514\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__30520\,
            I => \debug_CH3_20A_c\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__30517\,
            I => \debug_CH3_20A_c\
        );

    \I__5798\ : Odrv12
    port map (
            O => \N__30514\,
            I => \debug_CH3_20A_c\
        );

    \I__5797\ : IoInMux
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__30501\,
            I => \debug_CH3_20A_c_0\
        );

    \I__5794\ : InMux
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__30495\,
            I => \N__30491\
        );

    \I__5792\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30488\
        );

    \I__5791\ : Span4Mux_h
    port map (
            O => \N__30491\,
            I => \N__30485\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30488\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__30485\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__5788\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30476\
        );

    \I__5787\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30472\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30469\
        );

    \I__5785\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30466\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30463\
        );

    \I__5783\ : Span4Mux_v
    port map (
            O => \N__30469\,
            I => \N__30460\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30455\
        );

    \I__5781\ : Span12Mux_v
    port map (
            O => \N__30463\,
            I => \N__30455\
        );

    \I__5780\ : Span4Mux_h
    port map (
            O => \N__30460\,
            I => \N__30452\
        );

    \I__5779\ : Odrv12
    port map (
            O => \N__30455\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__5778\ : Odrv4
    port map (
            O => \N__30452\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__5777\ : InMux
    port map (
            O => \N__30447\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6\
        );

    \I__5776\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30440\
        );

    \I__5775\ : InMux
    port map (
            O => \N__30443\,
            I => \N__30437\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__30440\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__30437\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__5772\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30426\
        );

    \I__5771\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30426\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__5768\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30416\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__30416\,
            I => \N__30410\
        );

    \I__5765\ : Span4Mux_h
    port map (
            O => \N__30413\,
            I => \N__30407\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__30410\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__30407\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__5762\ : InMux
    port map (
            O => \N__30402\,
            I => \bfn_13_22_0_\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__30399\,
            I => \N__30396\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30392\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__30395\,
            I => \N__30389\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__30392\,
            I => \N__30386\
        );

    \I__5757\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30383\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__30386\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__30383\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30371\
        );

    \I__5753\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30368\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__30371\,
            I => \N__30365\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30360\
        );

    \I__5749\ : Span12Mux_v
    port map (
            O => \N__30365\,
            I => \N__30360\
        );

    \I__5748\ : Odrv12
    port map (
            O => \N__30360\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\
        );

    \I__5747\ : InMux
    port map (
            O => \N__30357\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__5745\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30347\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30344\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__30347\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__30344\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__5741\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30335\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30331\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N__30328\
        );

    \I__5738\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30325\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__30331\,
            I => \N__30320\
        );

    \I__5736\ : Span4Mux_h
    port map (
            O => \N__30328\,
            I => \N__30320\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30317\
        );

    \I__5734\ : Span4Mux_v
    port map (
            O => \N__30320\,
            I => \N__30314\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__30317\,
            I => \N__30311\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__30314\,
            I => \N__30308\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__30311\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__30308\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30303\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30293\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30293\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30290\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__30293\,
            I => \N__30287\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__30290\,
            I => \N__30284\
        );

    \I__5723\ : Sp12to4
    port map (
            O => \N__30287\,
            I => \N__30281\
        );

    \I__5722\ : Span4Mux_h
    port map (
            O => \N__30284\,
            I => \N__30278\
        );

    \I__5721\ : Span12Mux_v
    port map (
            O => \N__30281\,
            I => \N__30275\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__30278\,
            I => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\
        );

    \I__5719\ : Odrv12
    port map (
            O => \N__30275\,
            I => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30270\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_10\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30263\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30260\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30263\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30260\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30255\,
            I => \N__30251\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30247\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30244\
        );

    \I__5710\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30241\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__30247\,
            I => \N__30238\
        );

    \I__5708\ : Sp12to4
    port map (
            O => \N__30244\,
            I => \N__30233\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30241\,
            I => \N__30233\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__30238\,
            I => \N__30230\
        );

    \I__5705\ : Span12Mux_v
    port map (
            O => \N__30233\,
            I => \N__30227\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__30230\,
            I => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\
        );

    \I__5703\ : Odrv12
    port map (
            O => \N__30227\,
            I => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30222\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_11\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30216\,
            I => \N__30211\
        );

    \I__5699\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30206\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30206\
        );

    \I__5697\ : Span4Mux_h
    port map (
            O => \N__30211\,
            I => \N__30203\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__30206\,
            I => \N__30200\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__30203\,
            I => \N__30197\
        );

    \I__5694\ : Span12Mux_v
    port map (
            O => \N__30200\,
            I => \N__30194\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__30197\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__5692\ : Odrv12
    port map (
            O => \N__30194\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30189\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_12\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30180\
        );

    \I__5689\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30180\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30180\,
            I => \N__30176\
        );

    \I__5687\ : InMux
    port map (
            O => \N__30179\,
            I => \N__30173\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__30176\,
            I => \N__30170\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__30173\,
            I => \N__30167\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__30170\,
            I => \N__30164\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__30167\,
            I => \N__30159\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__30164\,
            I => \N__30159\
        );

    \I__5681\ : Odrv4
    port map (
            O => \N__30159\,
            I => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\
        );

    \I__5680\ : InMux
    port map (
            O => \N__30156\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_13\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__30144\,
            I => scaler_3_data_14
        );

    \I__5675\ : InMux
    port map (
            O => \N__30141\,
            I => \bfn_13_20_0_\
        );

    \I__5674\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30134\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30131\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30128\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30125\
        );

    \I__5670\ : Span4Mux_v
    port map (
            O => \N__30128\,
            I => \N__30120\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30120\
        );

    \I__5668\ : Span4Mux_h
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__30111\,
            I => \pid_alt.un1_pid_prereg_0\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30105\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__30105\,
            I => \pid_alt.error_i_acummZ0Z_1\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__30102\,
            I => \N__30098\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__30101\,
            I => \N__30095\
        );

    \I__5660\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30092\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30089\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30086\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30082\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__30086\,
            I => \N__30079\
        );

    \I__5655\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30076\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__30082\,
            I => \N__30073\
        );

    \I__5653\ : Sp12to4
    port map (
            O => \N__30079\,
            I => \N__30070\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__30076\,
            I => \N__30067\
        );

    \I__5651\ : Span4Mux_v
    port map (
            O => \N__30073\,
            I => \N__30064\
        );

    \I__5650\ : Span12Mux_v
    port map (
            O => \N__30070\,
            I => \N__30061\
        );

    \I__5649\ : Span4Mux_h
    port map (
            O => \N__30067\,
            I => \N__30058\
        );

    \I__5648\ : Span4Mux_h
    port map (
            O => \N__30064\,
            I => \N__30055\
        );

    \I__5647\ : Odrv12
    port map (
            O => \N__30061\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__30058\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__30055\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30048\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_0\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__30042\,
            I => \pid_alt.error_i_acummZ0Z_2\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30036\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__30036\,
            I => \N__30032\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30029\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__30032\,
            I => \N__30025\
        );

    \I__5637\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30022\
        );

    \I__5636\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30019\
        );

    \I__5635\ : Sp12to4
    port map (
            O => \N__30025\,
            I => \N__30014\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__30022\,
            I => \N__30014\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__30019\,
            I => \N__30009\
        );

    \I__5632\ : Span12Mux_v
    port map (
            O => \N__30014\,
            I => \N__30009\
        );

    \I__5631\ : Odrv12
    port map (
            O => \N__30009\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__5630\ : InMux
    port map (
            O => \N__30006\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_1\
        );

    \I__5629\ : InMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30000\,
            I => \pid_alt.error_i_acummZ0Z_3\
        );

    \I__5627\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29993\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__29993\,
            I => \N__29986\
        );

    \I__5624\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29983\
        );

    \I__5623\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29980\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__29986\,
            I => \N__29975\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__29983\,
            I => \N__29975\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__29980\,
            I => \N__29972\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__29975\,
            I => \N__29969\
        );

    \I__5618\ : Span4Mux_v
    port map (
            O => \N__29972\,
            I => \N__29964\
        );

    \I__5617\ : Span4Mux_v
    port map (
            O => \N__29969\,
            I => \N__29964\
        );

    \I__5616\ : Span4Mux_h
    port map (
            O => \N__29964\,
            I => \N__29961\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__29961\,
            I => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\
        );

    \I__5614\ : InMux
    port map (
            O => \N__29958\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_2\
        );

    \I__5613\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29952\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__29952\,
            I => \pid_alt.error_i_acummZ0Z_4\
        );

    \I__5611\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29940\
        );

    \I__5610\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29940\
        );

    \I__5609\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29940\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29937\
        );

    \I__5607\ : Span4Mux_h
    port map (
            O => \N__29937\,
            I => \N__29934\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__29934\,
            I => \N__29931\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__29931\,
            I => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\
        );

    \I__5604\ : InMux
    port map (
            O => \N__29928\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_3\
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__29925\,
            I => \N__29921\
        );

    \I__5602\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29918\
        );

    \I__5601\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__29918\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__29915\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__5598\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29907\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__29907\,
            I => \N__29902\
        );

    \I__5596\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29897\
        );

    \I__5595\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29897\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__29902\,
            I => \N__29894\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29891\
        );

    \I__5592\ : Sp12to4
    port map (
            O => \N__29894\,
            I => \N__29886\
        );

    \I__5591\ : Span12Mux_h
    port map (
            O => \N__29891\,
            I => \N__29886\
        );

    \I__5590\ : Odrv12
    port map (
            O => \N__29886\,
            I => \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\
        );

    \I__5589\ : InMux
    port map (
            O => \N__29883\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_4\
        );

    \I__5588\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29874\
        );

    \I__5587\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29874\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29871\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__29871\,
            I => \N__29867\
        );

    \I__5584\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29864\
        );

    \I__5583\ : Span4Mux_v
    port map (
            O => \N__29867\,
            I => \N__29861\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__29864\,
            I => \N__29858\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__29861\,
            I => \N__29855\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__29858\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__29855\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__5578\ : InMux
    port map (
            O => \N__29850\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5\
        );

    \I__5577\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29844\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__29844\,
            I => scaler_4_data_14
        );

    \I__5575\ : InMux
    port map (
            O => \N__29841\,
            I => \bfn_13_18_0_\
        );

    \I__5574\ : InMux
    port map (
            O => \N__29838\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__5573\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29831\
        );

    \I__5572\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29828\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__29831\,
            I => \N__29825\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29820\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__29825\,
            I => \N__29820\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__29820\,
            I => scaler_3_data_8
        );

    \I__5567\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29814\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__5565\ : Odrv12
    port map (
            O => \N__29811\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__5564\ : InMux
    port map (
            O => \N__29808\,
            I => \ppm_encoder_1.un1_elevator_cry_7\
        );

    \I__5563\ : InMux
    port map (
            O => \N__29805\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__5562\ : InMux
    port map (
            O => \N__29802\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__5561\ : InMux
    port map (
            O => \N__29799\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__5560\ : InMux
    port map (
            O => \N__29796\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__5559\ : InMux
    port map (
            O => \N__29793\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__5558\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29786\
        );

    \I__5557\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29783\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__29786\,
            I => scaler_4_data_6
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__29783\,
            I => scaler_4_data_6
        );

    \I__5554\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29774\
        );

    \I__5553\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29771\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__29774\,
            I => scaler_4_data_7
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__29771\,
            I => scaler_4_data_7
        );

    \I__5550\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__29763\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__5548\ : InMux
    port map (
            O => \N__29760\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__5547\ : InMux
    port map (
            O => \N__29757\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__5546\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29750\
        );

    \I__5545\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29747\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__29750\,
            I => scaler_4_data_9
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__29747\,
            I => scaler_4_data_9
        );

    \I__5542\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__29739\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__5540\ : InMux
    port map (
            O => \N__29736\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__5539\ : InMux
    port map (
            O => \N__29733\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__5538\ : InMux
    port map (
            O => \N__29730\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__5537\ : InMux
    port map (
            O => \N__29727\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__5536\ : InMux
    port map (
            O => \N__29724\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__5535\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29718\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__29715\,
            I => \N__29709\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29706\
        );

    \I__5531\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29701\
        );

    \I__5530\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29698\
        );

    \I__5529\ : Span4Mux_h
    port map (
            O => \N__29709\,
            I => \N__29695\
        );

    \I__5528\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29688\
        );

    \I__5527\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29688\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29688\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29683\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29683\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__29695\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__29688\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__29683\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5520\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29673\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__29673\,
            I => \N__29669\
        );

    \I__5518\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29664\
        );

    \I__5517\ : Span4Mux_v
    port map (
            O => \N__29669\,
            I => \N__29658\
        );

    \I__5516\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29654\
        );

    \I__5515\ : InMux
    port map (
            O => \N__29667\,
            I => \N__29651\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__29664\,
            I => \N__29648\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__29663\,
            I => \N__29644\
        );

    \I__5512\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29637\
        );

    \I__5511\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29637\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__29658\,
            I => \N__29634\
        );

    \I__5509\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29631\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__29654\,
            I => \N__29628\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__29651\,
            I => \N__29623\
        );

    \I__5506\ : Span4Mux_h
    port map (
            O => \N__29648\,
            I => \N__29623\
        );

    \I__5505\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29614\
        );

    \I__5504\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29614\
        );

    \I__5503\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29614\
        );

    \I__5502\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29614\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__29637\,
            I => uart_drone_data_rdy
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__29634\,
            I => uart_drone_data_rdy
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__29631\,
            I => uart_drone_data_rdy
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__29628\,
            I => uart_drone_data_rdy
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__29623\,
            I => uart_drone_data_rdy
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__29614\,
            I => uart_drone_data_rdy
        );

    \I__5495\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29597\
        );

    \I__5494\ : IoInMux
    port map (
            O => \N__29600\,
            I => \N__29594\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29591\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__29594\,
            I => \N__29587\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__29591\,
            I => \N__29584\
        );

    \I__5490\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29581\
        );

    \I__5489\ : Span12Mux_s2_v
    port map (
            O => \N__29587\,
            I => \N__29578\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__29584\,
            I => \N__29572\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29572\
        );

    \I__5486\ : Span12Mux_v
    port map (
            O => \N__29578\,
            I => \N__29569\
        );

    \I__5485\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29566\
        );

    \I__5484\ : Span4Mux_h
    port map (
            O => \N__29572\,
            I => \N__29563\
        );

    \I__5483\ : Odrv12
    port map (
            O => \N__29569\,
            I => \debug_CH1_0A_c\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__29566\,
            I => \debug_CH1_0A_c\
        );

    \I__5481\ : Odrv4
    port map (
            O => \N__29563\,
            I => \debug_CH1_0A_c\
        );

    \I__5480\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29547\
        );

    \I__5478\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29544\
        );

    \I__5477\ : InMux
    port map (
            O => \N__29551\,
            I => \N__29541\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__29550\,
            I => \N__29538\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__29547\,
            I => \N__29535\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__29544\,
            I => \N__29532\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29529\
        );

    \I__5472\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29526\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__29535\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__29532\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__29529\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__29526\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5467\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29514\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__29514\,
            I => \N__29509\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29506\
        );

    \I__5464\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29503\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__29509\,
            I => \N__29500\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29497\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29494\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__29500\,
            I => \N__29488\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__29497\,
            I => \N__29488\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__29494\,
            I => \N__29485\
        );

    \I__5457\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29482\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__29488\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__29485\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__29482\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5453\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29471\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__29474\,
            I => \N__29468\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__5450\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29462\
        );

    \I__5449\ : Odrv12
    port map (
            O => \N__29465\,
            I => scaler_4_data_4
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__29462\,
            I => scaler_4_data_4
        );

    \I__5447\ : IoInMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29450\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__29453\,
            I => \N__29447\
        );

    \I__5444\ : Span12Mux_s3_v
    port map (
            O => \N__29450\,
            I => \N__29444\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29441\
        );

    \I__5442\ : Odrv12
    port map (
            O => \N__29444\,
            I => ppm_output_c
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__29441\,
            I => ppm_output_c
        );

    \I__5440\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29432\
        );

    \I__5439\ : InMux
    port map (
            O => \N__29435\,
            I => \N__29429\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__29432\,
            I => \N__29424\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29429\,
            I => \N__29424\
        );

    \I__5436\ : Span4Mux_v
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__29421\,
            I => throttle_command_10
        );

    \I__5434\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29415\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5432\ : Odrv4
    port map (
            O => \N__29412\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29406\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__29406\,
            I => \N__29403\
        );

    \I__5429\ : Odrv12
    port map (
            O => \N__29403\,
            I => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29397\,
            I => \N__29393\
        );

    \I__5426\ : CascadeMux
    port map (
            O => \N__29396\,
            I => \N__29389\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__29393\,
            I => \N__29386\
        );

    \I__5424\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29383\
        );

    \I__5423\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29380\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__29386\,
            I => \N__29377\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__29383\,
            I => \N__29374\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__29380\,
            I => throttle_command_4
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__29377\,
            I => throttle_command_4
        );

    \I__5418\ : Odrv12
    port map (
            O => \N__29374\,
            I => throttle_command_4
        );

    \I__5417\ : InMux
    port map (
            O => \N__29367\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__5416\ : InMux
    port map (
            O => \N__29364\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__5415\ : InMux
    port map (
            O => \N__29361\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__5414\ : InMux
    port map (
            O => \N__29358\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__5413\ : InMux
    port map (
            O => \N__29355\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29352\,
            I => \ppm_encoder_1.un1_throttle_cry_13\
        );

    \I__5411\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29342\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__29345\,
            I => \N__29338\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__29342\,
            I => \N__29335\
        );

    \I__5407\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29332\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29329\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__29335\,
            I => \N__29324\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29332\,
            I => \N__29324\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__29329\,
            I => throttle_command_2
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__29324\,
            I => throttle_command_2
        );

    \I__5401\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__29313\,
            I => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__29304\,
            I => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29297\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__29300\,
            I => \N__29293\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__29297\,
            I => \N__29290\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29287\
        );

    \I__5391\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29284\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__29290\,
            I => \N__29281\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__29287\,
            I => \N__29278\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__29284\,
            I => throttle_command_1
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__29281\,
            I => throttle_command_1
        );

    \I__5386\ : Odrv4
    port map (
            O => \N__29278\,
            I => throttle_command_1
        );

    \I__5385\ : InMux
    port map (
            O => \N__29271\,
            I => \ppm_encoder_1.un1_throttle_cry_0\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29268\,
            I => \ppm_encoder_1.un1_throttle_cry_1\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29265\,
            I => \ppm_encoder_1.un1_throttle_cry_2\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29262\,
            I => \ppm_encoder_1.un1_throttle_cry_3\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29255\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29252\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29255\,
            I => \N__29249\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__29249\,
            I => \N__29243\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__29246\,
            I => \N__29240\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__29243\,
            I => throttle_command_5
        );

    \I__5374\ : Odrv4
    port map (
            O => \N__29240\,
            I => throttle_command_5
        );

    \I__5373\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__29232\,
            I => \N__29229\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__29229\,
            I => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29226\,
            I => \ppm_encoder_1.un1_throttle_cry_4\
        );

    \I__5369\ : InMux
    port map (
            O => \N__29223\,
            I => \ppm_encoder_1.un1_throttle_cry_5\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29220\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__5367\ : InMux
    port map (
            O => \N__29217\,
            I => \bfn_13_14_0_\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29211\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__29211\,
            I => \N__29208\
        );

    \I__5364\ : Odrv12
    port map (
            O => \N__29208\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__29205\,
            I => \N__29202\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29199\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29199\,
            I => \N__29196\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__29196\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__5359\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29190\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__29190\,
            I => \N__29187\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__29187\,
            I => \N__29184\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__29184\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29177\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__29180\,
            I => \N__29174\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29171\
        );

    \I__5352\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29168\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__29171\,
            I => scaler_2_data_4
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__29168\,
            I => scaler_2_data_4
        );

    \I__5349\ : InMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29160\,
            I => scaler_2_data_5
        );

    \I__5347\ : InMux
    port map (
            O => \N__29157\,
            I => \N__29153\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__29156\,
            I => \N__29150\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29150\,
            I => \N__29144\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__29147\,
            I => scaler_3_data_4
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29144\,
            I => scaler_3_data_4
        );

    \I__5341\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__29136\,
            I => scaler_3_data_5
        );

    \I__5339\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__29130\,
            I => scaler_4_data_5
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29120\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29117\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__29117\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__29114\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__5331\ : SRMux
    port map (
            O => \N__29109\,
            I => \N__29106\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__5329\ : Odrv12
    port map (
            O => \N__29103\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29097\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29097\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29091\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__29091\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__5324\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29085\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29085\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__5322\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29076\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__29081\,
            I => \N__29073\
        );

    \I__5320\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29070\
        );

    \I__5319\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29067\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29064\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29061\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__29070\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__29067\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5314\ : Odrv12
    port map (
            O => \N__29064\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29061\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__5312\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29048\
        );

    \I__5311\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29045\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__29048\,
            I => \N__29039\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__29045\,
            I => \N__29039\
        );

    \I__5308\ : InMux
    port map (
            O => \N__29044\,
            I => \N__29036\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__29039\,
            I => \N__29032\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29029\
        );

    \I__5305\ : InMux
    port map (
            O => \N__29035\,
            I => \N__29026\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__29032\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__29029\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__29026\,
            I => \frame_decoder_CH2data_0\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29011\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__29015\,
            I => \N__29008\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29014\,
            I => \N__29004\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__29011\,
            I => \N__29001\
        );

    \I__5296\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28996\
        );

    \I__5295\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28996\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__29004\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__29001\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__28996\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__5291\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28985\
        );

    \I__5290\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28975\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28975\
        );

    \I__5287\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28972\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__28980\,
            I => \N__28969\
        );

    \I__5285\ : Span4Mux_v
    port map (
            O => \N__28975\,
            I => \N__28966\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28963\
        );

    \I__5283\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28960\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__28966\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__28963\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__28960\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__5279\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28949\
        );

    \I__5278\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28946\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__28949\,
            I => \N__28939\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28939\
        );

    \I__5275\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28936\
        );

    \I__5274\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28933\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__28939\,
            I => \N__28930\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28927\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28924\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__28930\,
            I => \frame_decoder_CH3data_0\
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__28927\,
            I => \frame_decoder_CH3data_0\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__28924\,
            I => \frame_decoder_CH3data_0\
        );

    \I__5267\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N__28910\
        );

    \I__5265\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28906\
        );

    \I__5264\ : Span4Mux_v
    port map (
            O => \N__28910\,
            I => \N__28903\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__28909\,
            I => \N__28900\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28896\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__28903\,
            I => \N__28893\
        );

    \I__5260\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28888\
        );

    \I__5259\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28888\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__28896\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__28893\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__28888\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__28881\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__28878\,
            I => \N__28875\
        );

    \I__5253\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28871\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__28874\,
            I => \N__28868\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__28871\,
            I => \N__28865\
        );

    \I__5250\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28862\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__28865\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__28862\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__28857\,
            I => \N__28854\
        );

    \I__5246\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28850\
        );

    \I__5245\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28847\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__28850\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__28847\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28838\
        );

    \I__5241\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28835\
        );

    \I__5240\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28832\
        );

    \I__5239\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28829\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__28832\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__28829\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__28824\,
            I => \N__28821\
        );

    \I__5235\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28814\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__28817\,
            I => \N__28811\
        );

    \I__5232\ : Span4Mux_v
    port map (
            O => \N__28814\,
            I => \N__28808\
        );

    \I__5231\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28805\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__28808\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__28805\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__28800\,
            I => \N__28796\
        );

    \I__5227\ : CascadeMux
    port map (
            O => \N__28799\,
            I => \N__28793\
        );

    \I__5226\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28790\
        );

    \I__5225\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28787\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__28790\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__28787\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__28782\,
            I => \N__28778\
        );

    \I__5221\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__5220\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28772\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__28775\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__28772\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__5217\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28743\
        );

    \I__5216\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28743\
        );

    \I__5215\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28743\
        );

    \I__5214\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28743\
        );

    \I__5213\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28743\
        );

    \I__5212\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28743\
        );

    \I__5211\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28743\
        );

    \I__5210\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28743\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__28737\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__5206\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28729\
        );

    \I__5205\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28724\
        );

    \I__5204\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28724\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__28729\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__28724\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__5201\ : CascadeMux
    port map (
            O => \N__28719\,
            I => \N__28714\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__28718\,
            I => \N__28711\
        );

    \I__5199\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28708\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28714\,
            I => \N__28703\
        );

    \I__5197\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28703\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__28708\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__28703\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__5194\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28691\
        );

    \I__5193\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28691\
        );

    \I__5192\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28688\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__28691\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__28688\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__28683\,
            I => \N__28680\
        );

    \I__5188\ : InMux
    port map (
            O => \N__28680\,
            I => \N__28677\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__28677\,
            I => \pid_alt.m35_e_2\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28669\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__28673\,
            I => \N__28664\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__28672\,
            I => \N__28661\
        );

    \I__5183\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28649\
        );

    \I__5182\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28649\
        );

    \I__5181\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28649\
        );

    \I__5180\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28649\
        );

    \I__5179\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28649\
        );

    \I__5178\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28646\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__28649\,
            I => \pid_alt.N_62_mux\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__28646\,
            I => \pid_alt.N_62_mux\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__28641\,
            I => \N__28638\
        );

    \I__5174\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28633\
        );

    \I__5173\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28630\
        );

    \I__5172\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28627\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28621\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28621\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__28627\,
            I => \N__28618\
        );

    \I__5168\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28615\
        );

    \I__5167\ : Span4Mux_v
    port map (
            O => \N__28621\,
            I => \N__28608\
        );

    \I__5166\ : Span4Mux_v
    port map (
            O => \N__28618\,
            I => \N__28608\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__28615\,
            I => \N__28608\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__5163\ : Odrv4
    port map (
            O => \N__28605\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__5161\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__28596\,
            I => \N__28591\
        );

    \I__5159\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28588\
        );

    \I__5158\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28585\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__28591\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__28588\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__28585\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__5154\ : InMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28570\
        );

    \I__5152\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28565\
        );

    \I__5151\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28565\
        );

    \I__5150\ : Odrv4
    port map (
            O => \N__28570\,
            I => \pid_alt.N_9_0\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__28565\,
            I => \pid_alt.N_9_0\
        );

    \I__5148\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__5146\ : Span4Mux_h
    port map (
            O => \N__28554\,
            I => \N__28549\
        );

    \I__5145\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28544\
        );

    \I__5144\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28544\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__28549\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__28544\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__5141\ : CascadeMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28530\
        );

    \I__5139\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28530\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__28530\,
            I => \uart_pc.N_144_1\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__5136\ : InMux
    port map (
            O => \N__28524\,
            I => \N__28517\
        );

    \I__5135\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28508\
        );

    \I__5134\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28508\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28521\,
            I => \N__28508\
        );

    \I__5132\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28508\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28502\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__28508\,
            I => \N__28502\
        );

    \I__5129\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28499\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__28502\,
            I => \N__28494\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__28499\,
            I => \N__28494\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__28494\,
            I => \N__28491\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__28491\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__5124\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28484\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28481\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28478\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__28481\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__5120\ : Odrv4
    port map (
            O => \N__28478\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__5119\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28470\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__28470\,
            I => \pid_alt.m21_e_8\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__28467\,
            I => \N__28463\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__28466\,
            I => \N__28460\
        );

    \I__5115\ : InMux
    port map (
            O => \N__28463\,
            I => \N__28457\
        );

    \I__5114\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28454\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__28457\,
            I => \N__28451\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__28454\,
            I => \N__28448\
        );

    \I__5111\ : Span4Mux_v
    port map (
            O => \N__28451\,
            I => \N__28443\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__28448\,
            I => \N__28443\
        );

    \I__5109\ : Span4Mux_h
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__28440\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__5107\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__28431\,
            I => \pid_alt.m21_e_2\
        );

    \I__5104\ : CascadeMux
    port map (
            O => \N__28428\,
            I => \pid_alt.m21_e_10_cascade_\
        );

    \I__5103\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__28419\,
            I => \pid_alt.N_138\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28413\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__28413\,
            I => \N__28410\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__28410\,
            I => \pid_alt.m35_e_3\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__28407\,
            I => \pid_alt.N_62_mux_cascade_\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28392\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28392\
        );

    \I__5094\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28392\
        );

    \I__5093\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28392\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__28392\,
            I => \pid_alt.N_129\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28385\
        );

    \I__5090\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28382\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__28382\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__28379\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__28374\,
            I => \pid_alt.m21_e_0_cascade_\
        );

    \I__5085\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__28368\,
            I => \pid_alt.m21_e_9\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28365\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__28362\,
            I => \pid_alt.un1_reset_1_0_i_cascade_\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__5080\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__28350\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\
        );

    \I__5077\ : InMux
    port map (
            O => \N__28347\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28341\,
            I => \N__28335\
        );

    \I__5074\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28335\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__28335\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28332\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__28329\,
            I => \N__28326\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28320\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28320\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28320\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\
        );

    \I__5067\ : InMux
    port map (
            O => \N__28317\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__28314\,
            I => \N__28311\
        );

    \I__5065\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28305\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28305\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__28305\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\
        );

    \I__5062\ : InMux
    port map (
            O => \N__28302\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__5059\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28290\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28290\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\
        );

    \I__5057\ : InMux
    port map (
            O => \N__28287\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__28284\,
            I => \N__28281\
        );

    \I__5055\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28275\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28275\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__28275\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\
        );

    \I__5052\ : InMux
    port map (
            O => \N__28272\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28260\
        );

    \I__5049\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28260\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__28260\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28257\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28250\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28247\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__28250\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28247\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__28242\,
            I => \N__28239\
        );

    \I__5041\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__28236\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__5039\ : InMux
    port map (
            O => \N__28233\,
            I => \bfn_12_17_0_\
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28221\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28221\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__28221\,
            I => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28218\,
            I => \scaler_3.un2_source_data_0_cry_2\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28206\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28206\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__28206\,
            I => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28203\,
            I => \scaler_3.un2_source_data_0_cry_3\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28191\
        );

    \I__5026\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28191\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__28191\,
            I => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\
        );

    \I__5024\ : InMux
    port map (
            O => \N__28188\,
            I => \scaler_3.un2_source_data_0_cry_4\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28176\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28176\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__28176\,
            I => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28173\,
            I => \scaler_3.un2_source_data_0_cry_5\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28161\
        );

    \I__5016\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28161\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__28161\,
            I => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28158\,
            I => \scaler_3.un2_source_data_0_cry_6\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__5012\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28146\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28146\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28146\,
            I => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28143\,
            I => \scaler_3.un2_source_data_0_cry_7\
        );

    \I__5008\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28136\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28133\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28136\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28133\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__28128\,
            I => \N__28125\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__28122\,
            I => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28119\,
            I => \bfn_12_15_0_\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28116\,
            I => \scaler_3.un2_source_data_0_cry_9\
        );

    \I__4999\ : InMux
    port map (
            O => \N__28113\,
            I => \bfn_12_12_0_\
        );

    \I__4998\ : InMux
    port map (
            O => \N__28110\,
            I => \scaler_2.un3_source_data_0_cry_8\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28104\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28104\,
            I => \N__28100\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28097\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__28100\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28097\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28088\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28085\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__28088\,
            I => \frame_decoder_CH2data_7\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__28085\,
            I => \frame_decoder_CH2data_7\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28077\,
            I => \scaler_2.N_1227_i_l_ofxZ0\
        );

    \I__4986\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28069\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__28073\,
            I => \N__28062\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__28072\,
            I => \N__28059\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28054\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28051\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28048\
        );

    \I__4980\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28044\
        );

    \I__4979\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28032\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28032\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28032\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28032\
        );

    \I__4975\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28032\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__28054\,
            I => \N__28027\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__28051\,
            I => \N__28027\
        );

    \I__4972\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28022\
        );

    \I__4971\ : InMux
    port map (
            O => \N__28047\,
            I => \N__28022\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__28044\,
            I => \N__28019\
        );

    \I__4969\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28016\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28011\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__28027\,
            I => \N__28011\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28008\
        );

    \I__4965\ : Span4Mux_v
    port map (
            O => \N__28019\,
            I => \N__28005\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__28002\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__28011\,
            I => \N__27999\
        );

    \I__4962\ : Span4Mux_v
    port map (
            O => \N__28008\,
            I => \N__27992\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__28005\,
            I => \N__27992\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__28002\,
            I => \N__27992\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__27999\,
            I => \pid_alt.pid_preregZ0Z_30\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__27992\,
            I => \pid_alt.pid_preregZ0Z_30\
        );

    \I__4957\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__4955\ : Span4Mux_h
    port map (
            O => \N__27981\,
            I => \N__27972\
        );

    \I__4954\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27969\
        );

    \I__4953\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27958\
        );

    \I__4952\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27958\
        );

    \I__4951\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27958\
        );

    \I__4950\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27958\
        );

    \I__4949\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27958\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__27972\,
            I => \pid_alt.N_106\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__27969\,
            I => \pid_alt.N_106\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__27958\,
            I => \pid_alt.N_106\
        );

    \I__4945\ : InMux
    port map (
            O => \N__27951\,
            I => \N__27948\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__27948\,
            I => \N__27944\
        );

    \I__4943\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27941\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__27944\,
            I => \N__27937\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27934\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27931\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__27937\,
            I => \N__27928\
        );

    \I__4938\ : Span4Mux_h
    port map (
            O => \N__27934\,
            I => \N__27923\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27923\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__27928\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__27923\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__4934\ : CEMux
    port map (
            O => \N__27918\,
            I => \N__27914\
        );

    \I__4933\ : CEMux
    port map (
            O => \N__27917\,
            I => \N__27909\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27906\
        );

    \I__4931\ : CEMux
    port map (
            O => \N__27913\,
            I => \N__27903\
        );

    \I__4930\ : CEMux
    port map (
            O => \N__27912\,
            I => \N__27900\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__27909\,
            I => \N__27897\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__27906\,
            I => \N__27894\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27891\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27888\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__27897\,
            I => \N__27885\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__27894\,
            I => \pid_alt.N_96_i_1\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__27891\,
            I => \pid_alt.N_96_i_1\
        );

    \I__4922\ : Odrv12
    port map (
            O => \N__27888\,
            I => \pid_alt.N_96_i_1\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__27885\,
            I => \pid_alt.N_96_i_1\
        );

    \I__4920\ : SRMux
    port map (
            O => \N__27876\,
            I => \N__27872\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27866\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__27869\,
            I => \N__27859\
        );

    \I__4916\ : Span4Mux_v
    port map (
            O => \N__27866\,
            I => \N__27856\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__27865\,
            I => \N__27853\
        );

    \I__4914\ : SRMux
    port map (
            O => \N__27864\,
            I => \N__27850\
        );

    \I__4913\ : SRMux
    port map (
            O => \N__27863\,
            I => \N__27847\
        );

    \I__4912\ : SRMux
    port map (
            O => \N__27862\,
            I => \N__27844\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__27859\,
            I => \N__27841\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__27856\,
            I => \N__27838\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__27853\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__27850\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__27847\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__27844\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__27841\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__27838\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N__27822\
        );

    \I__4902\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__4900\ : Odrv12
    port map (
            O => \N__27816\,
            I => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\
        );

    \I__4899\ : InMux
    port map (
            O => \N__27813\,
            I => \scaler_3.un2_source_data_0_cry_1\
        );

    \I__4898\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__27807\,
            I => \frame_decoder_CH2data_1\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__4895\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27798\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__27798\,
            I => \frame_decoder_OFF2data_1\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27795\,
            I => \scaler_2.un3_source_data_0_cry_0\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27792\,
            I => \N__27789\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__27789\,
            I => \frame_decoder_CH2data_2\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4889\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27780\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__27780\,
            I => \frame_decoder_OFF2data_2\
        );

    \I__4887\ : InMux
    port map (
            O => \N__27777\,
            I => \scaler_2.un3_source_data_0_cry_1\
        );

    \I__4886\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__27771\,
            I => \frame_decoder_CH2data_3\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__4883\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__27762\,
            I => \frame_decoder_OFF2data_3\
        );

    \I__4881\ : InMux
    port map (
            O => \N__27759\,
            I => \scaler_2.un3_source_data_0_cry_2\
        );

    \I__4880\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27753\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__27753\,
            I => \frame_decoder_CH2data_4\
        );

    \I__4878\ : CascadeMux
    port map (
            O => \N__27750\,
            I => \N__27747\
        );

    \I__4877\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27744\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__27744\,
            I => \frame_decoder_OFF2data_4\
        );

    \I__4875\ : InMux
    port map (
            O => \N__27741\,
            I => \scaler_2.un3_source_data_0_cry_3\
        );

    \I__4874\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__27735\,
            I => \frame_decoder_CH2data_5\
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__27732\,
            I => \N__27729\
        );

    \I__4871\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27726\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__27726\,
            I => \frame_decoder_OFF2data_5\
        );

    \I__4869\ : InMux
    port map (
            O => \N__27723\,
            I => \scaler_2.un3_source_data_0_cry_4\
        );

    \I__4868\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__27717\,
            I => \frame_decoder_CH2data_6\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__27714\,
            I => \N__27711\
        );

    \I__4865\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__27708\,
            I => \frame_decoder_OFF2data_6\
        );

    \I__4863\ : InMux
    port map (
            O => \N__27705\,
            I => \scaler_2.un3_source_data_0_cry_5\
        );

    \I__4862\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__27699\,
            I => \scaler_2.un3_source_data_0_axb_7\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27696\,
            I => \scaler_2.un3_source_data_0_cry_6\
        );

    \I__4859\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__27690\,
            I => \N__27687\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__27684\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__4855\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__27678\,
            I => \N__27674\
        );

    \I__4853\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27670\
        );

    \I__4852\ : Span4Mux_h
    port map (
            O => \N__27674\,
            I => \N__27666\
        );

    \I__4851\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27663\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__27670\,
            I => \N__27659\
        );

    \I__4849\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27656\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__27666\,
            I => \N__27646\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27646\
        );

    \I__4846\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27643\
        );

    \I__4845\ : Span4Mux_v
    port map (
            O => \N__27659\,
            I => \N__27640\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27637\
        );

    \I__4843\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27634\
        );

    \I__4842\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27631\
        );

    \I__4841\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27628\
        );

    \I__4840\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27625\
        );

    \I__4839\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27622\
        );

    \I__4838\ : Sp12to4
    port map (
            O => \N__27646\,
            I => \N__27617\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27617\
        );

    \I__4836\ : Sp12to4
    port map (
            O => \N__27640\,
            I => \N__27610\
        );

    \I__4835\ : Sp12to4
    port map (
            O => \N__27637\,
            I => \N__27603\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__27634\,
            I => \N__27603\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27631\,
            I => \N__27603\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__27628\,
            I => \N__27600\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__27625\,
            I => \N__27595\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27595\
        );

    \I__4829\ : Span12Mux_v
    port map (
            O => \N__27617\,
            I => \N__27592\
        );

    \I__4828\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27587\
        );

    \I__4827\ : InMux
    port map (
            O => \N__27615\,
            I => \N__27587\
        );

    \I__4826\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27582\
        );

    \I__4825\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27582\
        );

    \I__4824\ : Odrv12
    port map (
            O => \N__27610\,
            I => uart_pc_data_0
        );

    \I__4823\ : Odrv12
    port map (
            O => \N__27603\,
            I => uart_pc_data_0
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__27600\,
            I => uart_pc_data_0
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__27595\,
            I => uart_pc_data_0
        );

    \I__4820\ : Odrv12
    port map (
            O => \N__27592\,
            I => uart_pc_data_0
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__27587\,
            I => uart_pc_data_0
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__27582\,
            I => uart_pc_data_0
        );

    \I__4817\ : CEMux
    port map (
            O => \N__27567\,
            I => \N__27564\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27561\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__27561\,
            I => \N__27558\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__27558\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__27555\,
            I => \N__27548\
        );

    \I__4812\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27544\
        );

    \I__4811\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27539\
        );

    \I__4810\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27539\
        );

    \I__4809\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27536\
        );

    \I__4808\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27531\
        );

    \I__4807\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27531\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__27544\,
            I => \uart_pc.N_143\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__27539\,
            I => \uart_pc.N_143\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__27536\,
            I => \uart_pc.N_143\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__27531\,
            I => \uart_pc.N_143\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__27522\,
            I => \uart_pc.N_145_cascade_\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27516\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__27516\,
            I => \N__27513\
        );

    \I__4799\ : Span4Mux_h
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__27510\,
            I => \uart_drone.data_Auxce_0_0_4\
        );

    \I__4797\ : InMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__27498\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__27495\,
            I => \N__27491\
        );

    \I__4792\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27487\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27482\
        );

    \I__4790\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27482\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__27487\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__27482\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__4787\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27474\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__27471\,
            I => \uart_pc.N_126_li_cascade_\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__27468\,
            I => \N__27464\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__27467\,
            I => \N__27459\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27454\
        );

    \I__4781\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27454\
        );

    \I__4780\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27449\
        );

    \I__4779\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27449\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__27454\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__27449\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__4776\ : InMux
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__27441\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \uart_pc.timer_Count_0_sqmuxa_cascade_\
        );

    \I__4773\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__27432\,
            I => \pid_alt.error_i_acumm_preregZ0Z_15\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__27429\,
            I => \pid_alt.m7_e_4_cascade_\
        );

    \I__4770\ : CascadeMux
    port map (
            O => \N__27426\,
            I => \pid_alt.N_238_cascade_\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__27420\,
            I => \pid_alt.error_i_acumm_preregZ0Z_18\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__4766\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__27411\,
            I => \pid_alt.error_i_acumm_preregZ0Z_19\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__27405\,
            I => \pid_alt.error_i_acumm_preregZ0Z_14\
        );

    \I__4762\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__27399\,
            I => \pid_alt.error_i_acumm_preregZ0Z_17\
        );

    \I__4760\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27393\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__27393\,
            I => \pid_alt.error_i_acumm_preregZ0Z_20\
        );

    \I__4758\ : InMux
    port map (
            O => \N__27390\,
            I => \bfn_11_17_0_\
        );

    \I__4757\ : InMux
    port map (
            O => \N__27387\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__27381\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__4754\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27372\
        );

    \I__4753\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27372\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__27372\,
            I => \frame_decoder_CH4data_7\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__27369\,
            I => \N__27366\
        );

    \I__4750\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27360\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27360\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__27357\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__4746\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__27351\,
            I => \scaler_4.N_1251_i_l_ofxZ0\
        );

    \I__4744\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__4742\ : Span4Mux_h
    port map (
            O => \N__27342\,
            I => \N__27338\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27335\
        );

    \I__4740\ : Span4Mux_v
    port map (
            O => \N__27338\,
            I => \N__27330\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__27335\,
            I => \N__27330\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__27330\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__4737\ : CEMux
    port map (
            O => \N__27327\,
            I => \N__27324\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__27324\,
            I => \N__27321\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__27321\,
            I => \N__27318\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__27318\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__4733\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__27312\,
            I => \pid_alt.error_i_acumm_preregZ0Z_16\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27306\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__27306\,
            I => \frame_decoder_CH4data_1\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__27303\,
            I => \N__27300\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27297\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27297\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27294\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__27288\,
            I => \frame_decoder_CH4data_2\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__4722\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__4720\ : Odrv12
    port map (
            O => \N__27276\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27273\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__4718\ : InMux
    port map (
            O => \N__27270\,
            I => \N__27267\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__27267\,
            I => \frame_decoder_CH4data_3\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__27264\,
            I => \N__27261\
        );

    \I__4715\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__27258\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27255\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27249\,
            I => \N__27246\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__27240\,
            I => \frame_decoder_CH4data_4\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__27231\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27228\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__27222\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4697\ : Span4Mux_h
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__27204\,
            I => \frame_decoder_CH4data_5\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27201\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__27195\,
            I => \frame_decoder_CH4data_6\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__27186\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__4689\ : InMux
    port map (
            O => \N__27183\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27180\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27167\
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__27170\,
            I => \N__27163\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__27167\,
            I => \N__27160\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27157\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27154\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__27160\,
            I => \N__27149\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__27157\,
            I => \N__27149\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27154\,
            I => \N__27144\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__27149\,
            I => \N__27144\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__27144\,
            I => \pid_alt.pid_preregZ0Z_7\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__27141\,
            I => \N__27137\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27133\
        );

    \I__4673\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27130\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__27136\,
            I => \N__27127\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__27133\,
            I => \N__27124\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27130\,
            I => \N__27121\
        );

    \I__4669\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27118\
        );

    \I__4668\ : Span4Mux_h
    port map (
            O => \N__27124\,
            I => \N__27115\
        );

    \I__4667\ : Span4Mux_h
    port map (
            O => \N__27121\,
            I => \N__27110\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__27118\,
            I => \N__27110\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__27115\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__27110\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27101\
        );

    \I__4662\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27098\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27101\,
            I => \N__27094\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27091\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27088\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__27094\,
            I => \N__27081\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__27091\,
            I => \N__27081\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27081\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__27081\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27072\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__27069\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_4\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27063\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27063\,
            I => \N__27060\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__27060\,
            I => \N__27056\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27059\,
            I => \N__27053\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__27056\,
            I => \N__27050\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__27053\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__27050\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27036\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__27044\,
            I => \N__27032\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__27043\,
            I => \N__27029\
        );

    \I__4640\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27023\
        );

    \I__4639\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27017\
        );

    \I__4638\ : InMux
    port map (
            O => \N__27040\,
            I => \N__27014\
        );

    \I__4637\ : InMux
    port map (
            O => \N__27039\,
            I => \N__27011\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__27036\,
            I => \N__27005\
        );

    \I__4635\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27000\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27000\
        );

    \I__4633\ : InMux
    port map (
            O => \N__27029\,
            I => \N__26993\
        );

    \I__4632\ : InMux
    port map (
            O => \N__27028\,
            I => \N__26993\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27027\,
            I => \N__26990\
        );

    \I__4630\ : CascadeMux
    port map (
            O => \N__27026\,
            I => \N__26986\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__26983\
        );

    \I__4628\ : InMux
    port map (
            O => \N__27022\,
            I => \N__26976\
        );

    \I__4627\ : InMux
    port map (
            O => \N__27021\,
            I => \N__26976\
        );

    \I__4626\ : InMux
    port map (
            O => \N__27020\,
            I => \N__26976\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__27017\,
            I => \N__26973\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__27014\,
            I => \N__26969\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__27011\,
            I => \N__26966\
        );

    \I__4622\ : InMux
    port map (
            O => \N__27010\,
            I => \N__26959\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27009\,
            I => \N__26959\
        );

    \I__4620\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26959\
        );

    \I__4619\ : Span4Mux_v
    port map (
            O => \N__27005\,
            I => \N__26954\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26954\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \N__26950\
        );

    \I__4616\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26947\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26942\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26942\
        );

    \I__4613\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26937\
        );

    \I__4612\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26937\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__26983\,
            I => \N__26934\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__26976\,
            I => \N__26929\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__26973\,
            I => \N__26929\
        );

    \I__4608\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26926\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__26969\,
            I => \N__26917\
        );

    \I__4606\ : Span4Mux_v
    port map (
            O => \N__26966\,
            I => \N__26917\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__26959\,
            I => \N__26917\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__26954\,
            I => \N__26917\
        );

    \I__4603\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26912\
        );

    \I__4602\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26912\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__26947\,
            I => uart_pc_data_rdy
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__26942\,
            I => uart_pc_data_rdy
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__26937\,
            I => uart_pc_data_rdy
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__26934\,
            I => uart_pc_data_rdy
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__26929\,
            I => uart_pc_data_rdy
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__26926\,
            I => uart_pc_data_rdy
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__26917\,
            I => uart_pc_data_rdy
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__26912\,
            I => uart_pc_data_rdy
        );

    \I__4593\ : InMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__26889\,
            I => \frame_decoder_CH3data_2\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__4589\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__26880\,
            I => \frame_decoder_OFF3data_2\
        );

    \I__4587\ : InMux
    port map (
            O => \N__26877\,
            I => \scaler_3.un3_source_data_0_cry_1\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__26868\,
            I => \frame_decoder_CH3data_3\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__4582\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__26859\,
            I => \frame_decoder_OFF3data_3\
        );

    \I__4580\ : InMux
    port map (
            O => \N__26856\,
            I => \scaler_3.un3_source_data_0_cry_2\
        );

    \I__4579\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26850\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__4577\ : Span4Mux_h
    port map (
            O => \N__26847\,
            I => \N__26844\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__26844\,
            I => \frame_decoder_CH3data_4\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__4574\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__26835\,
            I => \frame_decoder_OFF3data_4\
        );

    \I__4572\ : InMux
    port map (
            O => \N__26832\,
            I => \scaler_3.un3_source_data_0_cry_3\
        );

    \I__4571\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__4569\ : Span4Mux_h
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__26820\,
            I => \frame_decoder_CH3data_5\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__26817\,
            I => \N__26814\
        );

    \I__4566\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__26808\,
            I => \frame_decoder_OFF3data_5\
        );

    \I__4563\ : InMux
    port map (
            O => \N__26805\,
            I => \scaler_3.un3_source_data_0_cry_4\
        );

    \I__4562\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__26793\,
            I => \frame_decoder_CH3data_6\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__4557\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26784\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__26784\,
            I => \frame_decoder_OFF3data_6\
        );

    \I__4555\ : InMux
    port map (
            O => \N__26781\,
            I => \scaler_3.un3_source_data_0_cry_5\
        );

    \I__4554\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__26772\,
            I => \scaler_3.un3_source_data_0_axb_7\
        );

    \I__4551\ : InMux
    port map (
            O => \N__26769\,
            I => \scaler_3.un3_source_data_0_cry_6\
        );

    \I__4550\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__26760\,
            I => \scaler_3.N_1239_i_l_ofxZ0\
        );

    \I__4547\ : InMux
    port map (
            O => \N__26757\,
            I => \bfn_11_14_0_\
        );

    \I__4546\ : InMux
    port map (
            O => \N__26754\,
            I => \scaler_3.un3_source_data_0_cry_8\
        );

    \I__4545\ : CEMux
    port map (
            O => \N__26751\,
            I => \N__26748\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__4543\ : Sp12to4
    port map (
            O => \N__26745\,
            I => \N__26741\
        );

    \I__4542\ : CEMux
    port map (
            O => \N__26744\,
            I => \N__26738\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__26741\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__26738\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__4539\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__26730\,
            I => \frame_decoder_OFF3data_1\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__4536\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__4534\ : Span4Mux_v
    port map (
            O => \N__26718\,
            I => \N__26715\
        );

    \I__4533\ : Odrv4
    port map (
            O => \N__26715\,
            I => \frame_decoder_CH3data_1\
        );

    \I__4532\ : InMux
    port map (
            O => \N__26712\,
            I => \scaler_3.un3_source_data_0_cry_0\
        );

    \I__4531\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26705\
        );

    \I__4530\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26702\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__26705\,
            I => \N__26699\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26696\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__26699\,
            I => \N__26693\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__26696\,
            I => \N__26690\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__26693\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__26690\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__4523\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26681\
        );

    \I__4522\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26678\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__26681\,
            I => \N__26675\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__26678\,
            I => \frame_decoder_CH3data_7\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__26675\,
            I => \frame_decoder_CH3data_7\
        );

    \I__4518\ : CEMux
    port map (
            O => \N__26670\,
            I => \N__26667\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__26661\,
            I => \N__26658\
        );

    \I__4514\ : Odrv4
    port map (
            O => \N__26658\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__26655\,
            I => \N__26651\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26646\
        );

    \I__4511\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26639\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26639\
        );

    \I__4509\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26639\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__26646\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__26639\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__4506\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26629\
        );

    \I__4505\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26624\
        );

    \I__4504\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26624\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__26629\,
            I => \Commands_frame_decoder.countZ0Z_1\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__26624\,
            I => \Commands_frame_decoder.countZ0Z_1\
        );

    \I__4501\ : SRMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__4498\ : Sp12to4
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__4497\ : Odrv12
    port map (
            O => \N__26607\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__26604\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\
        );

    \I__4495\ : CEMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__26589\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__4490\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26581\
        );

    \I__4489\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26578\
        );

    \I__4488\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26575\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26569\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26569\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__26575\,
            I => \N__26566\
        );

    \I__4484\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26563\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__26569\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4482\ : Odrv12
    port map (
            O => \N__26566\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__26563\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4480\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__26553\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__4478\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__26547\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__4476\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__26541\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__26538\,
            I => \N__26532\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26529\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26526\
        );

    \I__4471\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26521\
        );

    \I__4470\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26521\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__26529\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__26526\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__26521\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26507\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26504\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26507\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__26504\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__4461\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26493\
        );

    \I__4460\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26493\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__26493\,
            I => \N__26490\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__26490\,
            I => \Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__26487\,
            I => \Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26477\
        );

    \I__4455\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26477\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26473\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26470\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26467\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__26473\,
            I => \N__26459\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__26470\,
            I => \N__26459\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__26467\,
            I => \N__26459\
        );

    \I__4448\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26456\
        );

    \I__4447\ : Span4Mux_h
    port map (
            O => \N__26459\,
            I => \N__26453\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__26456\,
            I => \Commands_frame_decoder.stateZ0Z_12\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__26453\,
            I => \Commands_frame_decoder.stateZ0Z_12\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26445\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26441\
        );

    \I__4442\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26438\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__26441\,
            I => \N__26433\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26433\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__26433\,
            I => \Commands_frame_decoder.N_330\
        );

    \I__4438\ : InMux
    port map (
            O => \N__26430\,
            I => \N__26427\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__26427\,
            I => \N__26424\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__26424\,
            I => \Commands_frame_decoder.state_ns_i_a4_2_0_0\
        );

    \I__4435\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__26418\,
            I => \uart_pc_sync.aux_3__0_Z0Z_0\
        );

    \I__4433\ : InMux
    port map (
            O => \N__26415\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__4432\ : InMux
    port map (
            O => \N__26412\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26409\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26403\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26403\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__4428\ : CEMux
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__26397\,
            I => \N__26393\
        );

    \I__4426\ : CEMux
    port map (
            O => \N__26396\,
            I => \N__26390\
        );

    \I__4425\ : Span4Mux_h
    port map (
            O => \N__26393\,
            I => \N__26387\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26384\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__26387\,
            I => \N__26378\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__26384\,
            I => \N__26378\
        );

    \I__4421\ : CEMux
    port map (
            O => \N__26383\,
            I => \N__26375\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__26378\,
            I => \N__26372\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26369\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__26372\,
            I => \N__26364\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__26369\,
            I => \N__26364\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__26364\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__4415\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26355\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__26355\,
            I => \Commands_frame_decoder.source_CH1data8lt7_0\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26349\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__26349\,
            I => \N__26346\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__26346\,
            I => \N__26342\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26339\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__26342\,
            I => \N__26336\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26333\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__26336\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__26333\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26324\
        );

    \I__4403\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26321\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__26324\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__26321\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26312\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__26315\,
            I => \N__26309\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26306\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26303\
        );

    \I__4396\ : Span4Mux_v
    port map (
            O => \N__26306\,
            I => \N__26300\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__26303\,
            I => \N__26297\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__26300\,
            I => \N__26294\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__26297\,
            I => \N__26291\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__26294\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__26291\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26283\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__26283\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24\
        );

    \I__4388\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26276\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26273\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26270\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__26273\,
            I => \N__26267\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__26270\,
            I => \N__26264\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__26267\,
            I => \N__26261\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__26264\,
            I => \N__26258\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__26261\,
            I => \N__26255\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__26258\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__26255\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__26244\,
            I => \N__26240\
        );

    \I__4375\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26237\
        );

    \I__4374\ : Span4Mux_h
    port map (
            O => \N__26240\,
            I => \N__26234\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__26234\,
            I => \N__26228\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__26231\,
            I => \N__26225\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__26228\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__26225\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26217\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26217\,
            I => \N__26214\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26211\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__26211\,
            I => \N__26208\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__26208\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23\
        );

    \I__4363\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26202\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__26202\,
            I => \N__26197\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26194\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26191\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__26197\,
            I => \N__26187\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26194\,
            I => \N__26184\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__26191\,
            I => \N__26181\
        );

    \I__4356\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26178\
        );

    \I__4355\ : Span4Mux_v
    port map (
            O => \N__26187\,
            I => \N__26175\
        );

    \I__4354\ : Span12Mux_v
    port map (
            O => \N__26184\,
            I => \N__26172\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__26181\,
            I => \N__26169\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26166\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__26175\,
            I => uart_drone_data_3
        );

    \I__4350\ : Odrv12
    port map (
            O => \N__26172\,
            I => uart_drone_data_3
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__26169\,
            I => uart_drone_data_3
        );

    \I__4348\ : Odrv4
    port map (
            O => \N__26166\,
            I => uart_drone_data_3
        );

    \I__4347\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26154\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26151\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__26151\,
            I => \dron_frame_decoder_1.drone_altitude_11\
        );

    \I__4344\ : CEMux
    port map (
            O => \N__26148\,
            I => \N__26144\
        );

    \I__4343\ : CEMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26135\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__26138\,
            I => \N__26132\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__26135\,
            I => \N__26129\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__26129\,
            I => \N__26123\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__26126\,
            I => \dron_frame_decoder_1.N_384_0\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__26123\,
            I => \dron_frame_decoder_1.N_384_0\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__4333\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26111\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26108\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26102\
        );

    \I__4329\ : Span12Mux_v
    port map (
            O => \N__26105\,
            I => \N__26099\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__26102\,
            I => \N__26096\
        );

    \I__4327\ : Odrv12
    port map (
            O => \N__26099\,
            I => \pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__26096\,
            I => \pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__26091\,
            I => \N__26088\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__4322\ : Span4Mux_h
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__26079\,
            I => \pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3\
        );

    \I__4320\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26070\
        );

    \I__4319\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26070\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__26064\,
            I => \N__26061\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__26061\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26052\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26052\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26052\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__26049\,
            I => \N__26045\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26042\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26039\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26036\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__26039\,
            I => \N__26033\
        );

    \I__4306\ : Span4Mux_h
    port map (
            O => \N__26036\,
            I => \N__26030\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__26033\,
            I => \N__26027\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__26030\,
            I => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__26027\,
            I => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__26022\,
            I => \N__26019\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26013\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26013\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__26013\,
            I => \pid_alt.error_d_reg_prevZ0Z_4\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26010\,
            I => \N__26007\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26007\,
            I => \N__26002\
        );

    \I__4296\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25997\
        );

    \I__4295\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25997\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__26002\,
            I => \N__25992\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25992\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__25992\,
            I => \N__25989\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__25989\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__4290\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25982\
        );

    \I__4289\ : InMux
    port map (
            O => \N__25985\,
            I => \N__25979\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__25982\,
            I => \N__25976\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25972\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25969\
        );

    \I__4285\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25966\
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__25972\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__25969\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__25966\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__4281\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25955\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__25958\,
            I => \N__25952\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__25955\,
            I => \N__25948\
        );

    \I__4278\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25945\
        );

    \I__4277\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25942\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__25948\,
            I => \N__25937\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__25945\,
            I => \N__25937\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__25942\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__25937\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__4272\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25929\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25924\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25919\
        );

    \I__4269\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25919\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__25924\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__25919\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__4266\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25911\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__25911\,
            I => \N__25908\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__25908\,
            I => \N__25901\
        );

    \I__4263\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25892\
        );

    \I__4262\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25892\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25892\
        );

    \I__4260\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25892\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__25901\,
            I => \pid_alt.N_91_1\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__25892\,
            I => \pid_alt.N_91_1\
        );

    \I__4257\ : InMux
    port map (
            O => \N__25887\,
            I => \N__25883\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25880\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__25883\,
            I => \N__25876\
        );

    \I__4254\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25871\
        );

    \I__4253\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25871\
        );

    \I__4252\ : Odrv12
    port map (
            O => \N__25876\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__25871\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__4250\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25863\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__25863\,
            I => \N__25859\
        );

    \I__4248\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25856\
        );

    \I__4247\ : Span4Mux_v
    port map (
            O => \N__25859\,
            I => \N__25853\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__25856\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__25853\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\
        );

    \I__4244\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25844\
        );

    \I__4243\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25841\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25836\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25836\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__25836\,
            I => \N__25833\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__4237\ : Odrv4
    port map (
            O => \N__25827\,
            I => \pid_alt.error_p_regZ0Z_5\
        );

    \I__4236\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25820\
        );

    \I__4235\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25817\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__25820\,
            I => \N__25812\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__25817\,
            I => \N__25812\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__25812\,
            I => \pid_alt.error_d_reg_prevZ0Z_5\
        );

    \I__4231\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25803\
        );

    \I__4230\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25803\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__25803\,
            I => \N__25799\
        );

    \I__4228\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25796\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__25799\,
            I => \N__25793\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25790\
        );

    \I__4225\ : Sp12to4
    port map (
            O => \N__25793\,
            I => \N__25785\
        );

    \I__4224\ : Span12Mux_v
    port map (
            O => \N__25790\,
            I => \N__25785\
        );

    \I__4223\ : Odrv12
    port map (
            O => \N__25785\,
            I => \pid_alt.error_d_regZ0Z_5\
        );

    \I__4222\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25776\
        );

    \I__4221\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25776\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__25776\,
            I => \N__25773\
        );

    \I__4219\ : Odrv4
    port map (
            O => \N__25773\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__25770\,
            I => \N__25766\
        );

    \I__4217\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25763\
        );

    \I__4216\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25760\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__25763\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__25760\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__25755\,
            I => \N__25751\
        );

    \I__4212\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25748\
        );

    \I__4211\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25745\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__25748\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__25745\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__4208\ : CEMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__25734\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\
        );

    \I__4204\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25724\
        );

    \I__4203\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25721\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__25724\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25721\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__4200\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25713\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__25710\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__25707\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \N__25700\
        );

    \I__4195\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25697\
        );

    \I__4194\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25694\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__25697\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__25694\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__25689\,
            I => \N__25685\
        );

    \I__4190\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25682\
        );

    \I__4189\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25679\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__25682\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__25679\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__25674\,
            I => \N__25670\
        );

    \I__4185\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__4184\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25664\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__25667\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__25664\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__25659\,
            I => \N__25655\
        );

    \I__4180\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25652\
        );

    \I__4179\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25649\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__25652\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__25649\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__4176\ : InMux
    port map (
            O => \N__25644\,
            I => \N__25640\
        );

    \I__4175\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__25640\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__25637\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__25632\,
            I => \N__25628\
        );

    \I__4171\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25625\
        );

    \I__4170\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25622\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__25625\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__25622\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__4167\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25612\
        );

    \I__4166\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25609\
        );

    \I__4165\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25606\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__25612\,
            I => \Commands_frame_decoder.N_320_0\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__25609\,
            I => \Commands_frame_decoder.N_320_0\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__25606\,
            I => \Commands_frame_decoder.N_320_0\
        );

    \I__4161\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__25596\,
            I => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__25593\,
            I => \Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_\
        );

    \I__4158\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__25587\,
            I => \Commands_frame_decoder.state_ns_0_a4_0_3_2\
        );

    \I__4156\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25578\
        );

    \I__4155\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25573\
        );

    \I__4154\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25573\
        );

    \I__4153\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25570\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__25578\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__25573\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__25570\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__4149\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25556\
        );

    \I__4148\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25556\
        );

    \I__4147\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25553\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__25556\,
            I => \Commands_frame_decoder.N_364\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__25553\,
            I => \Commands_frame_decoder.N_364\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__25548\,
            I => \Commands_frame_decoder.N_360_cascade_\
        );

    \I__4143\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25542\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__25542\,
            I => \Commands_frame_decoder.N_359\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__4140\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__25533\,
            I => \Commands_frame_decoder.state_ns_i_0_0\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__25530\,
            I => \N__25525\
        );

    \I__4137\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25519\
        );

    \I__4136\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25519\
        );

    \I__4135\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25516\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25513\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25519\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__25516\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25513\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__25497\,
            I => \N__25494\
        );

    \I__4126\ : Sp12to4
    port map (
            O => \N__25494\,
            I => \N__25490\
        );

    \I__4125\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__4124\ : Span12Mux_s10_h
    port map (
            O => \N__25490\,
            I => \N__25484\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__25487\,
            I => alt_kp_4
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__25484\,
            I => alt_kp_4
        );

    \I__4121\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25475\
        );

    \I__4120\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25472\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__25475\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__25472\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__4117\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__25464\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__4115\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__25458\,
            I => \uart_pc_sync.aux_2__0_Z0Z_0\
        );

    \I__4113\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__25449\,
            I => \uart_pc_sync.aux_0__0_Z0Z_0\
        );

    \I__4110\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__25443\,
            I => \uart_pc_sync.aux_1__0_Z0Z_0\
        );

    \I__4108\ : SRMux
    port map (
            O => \N__25440\,
            I => \N__25436\
        );

    \I__4107\ : SRMux
    port map (
            O => \N__25439\,
            I => \N__25433\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__25436\,
            I => \Commands_frame_decoder.un1_state53_iZ0\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25433\,
            I => \Commands_frame_decoder.un1_state53_iZ0\
        );

    \I__4104\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25422\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25417\
        );

    \I__4102\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25417\
        );

    \I__4101\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25414\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__25422\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__25417\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__25414\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4097\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25401\
        );

    \I__4096\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25398\
        );

    \I__4095\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25395\
        );

    \I__4094\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25392\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__25401\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__25398\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25395\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__25392\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25377\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25374\
        );

    \I__4087\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25371\
        );

    \I__4086\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25368\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__25377\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__25374\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__25371\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__25368\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25355\
        );

    \I__4080\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25351\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__25355\,
            I => \N__25348\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25343\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25340\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__25348\,
            I => \N__25337\
        );

    \I__4075\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25334\
        );

    \I__4074\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25331\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__25343\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__25340\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__25337\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__25334\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25331\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__25320\,
            I => \Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25312\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25309\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25304\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__25312\,
            I => \N__25299\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__25309\,
            I => \N__25299\
        );

    \I__4062\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25296\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25293\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25304\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__25299\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25296\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__25293\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__25278\,
            I => \Commands_frame_decoder.state_0_sqmuxacf0\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__25275\,
            I => \N__25272\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25263\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25256\
        );

    \I__4049\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25256\
        );

    \I__4048\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25256\
        );

    \I__4047\ : Odrv12
    port map (
            O => \N__25263\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__25256\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__4045\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25248\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__25245\,
            I => \Commands_frame_decoder.count_1_sqmuxa\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25239\,
            I => \N__25235\
        );

    \I__4040\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__25235\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__25232\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__4036\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__25221\,
            I => \Commands_frame_decoder.state_ns_0_a4_0_1_1\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25213\
        );

    \I__4033\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25210\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25206\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__25213\,
            I => \N__25201\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25201\
        );

    \I__4029\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25198\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__25206\,
            I => \N__25195\
        );

    \I__4027\ : Span12Mux_v
    port map (
            O => \N__25201\,
            I => \N__25192\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__25198\,
            I => \N__25187\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__25195\,
            I => \N__25187\
        );

    \I__4024\ : Odrv12
    port map (
            O => \N__25192\,
            I => uart_drone_data_4
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__25187\,
            I => uart_drone_data_4
        );

    \I__4022\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25179\,
            I => drone_altitude_12
        );

    \I__4020\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25171\
        );

    \I__4019\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25168\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25174\,
            I => \N__25165\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__25171\,
            I => \N__25160\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25168\,
            I => \N__25160\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__25165\,
            I => \N__25157\
        );

    \I__4014\ : Span12Mux_v
    port map (
            O => \N__25160\,
            I => \N__25154\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__25157\,
            I => \N__25151\
        );

    \I__4012\ : Odrv12
    port map (
            O => \N__25154\,
            I => uart_drone_data_5
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__25151\,
            I => uart_drone_data_5
        );

    \I__4010\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25143\,
            I => drone_altitude_13
        );

    \I__4008\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25134\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25131\
        );

    \I__4006\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25128\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \N__25125\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__25134\,
            I => \N__25120\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__25131\,
            I => \N__25120\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__25128\,
            I => \N__25117\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25114\
        );

    \I__4000\ : Span12Mux_v
    port map (
            O => \N__25120\,
            I => \N__25111\
        );

    \I__3999\ : Span4Mux_h
    port map (
            O => \N__25117\,
            I => \N__25108\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__25114\,
            I => \N__25105\
        );

    \I__3997\ : Odrv12
    port map (
            O => \N__25111\,
            I => uart_drone_data_6
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__25108\,
            I => uart_drone_data_6
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__25105\,
            I => uart_drone_data_6
        );

    \I__3994\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25095\,
            I => drone_altitude_14
        );

    \I__3992\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25087\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25084\
        );

    \I__3990\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25081\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__25087\,
            I => \N__25076\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__25084\,
            I => \N__25076\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25073\
        );

    \I__3986\ : Span12Mux_v
    port map (
            O => \N__25076\,
            I => \N__25070\
        );

    \I__3985\ : Span4Mux_h
    port map (
            O => \N__25073\,
            I => \N__25067\
        );

    \I__3984\ : Odrv12
    port map (
            O => \N__25070\,
            I => uart_drone_data_7
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__25067\,
            I => uart_drone_data_7
        );

    \I__3982\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25059\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__25056\,
            I => drone_altitude_15
        );

    \I__3979\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25050\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__25050\,
            I => \N__25046\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25049\,
            I => \N__25043\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__25046\,
            I => \N__25037\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__25043\,
            I => \N__25037\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25034\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__25037\,
            I => \N__25031\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__25034\,
            I => \N__25028\
        );

    \I__3971\ : Span4Mux_v
    port map (
            O => \N__25031\,
            I => \N__25023\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__25028\,
            I => \N__25023\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__25023\,
            I => uart_drone_data_0
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__25014\,
            I => \dron_frame_decoder_1.drone_altitude_8\
        );

    \I__3965\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25006\
        );

    \I__3964\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25003\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25009\,
            I => \N__24999\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24994\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__24994\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24991\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24988\
        );

    \I__3958\ : Span12Mux_v
    port map (
            O => \N__24994\,
            I => \N__24985\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24982\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__24988\,
            I => \N__24979\
        );

    \I__3955\ : Odrv12
    port map (
            O => \N__24985\,
            I => uart_drone_data_1
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__24982\,
            I => uart_drone_data_1
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__24979\,
            I => uart_drone_data_1
        );

    \I__3952\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__24969\,
            I => \dron_frame_decoder_1.drone_altitude_9\
        );

    \I__3950\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__24963\,
            I => \N__24958\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N__24954\
        );

    \I__3947\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24951\
        );

    \I__3946\ : Span4Mux_s3_v
    port map (
            O => \N__24958\,
            I => \N__24947\
        );

    \I__3945\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24942\
        );

    \I__3944\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24942\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__24951\,
            I => \N__24939\
        );

    \I__3942\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24936\
        );

    \I__3941\ : Span4Mux_v
    port map (
            O => \N__24947\,
            I => \N__24933\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__24942\,
            I => \N__24930\
        );

    \I__3939\ : Span4Mux_v
    port map (
            O => \N__24939\,
            I => \N__24927\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24922\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__24933\,
            I => \N__24922\
        );

    \I__3936\ : Span4Mux_h
    port map (
            O => \N__24930\,
            I => \N__24919\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__24927\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__24922\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__24919\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__3932\ : IoInMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__3930\ : Span4Mux_s2_v
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__24903\,
            I => \pid_alt.state_0_0\
        );

    \I__3928\ : CEMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__24897\,
            I => \N__24894\
        );

    \I__3926\ : Span12Mux_h
    port map (
            O => \N__24894\,
            I => \N__24891\
        );

    \I__3925\ : Odrv12
    port map (
            O => \N__24891\,
            I => \dron_frame_decoder_1.N_392_0\
        );

    \I__3924\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24885\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__24885\,
            I => \N__24882\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__24882\,
            I => \N__24878\
        );

    \I__3921\ : InMux
    port map (
            O => \N__24881\,
            I => \N__24875\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__24878\,
            I => \N__24870\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24870\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__24870\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__3917\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24850\
        );

    \I__3915\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24845\
        );

    \I__3914\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24845\
        );

    \I__3913\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24838\
        );

    \I__3912\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24838\
        );

    \I__3911\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24838\
        );

    \I__3910\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24825\
        );

    \I__3909\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24825\
        );

    \I__3908\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24825\
        );

    \I__3907\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24825\
        );

    \I__3906\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24825\
        );

    \I__3905\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24825\
        );

    \I__3904\ : Odrv12
    port map (
            O => \N__24850\,
            I => \Commands_frame_decoder.N_358\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__24845\,
            I => \Commands_frame_decoder.N_358\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__24838\,
            I => \Commands_frame_decoder.N_358\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__24825\,
            I => \Commands_frame_decoder.N_358\
        );

    \I__3900\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24813\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__24813\,
            I => \dron_frame_decoder_1.drone_altitude_4\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__24810\,
            I => \N__24807\
        );

    \I__3897\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__24801\,
            I => drone_altitude_i_4
        );

    \I__3894\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__24795\,
            I => \dron_frame_decoder_1.drone_altitude_5\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__3891\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__24783\,
            I => drone_altitude_i_5
        );

    \I__3888\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__24777\,
            I => \dron_frame_decoder_1.drone_altitude_6\
        );

    \I__3886\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24771\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__24771\,
            I => \N__24768\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__24768\,
            I => drone_altitude_i_6
        );

    \I__3883\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24762\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__24762\,
            I => \dron_frame_decoder_1.drone_altitude_7\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__3880\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__24750\,
            I => drone_altitude_i_7
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__3876\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__24738\,
            I => \N__24735\
        );

    \I__3873\ : Odrv4
    port map (
            O => \N__24735\,
            I => drone_altitude_i_8
        );

    \I__3872\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24727\
        );

    \I__3871\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24724\
        );

    \I__3870\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24721\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__24727\,
            I => \N__24718\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__24724\,
            I => \N__24713\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24713\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__24718\,
            I => \N__24710\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__24713\,
            I => uart_drone_data_2
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__24710\,
            I => uart_drone_data_2
        );

    \I__3863\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__24702\,
            I => \dron_frame_decoder_1.drone_altitude_10\
        );

    \I__3861\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24693\
        );

    \I__3860\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24693\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__24693\,
            I => \pid_alt.error_d_reg_prevZ0Z_24\
        );

    \I__3858\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24681\
        );

    \I__3857\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24681\
        );

    \I__3856\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24681\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__3854\ : Span4Mux_v
    port map (
            O => \N__24678\,
            I => \N__24675\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__3852\ : Span4Mux_h
    port map (
            O => \N__24672\,
            I => \N__24669\
        );

    \I__3851\ : Span4Mux_v
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__24666\,
            I => \pid_alt.error_d_regZ0Z_24\
        );

    \I__3849\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24654\
        );

    \I__3848\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24651\
        );

    \I__3847\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24648\
        );

    \I__3846\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24643\
        );

    \I__3845\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24643\
        );

    \I__3844\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24638\
        );

    \I__3843\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24638\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24623\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24623\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24623\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__24643\,
            I => \N__24623\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__24638\,
            I => \N__24623\
        );

    \I__3837\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24615\
        );

    \I__3836\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24615\
        );

    \I__3835\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24615\
        );

    \I__3834\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24609\
        );

    \I__3833\ : Span4Mux_v
    port map (
            O => \N__24623\,
            I => \N__24605\
        );

    \I__3832\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24602\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24599\
        );

    \I__3830\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24596\
        );

    \I__3829\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24591\
        );

    \I__3828\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24591\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__24609\,
            I => \N__24588\
        );

    \I__3826\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24585\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__24605\,
            I => \N__24580\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__24602\,
            I => \N__24580\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__24599\,
            I => \N__24573\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24573\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24573\
        );

    \I__3820\ : Span4Mux_h
    port map (
            O => \N__24588\,
            I => \N__24568\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24568\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__24580\,
            I => \N__24565\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__24573\,
            I => \N__24560\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__24568\,
            I => \N__24560\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__24565\,
            I => \N__24557\
        );

    \I__3814\ : Span4Mux_v
    port map (
            O => \N__24560\,
            I => \N__24554\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__24557\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__24554\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3811\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24543\
        );

    \I__3810\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24543\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__24543\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24\
        );

    \I__3808\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24536\
        );

    \I__3807\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24533\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24530\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__24533\,
            I => \N__24527\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__24530\,
            I => \N__24524\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__24527\,
            I => \N__24521\
        );

    \I__3802\ : Span4Mux_h
    port map (
            O => \N__24524\,
            I => \N__24516\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__24521\,
            I => \N__24516\
        );

    \I__3800\ : Span4Mux_h
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__24513\,
            I => \pid_alt.error_p_regZ0Z_6\
        );

    \I__3798\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24506\
        );

    \I__3797\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24503\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24500\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24503\,
            I => \pid_alt.error_d_reg_prevZ0Z_6\
        );

    \I__3794\ : Odrv12
    port map (
            O => \N__24500\,
            I => \pid_alt.error_d_reg_prevZ0Z_6\
        );

    \I__3793\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24491\
        );

    \I__3792\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24488\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24482\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__24488\,
            I => \N__24482\
        );

    \I__3789\ : InMux
    port map (
            O => \N__24487\,
            I => \N__24479\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__24482\,
            I => \N__24474\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24474\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__24474\,
            I => \N__24471\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__24468\,
            I => \N__24465\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__24465\,
            I => \pid_alt.error_d_regZ0Z_6\
        );

    \I__3782\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24455\
        );

    \I__3780\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24452\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__24455\,
            I => \N__24448\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__24452\,
            I => \N__24445\
        );

    \I__3777\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24442\
        );

    \I__3776\ : Span4Mux_h
    port map (
            O => \N__24448\,
            I => \N__24439\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__24445\,
            I => \N__24436\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24442\,
            I => \N__24433\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__24439\,
            I => \N__24430\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__24436\,
            I => \N__24425\
        );

    \I__3771\ : Span4Mux_v
    port map (
            O => \N__24433\,
            I => \N__24425\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__24430\,
            I => \N__24422\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__24425\,
            I => \N__24419\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__24422\,
            I => \N__24415\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__24419\,
            I => \N__24412\
        );

    \I__3766\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24409\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__24415\,
            I => drone_altitude_0
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__24412\,
            I => drone_altitude_0
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__24409\,
            I => drone_altitude_0
        );

    \I__3762\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24399\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__24399\,
            I => drone_altitude_1
        );

    \I__3760\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__24393\,
            I => drone_altitude_2
        );

    \I__3758\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__24387\,
            I => drone_altitude_3
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3755\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__3753\ : Span4Mux_h
    port map (
            O => \N__24375\,
            I => \N__24372\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__24372\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25\
        );

    \I__3751\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24363\
        );

    \I__3750\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24363\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__24363\,
            I => \pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26\
        );

    \I__3748\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24354\
        );

    \I__3747\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24354\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__24354\,
            I => \pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__24351\,
            I => \N__24348\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24344\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__24347\,
            I => \N__24341\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24344\,
            I => \N__24338\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24335\
        );

    \I__3740\ : Span4Mux_v
    port map (
            O => \N__24338\,
            I => \N__24332\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24329\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__24332\,
            I => \pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__24329\,
            I => \pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__24315\,
            I => \pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24308\
        );

    \I__3731\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24305\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24308\,
            I => \pid_alt.error_d_reg_prevZ0Z_25\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__24305\,
            I => \pid_alt.error_d_reg_prevZ0Z_25\
        );

    \I__3728\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24295\
        );

    \I__3727\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24290\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24290\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24295\,
            I => \N__24285\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__24290\,
            I => \N__24285\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__3722\ : Span4Mux_h
    port map (
            O => \N__24282\,
            I => \N__24279\
        );

    \I__3721\ : Span4Mux_h
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__3720\ : Span4Mux_v
    port map (
            O => \N__24276\,
            I => \N__24273\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__24273\,
            I => \pid_alt.error_d_regZ0Z_25\
        );

    \I__3718\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24267\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24267\,
            I => \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__24264\,
            I => \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__24261\,
            I => \N__24257\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24254\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24248\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24251\,
            I => \pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__24248\,
            I => \pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__24243\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__24240\,
            I => \N__24236\
        );

    \I__3707\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24233\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24230\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24227\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24224\
        );

    \I__3703\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24221\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__24224\,
            I => \pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__24221\,
            I => \pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23\
        );

    \I__3700\ : InMux
    port map (
            O => \N__24216\,
            I => \N__24213\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__24210\,
            I => \pid_alt.un9lto29_i_a2_0_and\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24204\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__24204\,
            I => \N__24201\
        );

    \I__3695\ : Odrv4
    port map (
            O => \N__24201\,
            I => \pid_alt.N_96\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__24198\,
            I => \N__24192\
        );

    \I__3693\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24185\
        );

    \I__3692\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24185\
        );

    \I__3691\ : InMux
    port map (
            O => \N__24195\,
            I => \N__24185\
        );

    \I__3690\ : InMux
    port map (
            O => \N__24192\,
            I => \N__24182\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24179\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__24182\,
            I => \N__24176\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__24179\,
            I => \N__24173\
        );

    \I__3686\ : Odrv12
    port map (
            O => \N__24176\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__24173\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__3684\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24158\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24158\
        );

    \I__3682\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24158\
        );

    \I__3681\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24155\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24152\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__24155\,
            I => \N__24147\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__24152\,
            I => \N__24147\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__24147\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__3674\ : Odrv12
    port map (
            O => \N__24138\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_4\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24132\,
            I => \N__24129\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__24129\,
            I => \N__24125\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24122\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__24125\,
            I => \N__24119\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__24122\,
            I => \N__24116\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__24119\,
            I => \N__24113\
        );

    \I__3666\ : Span12Mux_s9_h
    port map (
            O => \N__24116\,
            I => \N__24110\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__24113\,
            I => \N__24107\
        );

    \I__3664\ : Odrv12
    port map (
            O => \N__24110\,
            I => \pid_alt.state_RNIFCSD1Z0Z_0\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__24107\,
            I => \pid_alt.state_RNIFCSD1Z0Z_0\
        );

    \I__3662\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24096\
        );

    \I__3661\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24089\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24089\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24089\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24096\,
            I => \N__24086\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24083\
        );

    \I__3656\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24080\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__24083\,
            I => \N__24077\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__24080\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__24077\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24066\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24066\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__24066\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\
        );

    \I__3649\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24057\
        );

    \I__3648\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24057\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24054\
        );

    \I__3646\ : Span12Mux_v
    port map (
            O => \N__24054\,
            I => \N__24051\
        );

    \I__3645\ : Odrv12
    port map (
            O => \N__24051\,
            I => \pid_alt.error_p_regZ0Z_4\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__24048\,
            I => \pid_alt.un1_reset_0_i_cascade_\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24039\
        );

    \I__3641\ : Span4Mux_h
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__24036\,
            I => \pid_alt.pid_preregZ0Z_26\
        );

    \I__3639\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24027\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__24024\,
            I => \pid_alt.pid_preregZ0Z_25\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24015\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__24012\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__24012\,
            I => \N__24009\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__24009\,
            I => \pid_alt.pid_preregZ0Z_27\
        );

    \I__3630\ : InMux
    port map (
            O => \N__24006\,
            I => \N__24003\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__3628\ : Span4Mux_h
    port map (
            O => \N__24000\,
            I => \N__23997\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__23997\,
            I => \pid_alt.pid_preregZ0Z_24\
        );

    \I__3626\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23991\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23987\
        );

    \I__3624\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__23987\,
            I => \pid_alt.un9lto29_i_a2_5_and\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__23984\,
            I => \pid_alt.un9lto29_i_a2_5_and\
        );

    \I__3621\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23976\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__23976\,
            I => \N__23969\
        );

    \I__3619\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23966\
        );

    \I__3618\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23961\
        );

    \I__3617\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23961\
        );

    \I__3616\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23958\
        );

    \I__3615\ : Span4Mux_v
    port map (
            O => \N__23969\,
            I => \N__23953\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__23966\,
            I => \N__23953\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__23961\,
            I => \N__23950\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__23958\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__23953\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__23950\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__3609\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23936\
        );

    \I__3608\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23936\
        );

    \I__3607\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23933\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__23936\,
            I => \N__23930\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__23933\,
            I => \pid_alt.N_124\
        );

    \I__3604\ : Odrv12
    port map (
            O => \N__23930\,
            I => \pid_alt.N_124\
        );

    \I__3603\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23922\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23917\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23912\
        );

    \I__3600\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23912\
        );

    \I__3599\ : Span4Mux_v
    port map (
            O => \N__23917\,
            I => \N__23907\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23907\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__23907\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__23904\,
            I => \N__23901\
        );

    \I__3595\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23898\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__23898\,
            I => \N__23895\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__23895\,
            I => \pid_alt.N_12_i\
        );

    \I__3592\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23888\
        );

    \I__3591\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23885\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23882\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__23885\,
            I => \pid_alt.un9lto29_i_a2_3_and\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__23882\,
            I => \pid_alt.un9lto29_i_a2_3_and\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__3586\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__23868\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_0\
        );

    \I__3583\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23861\
        );

    \I__3582\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23858\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23855\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__23858\,
            I => \pid_alt.un9lto29_i_a2_4_and\
        );

    \I__3579\ : Odrv4
    port map (
            O => \N__23855\,
            I => \pid_alt.un9lto29_i_a2_4_and\
        );

    \I__3578\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__23847\,
            I => \N__23844\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__23844\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_5\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__23841\,
            I => \pid_alt.N_123_cascade_\
        );

    \I__3574\ : InMux
    port map (
            O => \N__23838\,
            I => \N__23835\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__23835\,
            I => \N__23832\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__23832\,
            I => \N__23826\
        );

    \I__3571\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23819\
        );

    \I__3570\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23819\
        );

    \I__3569\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23819\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__23826\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__23819\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__3566\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23807\
        );

    \I__3565\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23807\
        );

    \I__3564\ : InMux
    port map (
            O => \N__23812\,
            I => \N__23804\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__23807\,
            I => \pid_alt.N_123\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__23804\,
            I => \pid_alt.N_123\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__23799\,
            I => \pid_alt.N_106_cascade_\
        );

    \I__3560\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23793\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__23793\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0\
        );

    \I__3558\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23787\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__23787\,
            I => \pid_alt.N_100\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__23784\,
            I => \pid_alt.N_91_1_cascade_\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__23781\,
            I => \Commands_frame_decoder.N_358_cascade_\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \N__23773\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__23777\,
            I => \N__23770\
        );

    \I__3552\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23765\
        );

    \I__3551\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23765\
        );

    \I__3550\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23762\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__23765\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__23762\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__3547\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__23754\,
            I => \N__23750\
        );

    \I__3545\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23747\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__23750\,
            I => \N__23744\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__23747\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__23744\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__3541\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23733\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__23730\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__3537\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__23724\,
            I => \Commands_frame_decoder.N_327\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__23721\,
            I => \N__23718\
        );

    \I__3534\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23712\
        );

    \I__3533\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23712\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__23712\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__3531\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23705\
        );

    \I__3530\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23702\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23698\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23695\
        );

    \I__3527\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23692\
        );

    \I__3526\ : Span4Mux_h
    port map (
            O => \N__23698\,
            I => \N__23687\
        );

    \I__3525\ : Span4Mux_v
    port map (
            O => \N__23695\,
            I => \N__23687\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__23692\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__23687\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3521\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23675\
        );

    \I__3520\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23672\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__23675\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__23672\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__3517\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23664\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23660\
        );

    \I__3515\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23657\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__23660\,
            I => \N__23652\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23652\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__23652\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__3511\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23644\
        );

    \I__3510\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23639\
        );

    \I__3509\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23639\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__23644\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__23639\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__3506\ : InMux
    port map (
            O => \N__23634\,
            I => \bfn_9_6_0_\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__23631\,
            I => \N__23626\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \N__23623\
        );

    \I__3503\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23620\
        );

    \I__3502\ : InMux
    port map (
            O => \N__23626\,
            I => \N__23615\
        );

    \I__3501\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23615\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__23620\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__23615\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__3498\ : InMux
    port map (
            O => \N__23610\,
            I => \Commands_frame_decoder.un1_WDT_cry_8\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__23607\,
            I => \N__23602\
        );

    \I__3496\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23599\
        );

    \I__3495\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23594\
        );

    \I__3494\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23594\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__23599\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__23594\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__3491\ : InMux
    port map (
            O => \N__23589\,
            I => \Commands_frame_decoder.un1_WDT_cry_9\
        );

    \I__3490\ : InMux
    port map (
            O => \N__23586\,
            I => \Commands_frame_decoder.un1_WDT_cry_10\
        );

    \I__3489\ : InMux
    port map (
            O => \N__23583\,
            I => \Commands_frame_decoder.un1_WDT_cry_11\
        );

    \I__3488\ : InMux
    port map (
            O => \N__23580\,
            I => \Commands_frame_decoder.un1_WDT_cry_12\
        );

    \I__3487\ : InMux
    port map (
            O => \N__23577\,
            I => \Commands_frame_decoder.un1_WDT_cry_13\
        );

    \I__3486\ : InMux
    port map (
            O => \N__23574\,
            I => \Commands_frame_decoder.un1_WDT_cry_14\
        );

    \I__3485\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23568\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__23568\,
            I => uart_input_pc_c
        );

    \I__3483\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23561\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__3480\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23552\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__23555\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__23552\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3477\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__23544\,
            I => \Commands_frame_decoder.WDTZ0Z_0\
        );

    \I__3475\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__23538\,
            I => \Commands_frame_decoder.WDTZ0Z_1\
        );

    \I__3473\ : InMux
    port map (
            O => \N__23535\,
            I => \Commands_frame_decoder.un1_WDT_cry_0\
        );

    \I__3472\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23529\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__23529\,
            I => \Commands_frame_decoder.WDTZ0Z_2\
        );

    \I__3470\ : InMux
    port map (
            O => \N__23526\,
            I => \Commands_frame_decoder.un1_WDT_cry_1\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__23520\,
            I => \Commands_frame_decoder.WDTZ0Z_3\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23517\,
            I => \Commands_frame_decoder.un1_WDT_cry_2\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23514\,
            I => \N__23509\
        );

    \I__3465\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23504\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23504\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__23509\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23504\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__3461\ : InMux
    port map (
            O => \N__23499\,
            I => \Commands_frame_decoder.un1_WDT_cry_3\
        );

    \I__3460\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23491\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23486\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23486\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__23491\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__23486\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__3455\ : InMux
    port map (
            O => \N__23481\,
            I => \Commands_frame_decoder.un1_WDT_cry_4\
        );

    \I__3454\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23473\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23470\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23467\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__23473\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__23470\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__23467\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23460\,
            I => \Commands_frame_decoder.un1_WDT_cry_5\
        );

    \I__3447\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23452\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23449\
        );

    \I__3445\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23446\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__23452\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__23449\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__23446\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23439\,
            I => \Commands_frame_decoder.un1_WDT_cry_6\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__3439\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__23430\,
            I => \pid_alt.error_axbZ0Z_1\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__3436\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__23421\,
            I => \pid_alt.error_axbZ0Z_12\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__3433\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__23412\,
            I => \pid_alt.error_axbZ0Z_13\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__3430\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__23403\,
            I => \pid_alt.error_axbZ0Z_14\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__23400\,
            I => \N__23397\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__23394\,
            I => \pid_alt.error_axbZ0Z_2\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__3422\ : Sp12to4
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__3421\ : Span12Mux_s9_h
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__3420\ : Odrv12
    port map (
            O => \N__23376\,
            I => alt_ki_0
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__3418\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__23367\,
            I => drone_altitude_i_9
        );

    \I__3416\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23360\
        );

    \I__3415\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23357\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__23357\,
            I => alt_command_0
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__23354\,
            I => alt_command_0
        );

    \I__3411\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__3409\ : Span4Mux_h
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__23340\,
            I => \N__23337\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__23337\,
            I => \pid_alt.O_1_9\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__23334\,
            I => \N__23331\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23325\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23325\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__23325\,
            I => \pid_alt.error_d_reg_prevZ0Z_21\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23313\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23313\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23320\,
            I => \N__23313\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__3398\ : Span4Mux_h
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__3396\ : Sp12to4
    port map (
            O => \N__23304\,
            I => \N__23301\
        );

    \I__3395\ : Odrv12
    port map (
            O => \N__23301\,
            I => \pid_alt.error_d_regZ0Z_21\
        );

    \I__3394\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23295\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__23295\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__23292\,
            I => \N__23288\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23285\
        );

    \I__3390\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23282\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23285\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__23282\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23271\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23271\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__3384\ : Span4Mux_h
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__3383\ : Span4Mux_h
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__23262\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__23259\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__23247\,
            I => \pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__23244\,
            I => \N__23240\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23237\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23234\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23237\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__23234\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__23229\,
            I => \N__23226\
        );

    \I__3370\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23223\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__23223\,
            I => \pid_alt.error_axbZ0Z_3\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__23220\,
            I => \N__23217\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23214\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__23214\,
            I => drone_altitude_i_10
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__23211\,
            I => \N__23208\
        );

    \I__3364\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23205\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__23205\,
            I => drone_altitude_i_11
        );

    \I__3362\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__3360\ : Span4Mux_h
    port map (
            O => \N__23196\,
            I => \N__23192\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23189\
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__23192\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__23189\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23184\,
            I => \N__23181\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__23181\,
            I => \N__23178\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__23178\,
            I => \N__23175\
        );

    \I__3353\ : Span4Mux_h
    port map (
            O => \N__23175\,
            I => \N__23171\
        );

    \I__3352\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23168\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__23171\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23168\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23163\,
            I => \N__23160\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23157\
        );

    \I__3347\ : Odrv12
    port map (
            O => \N__23157\,
            I => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\
        );

    \I__3346\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23150\
        );

    \I__3345\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23147\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__23147\,
            I => \pid_alt.error_d_reg_prevZ0Z_26\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__23144\,
            I => \pid_alt.error_d_reg_prevZ0Z_26\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23133\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23133\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23129\
        );

    \I__3338\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23126\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__23129\,
            I => \N__23123\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23120\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__23123\,
            I => \N__23117\
        );

    \I__3334\ : Span4Mux_h
    port map (
            O => \N__23120\,
            I => \N__23114\
        );

    \I__3333\ : Span4Mux_v
    port map (
            O => \N__23117\,
            I => \N__23111\
        );

    \I__3332\ : Sp12to4
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__3331\ : Sp12to4
    port map (
            O => \N__23111\,
            I => \N__23103\
        );

    \I__3330\ : Span12Mux_v
    port map (
            O => \N__23108\,
            I => \N__23103\
        );

    \I__3329\ : Odrv12
    port map (
            O => \N__23103\,
            I => \pid_alt.error_d_regZ0Z_26\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23097\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23097\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\
        );

    \I__3326\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23090\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23087\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__23090\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__23087\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__23082\,
            I => \N__23078\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__23081\,
            I => \N__23075\
        );

    \I__3320\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23072\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23069\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23066\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23063\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__23066\,
            I => \N__23060\
        );

    \I__3315\ : Span4Mux_h
    port map (
            O => \N__23063\,
            I => \N__23057\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__23060\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__23057\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__23046\
        );

    \I__3310\ : Span4Mux_v
    port map (
            O => \N__23046\,
            I => \N__23042\
        );

    \I__3309\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23039\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__23042\,
            I => \pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__23039\,
            I => \pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__23031\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23022\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23022\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__3301\ : Span4Mux_h
    port map (
            O => \N__23019\,
            I => \N__23016\
        );

    \I__3300\ : Odrv4
    port map (
            O => \N__23016\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__23013\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__3297\ : InMux
    port map (
            O => \N__23007\,
            I => \N__23004\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__23001\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21\
        );

    \I__3294\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22994\
        );

    \I__3293\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22991\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__22994\,
            I => \N__22988\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__22991\,
            I => \pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__22988\,
            I => \pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__22983\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\
        );

    \I__3288\ : InMux
    port map (
            O => \N__22980\,
            I => \N__22977\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__22977\,
            I => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\
        );

    \I__3286\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__22971\,
            I => \N__22967\
        );

    \I__3284\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22964\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__22967\,
            I => \N__22959\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__22964\,
            I => \N__22959\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__22959\,
            I => \N__22956\
        );

    \I__3280\ : Span4Mux_h
    port map (
            O => \N__22956\,
            I => \N__22953\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__22953\,
            I => \pid_alt.error_p_regZ0Z_10\
        );

    \I__3278\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22943\
        );

    \I__3276\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22940\
        );

    \I__3275\ : Span4Mux_v
    port map (
            O => \N__22943\,
            I => \N__22937\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__22940\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__22937\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3272\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22927\
        );

    \I__3271\ : InMux
    port map (
            O => \N__22931\,
            I => \N__22922\
        );

    \I__3270\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22922\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__22927\,
            I => \N__22919\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__22919\,
            I => \N__22913\
        );

    \I__3266\ : Span4Mux_h
    port map (
            O => \N__22916\,
            I => \N__22910\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22907\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__22910\,
            I => \pid_alt.error_d_regZ0Z_10\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__22907\,
            I => \pid_alt.error_d_regZ0Z_10\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__22902\,
            I => \N__22898\
        );

    \I__3261\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22895\
        );

    \I__3260\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22892\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__22895\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__22892\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__3257\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22881\
        );

    \I__3256\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22881\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__3254\ : Span4Mux_h
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__3253\ : Span4Mux_v
    port map (
            O => \N__22875\,
            I => \N__22872\
        );

    \I__3252\ : Span4Mux_h
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__22869\,
            I => \pid_alt.error_p_regZ0Z_9\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__3249\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22857\
        );

    \I__3248\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22857\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__22857\,
            I => \pid_alt.error_d_reg_prevZ0Z_9\
        );

    \I__3246\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22845\
        );

    \I__3245\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22845\
        );

    \I__3244\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22845\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__3242\ : Span4Mux_v
    port map (
            O => \N__22842\,
            I => \N__22839\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__22833\,
            I => \pid_alt.error_d_regZ0Z_9\
        );

    \I__3238\ : InMux
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__22827\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\
        );

    \I__3236\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22818\
        );

    \I__3235\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22818\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__22812\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\
        );

    \I__3231\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22805\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \N__22802\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__22805\,
            I => \N__22799\
        );

    \I__3228\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22796\
        );

    \I__3227\ : Span4Mux_v
    port map (
            O => \N__22799\,
            I => \N__22793\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22790\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__22793\,
            I => \N__22785\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__22790\,
            I => \N__22785\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__22785\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__22782\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\
        );

    \I__3221\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__22776\,
            I => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__22773\,
            I => \N__22769\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__22772\,
            I => \N__22766\
        );

    \I__3217\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22763\
        );

    \I__3216\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22760\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22755\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__22760\,
            I => \N__22755\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__22755\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\
        );

    \I__3212\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__3210\ : Span4Mux_h
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__22743\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__22740\,
            I => \N__22736\
        );

    \I__3207\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22733\
        );

    \I__3206\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22730\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22727\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22724\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__22727\,
            I => \N__22719\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__22724\,
            I => \N__22719\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__22719\,
            I => \pid_alt.pid_preregZ0Z_29\
        );

    \I__3200\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22710\
        );

    \I__3199\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22710\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__22710\,
            I => \pid_alt.pid_preregZ0Z_14\
        );

    \I__3197\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__22704\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__22701\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\
        );

    \I__3194\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__22695\,
            I => \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \N__22688\
        );

    \I__3191\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22685\
        );

    \I__3190\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22682\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__22685\,
            I => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__22682\,
            I => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\
        );

    \I__3187\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22674\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__22674\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__22671\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_\
        );

    \I__3184\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__22665\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__22662\,
            I => \N__22659\
        );

    \I__3181\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__22656\,
            I => \pid_alt.N_232_i\
        );

    \I__3179\ : InMux
    port map (
            O => \N__22653\,
            I => \bfn_8_12_0_\
        );

    \I__3178\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22644\
        );

    \I__3177\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22641\
        );

    \I__3176\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22636\
        );

    \I__3175\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22636\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__22644\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__22641\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__22636\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__3171\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__22626\,
            I => \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\
        );

    \I__3169\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22620\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22617\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__22617\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3166\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22611\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22608\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__22608\,
            I => \pid_alt.pid_preregZ0Z_21\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__22605\,
            I => \N__22602\
        );

    \I__3162\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__22596\,
            I => \pid_alt.pid_preregZ0Z_23\
        );

    \I__3159\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__22587\,
            I => \pid_alt.pid_preregZ0Z_20\
        );

    \I__3156\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__22578\,
            I => \pid_alt.source_pid10lt4_0\
        );

    \I__3153\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__22569\,
            I => \pid_alt.un9lto29_i_a2_2_and\
        );

    \I__3150\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22562\
        );

    \I__3149\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22559\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22556\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__3146\ : Odrv12
    port map (
            O => \N__22556\,
            I => \pid_alt.pid_preregZ0Z_28\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__22553\,
            I => \pid_alt.pid_preregZ0Z_28\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__3143\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22539\
        );

    \I__3142\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22539\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__22539\,
            I => \N__22536\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__22536\,
            I => \pid_alt.pid_preregZ0Z_15\
        );

    \I__3139\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22522\
        );

    \I__3138\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22522\
        );

    \I__3137\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22522\
        );

    \I__3136\ : InMux
    port map (
            O => \N__22530\,
            I => \N__22517\
        );

    \I__3135\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22517\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22509\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__22517\,
            I => \N__22509\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22502\
        );

    \I__3131\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22502\
        );

    \I__3130\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22502\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__22509\,
            I => \N__22497\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22502\,
            I => \N__22497\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__22497\,
            I => \dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15\
        );

    \I__3126\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22485\
        );

    \I__3125\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22485\
        );

    \I__3124\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22485\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__22485\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__3122\ : CEMux
    port map (
            O => \N__22482\,
            I => \N__22478\
        );

    \I__3121\ : CEMux
    port map (
            O => \N__22481\,
            I => \N__22475\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__22478\,
            I => \N__22467\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22467\
        );

    \I__3118\ : CEMux
    port map (
            O => \N__22474\,
            I => \N__22464\
        );

    \I__3117\ : CEMux
    port map (
            O => \N__22473\,
            I => \N__22461\
        );

    \I__3116\ : CEMux
    port map (
            O => \N__22472\,
            I => \N__22458\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__22467\,
            I => \N__22451\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__22464\,
            I => \N__22451\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22451\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22448\
        );

    \I__3111\ : Span4Mux_v
    port map (
            O => \N__22451\,
            I => \N__22443\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__22448\,
            I => \N__22443\
        );

    \I__3109\ : Span4Mux_v
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__22440\,
            I => \N__22437\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__22434\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__3104\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__22422\,
            I => \Commands_frame_decoder.N_354\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__22416\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__3099\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22407\
        );

    \I__3098\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22407\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__22407\,
            I => \Commands_frame_decoder.stateZ0Z_8\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__3095\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22398\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__22398\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__22395\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_\
        );

    \I__3092\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22386\
        );

    \I__3091\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22383\
        );

    \I__3090\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22378\
        );

    \I__3089\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22378\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__22386\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__22383\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22378\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__3084\ : InMux
    port map (
            O => \N__22368\,
            I => \N__22363\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22358\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22358\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__22363\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__22358\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__22353\,
            I => \Commands_frame_decoder.WDT8lt12_0_cascade_\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22347\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22347\,
            I => \Commands_frame_decoder.state_0_sqmuxacf1\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22341\,
            I => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__22332\,
            I => \uart_drone_sync.aux_2__0__0_0\
        );

    \I__3071\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__22326\,
            I => \uart_drone_sync.aux_3__0__0_0\
        );

    \I__3069\ : SRMux
    port map (
            O => \N__22323\,
            I => \N__22319\
        );

    \I__3068\ : SRMux
    port map (
            O => \N__22322\,
            I => \N__22316\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22313\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22310\
        );

    \I__3065\ : Span4Mux_h
    port map (
            O => \N__22313\,
            I => \N__22307\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__22310\,
            I => \N__22304\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__22307\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__22304\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__22299\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__22296\,
            I => \Commands_frame_decoder.N_322_0_cascade_\
        );

    \I__3059\ : IoInMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__3057\ : Span4Mux_s1_v
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__22284\,
            I => \pid_alt.N_410_0\
        );

    \I__3055\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22278\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__22278\,
            I => \uart_drone_sync.aux_1__0__0_0\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22272\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22269\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__22269\,
            I => uart_input_drone_c
        );

    \I__3050\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22263\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22263\,
            I => \uart_drone_sync.aux_0__0__0_0\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__22260\,
            I => \Commands_frame_decoder.WDT8lto13_1_cascade_\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__22254\,
            I => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \Commands_frame_decoder.WDT8lto9_3_cascade_\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22244\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22240\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22237\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22234\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22231\
        );

    \I__3039\ : Span12Mux_s6_h
    port map (
            O => \N__22237\,
            I => \N__22228\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22225\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__22231\,
            I => \N__22222\
        );

    \I__3036\ : Span12Mux_h
    port map (
            O => \N__22228\,
            I => \N__22217\
        );

    \I__3035\ : Span12Mux_s7_h
    port map (
            O => \N__22225\,
            I => \N__22217\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__22222\,
            I => \N__22214\
        );

    \I__3033\ : Odrv12
    port map (
            O => \N__22217\,
            I => \pid_alt.error_13\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__22214\,
            I => \pid_alt.error_13\
        );

    \I__3031\ : InMux
    port map (
            O => \N__22209\,
            I => \pid_alt.error_cry_12\
        );

    \I__3030\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__3028\ : Span4Mux_s2_h
    port map (
            O => \N__22200\,
            I => \N__22197\
        );

    \I__3027\ : Span4Mux_h
    port map (
            O => \N__22197\,
            I => \N__22193\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22190\
        );

    \I__3025\ : Span4Mux_h
    port map (
            O => \N__22193\,
            I => \N__22186\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22183\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22180\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__22186\,
            I => \N__22177\
        );

    \I__3021\ : Span4Mux_s3_h
    port map (
            O => \N__22183\,
            I => \N__22174\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__22180\,
            I => \N__22171\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__22177\,
            I => \N__22166\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__22174\,
            I => \N__22166\
        );

    \I__3017\ : Span4Mux_s3_h
    port map (
            O => \N__22171\,
            I => \N__22163\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__22166\,
            I => \N__22158\
        );

    \I__3015\ : Span4Mux_h
    port map (
            O => \N__22163\,
            I => \N__22158\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__22158\,
            I => \pid_alt.error_14\
        );

    \I__3013\ : InMux
    port map (
            O => \N__22155\,
            I => \pid_alt.error_cry_13\
        );

    \I__3012\ : InMux
    port map (
            O => \N__22152\,
            I => \pid_alt.error_cry_14\
        );

    \I__3011\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__3009\ : Span4Mux_s2_h
    port map (
            O => \N__22143\,
            I => \N__22140\
        );

    \I__3008\ : Span4Mux_h
    port map (
            O => \N__22140\,
            I => \N__22136\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22133\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__22136\,
            I => \N__22129\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__22133\,
            I => \N__22126\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22123\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__22129\,
            I => \N__22120\
        );

    \I__3002\ : Span4Mux_s3_h
    port map (
            O => \N__22126\,
            I => \N__22117\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22123\,
            I => \N__22114\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__22120\,
            I => \N__22109\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__22117\,
            I => \N__22109\
        );

    \I__2998\ : Span4Mux_s3_h
    port map (
            O => \N__22114\,
            I => \N__22106\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__22109\,
            I => \N__22101\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__22106\,
            I => \N__22101\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__22101\,
            I => \pid_alt.error_15\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22095\,
            I => alt_command_4
        );

    \I__2992\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__22086\,
            I => alt_command_5
        );

    \I__2989\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__22077\,
            I => alt_command_6
        );

    \I__2986\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__22071\,
            I => alt_command_7
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22059\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__22056\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__22053\,
            I => \N__22048\
        );

    \I__2978\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22044\
        );

    \I__2977\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22041\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22038\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22035\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__22044\,
            I => \N__22030\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22030\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__22038\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22035\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27\
        );

    \I__2970\ : Odrv12
    port map (
            O => \N__22030\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__2968\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22016\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22010\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22010\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22005\
        );

    \I__2964\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__22002\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21997\
        );

    \I__2962\ : InMux
    port map (
            O => \N__22008\,
            I => \N__21997\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__22005\,
            I => \pid_alt.un1_pid_prereg_296_1\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__22002\,
            I => \pid_alt.un1_pid_prereg_296_1\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__21997\,
            I => \pid_alt.un1_pid_prereg_296_1\
        );

    \I__2958\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__21984\,
            I => \N__21981\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__21981\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21974\
        );

    \I__2953\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21971\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21968\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__21971\,
            I => alt_command_1
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__21968\,
            I => alt_command_1
        );

    \I__2949\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__2947\ : Span4Mux_s2_h
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__21954\,
            I => \N__21950\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21953\,
            I => \N__21947\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__21950\,
            I => \N__21943\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21940\
        );

    \I__2942\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21937\
        );

    \I__2941\ : Span4Mux_h
    port map (
            O => \N__21943\,
            I => \N__21934\
        );

    \I__2940\ : Span4Mux_s3_h
    port map (
            O => \N__21940\,
            I => \N__21931\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__21937\,
            I => \N__21928\
        );

    \I__2938\ : Span4Mux_h
    port map (
            O => \N__21934\,
            I => \N__21923\
        );

    \I__2937\ : Span4Mux_h
    port map (
            O => \N__21931\,
            I => \N__21923\
        );

    \I__2936\ : Span4Mux_s3_h
    port map (
            O => \N__21928\,
            I => \N__21920\
        );

    \I__2935\ : Span4Mux_v
    port map (
            O => \N__21923\,
            I => \N__21915\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__21920\,
            I => \N__21915\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__21915\,
            I => \pid_alt.error_5\
        );

    \I__2932\ : InMux
    port map (
            O => \N__21912\,
            I => \pid_alt.error_cry_4\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__21909\,
            I => \N__21905\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__21908\,
            I => \N__21902\
        );

    \I__2929\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21899\
        );

    \I__2928\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21896\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__21899\,
            I => alt_command_2
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__21896\,
            I => alt_command_2
        );

    \I__2925\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21886\
        );

    \I__2924\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21883\
        );

    \I__2923\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21880\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__21886\,
            I => \N__21877\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21874\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21871\
        );

    \I__2919\ : Span12Mux_s6_h
    port map (
            O => \N__21877\,
            I => \N__21868\
        );

    \I__2918\ : Span4Mux_s3_h
    port map (
            O => \N__21874\,
            I => \N__21865\
        );

    \I__2917\ : Span12Mux_s7_h
    port map (
            O => \N__21871\,
            I => \N__21860\
        );

    \I__2916\ : Span12Mux_h
    port map (
            O => \N__21868\,
            I => \N__21860\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__21865\,
            I => \N__21857\
        );

    \I__2914\ : Odrv12
    port map (
            O => \N__21860\,
            I => \pid_alt.error_6\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__21857\,
            I => \pid_alt.error_6\
        );

    \I__2912\ : InMux
    port map (
            O => \N__21852\,
            I => \pid_alt.error_cry_5\
        );

    \I__2911\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21845\
        );

    \I__2910\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21842\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__21845\,
            I => alt_command_3
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__21842\,
            I => alt_command_3
        );

    \I__2907\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__21834\,
            I => \N__21831\
        );

    \I__2905\ : Span4Mux_s2_h
    port map (
            O => \N__21831\,
            I => \N__21827\
        );

    \I__2904\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21824\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__21827\,
            I => \N__21821\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21817\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__21821\,
            I => \N__21814\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21811\
        );

    \I__2899\ : Span4Mux_s3_h
    port map (
            O => \N__21817\,
            I => \N__21808\
        );

    \I__2898\ : Span4Mux_h
    port map (
            O => \N__21814\,
            I => \N__21805\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21802\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__21808\,
            I => \N__21799\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__21805\,
            I => \N__21796\
        );

    \I__2894\ : Span4Mux_s3_h
    port map (
            O => \N__21802\,
            I => \N__21793\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__21799\,
            I => \N__21786\
        );

    \I__2892\ : Span4Mux_v
    port map (
            O => \N__21796\,
            I => \N__21786\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__21793\,
            I => \N__21786\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__21786\,
            I => \pid_alt.error_7\
        );

    \I__2889\ : InMux
    port map (
            O => \N__21783\,
            I => \pid_alt.error_cry_6\
        );

    \I__2888\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__2886\ : Span4Mux_s2_h
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__21771\,
            I => \N__21767\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21764\
        );

    \I__2883\ : Span4Mux_h
    port map (
            O => \N__21767\,
            I => \N__21760\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21757\
        );

    \I__2881\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21754\
        );

    \I__2880\ : Span4Mux_h
    port map (
            O => \N__21760\,
            I => \N__21751\
        );

    \I__2879\ : Span4Mux_s3_h
    port map (
            O => \N__21757\,
            I => \N__21748\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21745\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__21751\,
            I => \N__21740\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__21748\,
            I => \N__21740\
        );

    \I__2875\ : Span4Mux_s3_h
    port map (
            O => \N__21745\,
            I => \N__21737\
        );

    \I__2874\ : Span4Mux_v
    port map (
            O => \N__21740\,
            I => \N__21732\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__21737\,
            I => \N__21732\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__21732\,
            I => \pid_alt.error_8\
        );

    \I__2871\ : InMux
    port map (
            O => \N__21729\,
            I => \bfn_7_20_0_\
        );

    \I__2870\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__2868\ : Span4Mux_s2_h
    port map (
            O => \N__21720\,
            I => \N__21717\
        );

    \I__2867\ : Span4Mux_h
    port map (
            O => \N__21717\,
            I => \N__21713\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21710\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21706\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21703\
        );

    \I__2863\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21700\
        );

    \I__2862\ : Span4Mux_h
    port map (
            O => \N__21706\,
            I => \N__21697\
        );

    \I__2861\ : Span4Mux_s3_h
    port map (
            O => \N__21703\,
            I => \N__21694\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N__21691\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__21697\,
            I => \N__21686\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__21694\,
            I => \N__21686\
        );

    \I__2857\ : Span4Mux_s3_h
    port map (
            O => \N__21691\,
            I => \N__21683\
        );

    \I__2856\ : Span4Mux_v
    port map (
            O => \N__21686\,
            I => \N__21678\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__21683\,
            I => \N__21678\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__21678\,
            I => \pid_alt.error_9\
        );

    \I__2853\ : InMux
    port map (
            O => \N__21675\,
            I => \pid_alt.error_cry_8\
        );

    \I__2852\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__21669\,
            I => \N__21665\
        );

    \I__2850\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21661\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__21665\,
            I => \N__21658\
        );

    \I__2848\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21655\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21652\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__21658\,
            I => \N__21647\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__21655\,
            I => \N__21647\
        );

    \I__2844\ : Span12Mux_s10_v
    port map (
            O => \N__21652\,
            I => \N__21644\
        );

    \I__2843\ : Span4Mux_h
    port map (
            O => \N__21647\,
            I => \N__21641\
        );

    \I__2842\ : Span12Mux_h
    port map (
            O => \N__21644\,
            I => \N__21638\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__21641\,
            I => \N__21635\
        );

    \I__2840\ : Odrv12
    port map (
            O => \N__21638\,
            I => \pid_alt.error_10\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__21635\,
            I => \pid_alt.error_10\
        );

    \I__2838\ : InMux
    port map (
            O => \N__21630\,
            I => \pid_alt.error_cry_9\
        );

    \I__2837\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__2835\ : Span4Mux_s1_h
    port map (
            O => \N__21621\,
            I => \N__21617\
        );

    \I__2834\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21613\
        );

    \I__2833\ : Sp12to4
    port map (
            O => \N__21617\,
            I => \N__21610\
        );

    \I__2832\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21607\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__21613\,
            I => \N__21604\
        );

    \I__2830\ : Span12Mux_s10_v
    port map (
            O => \N__21610\,
            I => \N__21601\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__21607\,
            I => \N__21598\
        );

    \I__2828\ : Span4Mux_s3_h
    port map (
            O => \N__21604\,
            I => \N__21595\
        );

    \I__2827\ : Span12Mux_h
    port map (
            O => \N__21601\,
            I => \N__21590\
        );

    \I__2826\ : Span12Mux_s10_v
    port map (
            O => \N__21598\,
            I => \N__21590\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__21595\,
            I => \N__21587\
        );

    \I__2824\ : Odrv12
    port map (
            O => \N__21590\,
            I => \pid_alt.error_11\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__21587\,
            I => \pid_alt.error_11\
        );

    \I__2822\ : InMux
    port map (
            O => \N__21582\,
            I => \pid_alt.error_cry_10\
        );

    \I__2821\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21576\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__2819\ : Span4Mux_v
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__21570\,
            I => \N__21566\
        );

    \I__2817\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21563\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__21566\,
            I => \N__21559\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21556\
        );

    \I__2814\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21553\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__21559\,
            I => \N__21550\
        );

    \I__2812\ : Span4Mux_v
    port map (
            O => \N__21556\,
            I => \N__21547\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__21553\,
            I => \N__21544\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__21550\,
            I => \N__21541\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__21547\,
            I => \N__21536\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__21544\,
            I => \N__21536\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__21541\,
            I => \N__21531\
        );

    \I__2806\ : Span4Mux_h
    port map (
            O => \N__21536\,
            I => \N__21531\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__21531\,
            I => \pid_alt.error_12\
        );

    \I__2804\ : InMux
    port map (
            O => \N__21528\,
            I => \pid_alt.error_cry_11\
        );

    \I__2803\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21516\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21516\
        );

    \I__2801\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21516\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__21516\,
            I => \N__21513\
        );

    \I__2799\ : Span4Mux_h
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__2798\ : Span4Mux_h
    port map (
            O => \N__21510\,
            I => \N__21507\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__21501\,
            I => \pid_alt.error_d_regZ0Z_27\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2793\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21489\
        );

    \I__2792\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21489\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__21489\,
            I => \pid_alt.error_d_reg_prevZ0Z_27\
        );

    \I__2790\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21482\
        );

    \I__2789\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21479\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__21482\,
            I => \N__21476\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21473\
        );

    \I__2786\ : Span4Mux_v
    port map (
            O => \N__21476\,
            I => \N__21469\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__21473\,
            I => \N__21466\
        );

    \I__2784\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21463\
        );

    \I__2783\ : Span4Mux_h
    port map (
            O => \N__21469\,
            I => \N__21460\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__21466\,
            I => \N__21455\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21455\
        );

    \I__2780\ : Sp12to4
    port map (
            O => \N__21460\,
            I => \N__21452\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__21455\,
            I => \N__21449\
        );

    \I__2778\ : Span12Mux_h
    port map (
            O => \N__21452\,
            I => \N__21446\
        );

    \I__2777\ : Span4Mux_h
    port map (
            O => \N__21449\,
            I => \N__21443\
        );

    \I__2776\ : Odrv12
    port map (
            O => \N__21446\,
            I => \pid_alt.error_1\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__21443\,
            I => \pid_alt.error_1\
        );

    \I__2774\ : InMux
    port map (
            O => \N__21438\,
            I => \pid_alt.error_cry_0\
        );

    \I__2773\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21431\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21427\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21424\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21421\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21418\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__21424\,
            I => \N__21415\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21412\
        );

    \I__2766\ : Span12Mux_s11_v
    port map (
            O => \N__21418\,
            I => \N__21409\
        );

    \I__2765\ : Span4Mux_v
    port map (
            O => \N__21415\,
            I => \N__21404\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__21412\,
            I => \N__21404\
        );

    \I__2763\ : Span12Mux_h
    port map (
            O => \N__21409\,
            I => \N__21401\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__21404\,
            I => \N__21398\
        );

    \I__2761\ : Odrv12
    port map (
            O => \N__21401\,
            I => \pid_alt.error_2\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__21398\,
            I => \pid_alt.error_2\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21393\,
            I => \pid_alt.error_cry_1\
        );

    \I__2758\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__21387\,
            I => \N__21384\
        );

    \I__2756\ : Span4Mux_v
    port map (
            O => \N__21384\,
            I => \N__21380\
        );

    \I__2755\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21376\
        );

    \I__2754\ : Span4Mux_h
    port map (
            O => \N__21380\,
            I => \N__21373\
        );

    \I__2753\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21370\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21367\
        );

    \I__2751\ : Sp12to4
    port map (
            O => \N__21373\,
            I => \N__21364\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__21370\,
            I => \N__21361\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__21367\,
            I => \N__21358\
        );

    \I__2748\ : Span12Mux_h
    port map (
            O => \N__21364\,
            I => \N__21355\
        );

    \I__2747\ : Span12Mux_s11_v
    port map (
            O => \N__21361\,
            I => \N__21352\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__21358\,
            I => \N__21349\
        );

    \I__2745\ : Odrv12
    port map (
            O => \N__21355\,
            I => \pid_alt.error_3\
        );

    \I__2744\ : Odrv12
    port map (
            O => \N__21352\,
            I => \pid_alt.error_3\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__21349\,
            I => \pid_alt.error_3\
        );

    \I__2742\ : InMux
    port map (
            O => \N__21342\,
            I => \pid_alt.error_cry_2\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2739\ : Span4Mux_s2_h
    port map (
            O => \N__21333\,
            I => \N__21330\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__21330\,
            I => \N__21326\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21323\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__21326\,
            I => \N__21319\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21316\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21313\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__21319\,
            I => \N__21310\
        );

    \I__2732\ : Span4Mux_s3_h
    port map (
            O => \N__21316\,
            I => \N__21307\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21313\,
            I => \N__21304\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__21310\,
            I => \N__21299\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__21307\,
            I => \N__21299\
        );

    \I__2728\ : Span4Mux_s3_h
    port map (
            O => \N__21304\,
            I => \N__21296\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__21299\,
            I => \N__21291\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__21296\,
            I => \N__21291\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__21291\,
            I => \pid_alt.error_4\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21288\,
            I => \pid_alt.error_cry_3\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21285\,
            I => \pid_alt.un1_pid_prereg_0_cry_28\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21282\,
            I => \pid_alt.un1_pid_prereg_0_cry_29\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21276\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__21276\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__21273\,
            I => \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21267\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__21264\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26\
        );

    \I__2715\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21257\
        );

    \I__2714\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21254\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__21257\,
            I => \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__21254\,
            I => \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__21249\,
            I => \pid_alt.un1_pid_prereg_296_1_cascade_\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__21246\,
            I => \N__21243\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21240\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21240\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__2705\ : Odrv12
    port map (
            O => \N__21231\,
            I => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__21228\,
            I => \N__21224\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__21227\,
            I => \N__21221\
        );

    \I__2702\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21218\
        );

    \I__2701\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21215\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21212\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21215\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__21212\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21207\,
            I => \pid_alt.un1_pid_prereg_0_cry_19\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21204\,
            I => \pid_alt.un1_pid_prereg_0_cry_20\
        );

    \I__2695\ : InMux
    port map (
            O => \N__21201\,
            I => \pid_alt.un1_pid_prereg_0_cry_21\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \N__21195\
        );

    \I__2693\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__21186\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21183\,
            I => \bfn_7_16_0_\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21180\,
            I => \pid_alt.un1_pid_prereg_0_cry_23\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21177\,
            I => \pid_alt.un1_pid_prereg_0_cry_24\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21174\,
            I => \pid_alt.un1_pid_prereg_0_cry_25\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21171\,
            I => \pid_alt.un1_pid_prereg_0_cry_26\
        );

    \I__2684\ : InMux
    port map (
            O => \N__21168\,
            I => \pid_alt.un1_pid_prereg_0_cry_27\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21159\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__21159\,
            I => \pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__21156\,
            I => \N__21153\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21147\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__21147\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21144\,
            I => \pid_alt.un1_pid_prereg_0_cry_11\
        );

    \I__2675\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__2672\ : Span4Mux_h
    port map (
            O => \N__21132\,
            I => \N__21129\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__21129\,
            I => \pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21116\
        );

    \I__2667\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21113\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__21116\,
            I => \N__21110\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__21113\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__21110\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21105\,
            I => \pid_alt.un1_pid_prereg_0_cry_12\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21096\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__21096\,
            I => \N__21093\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__21093\,
            I => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21083\
        );

    \I__2656\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21080\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21077\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21074\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__21077\,
            I => \N__21071\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__21074\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__21071\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__2650\ : InMux
    port map (
            O => \N__21066\,
            I => \pid_alt.un1_pid_prereg_0_cry_13\
        );

    \I__2649\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__21060\,
            I => \N__21057\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__21054\,
            I => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21044\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__21047\,
            I => \N__21041\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21038\
        );

    \I__2641\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21035\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__21038\,
            I => \N__21032\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__21035\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__21032\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21027\,
            I => \bfn_7_15_0_\
        );

    \I__2636\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__21021\,
            I => \N__21018\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__21018\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__21015\,
            I => \N__21012\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21008\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21005\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__21008\,
            I => \N__21002\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20999\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__21002\,
            I => \N__20996\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__20999\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__20996\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\
        );

    \I__2625\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__20985\,
            I => \pid_alt.pid_preregZ0Z_16\
        );

    \I__2622\ : InMux
    port map (
            O => \N__20982\,
            I => \pid_alt.un1_pid_prereg_0_cry_15\
        );

    \I__2621\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20976\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__20976\,
            I => \N__20973\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__20973\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__20970\,
            I => \N__20967\
        );

    \I__2617\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20963\
        );

    \I__2616\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20960\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__20963\,
            I => \N__20957\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__20960\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__20957\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__2612\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20949\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20946\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__20946\,
            I => \pid_alt.pid_preregZ0Z_17\
        );

    \I__2609\ : InMux
    port map (
            O => \N__20943\,
            I => \pid_alt.un1_pid_prereg_0_cry_16\
        );

    \I__2608\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__20937\,
            I => \N__20934\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__20934\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__20931\,
            I => \N__20927\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \N__20924\
        );

    \I__2603\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20921\
        );

    \I__2602\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20918\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__20921\,
            I => \N__20915\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__20918\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__20915\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__2598\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20907\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__20904\,
            I => \pid_alt.pid_preregZ0Z_18\
        );

    \I__2595\ : InMux
    port map (
            O => \N__20901\,
            I => \pid_alt.un1_pid_prereg_0_cry_17\
        );

    \I__2594\ : InMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__20892\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__20889\,
            I => \N__20885\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__2589\ : InMux
    port map (
            O => \N__20885\,
            I => \N__20879\
        );

    \I__2588\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20876\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20873\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__20876\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__20873\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__2583\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__2581\ : Odrv4
    port map (
            O => \N__20859\,
            I => \pid_alt.pid_preregZ0Z_19\
        );

    \I__2580\ : InMux
    port map (
            O => \N__20856\,
            I => \pid_alt.un1_pid_prereg_0_cry_18\
        );

    \I__2579\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__20847\,
            I => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\
        );

    \I__2576\ : InMux
    port map (
            O => \N__20844\,
            I => \pid_alt.un1_pid_prereg_0_cry_2\
        );

    \I__2575\ : InMux
    port map (
            O => \N__20841\,
            I => \pid_alt.un1_pid_prereg_0_cry_3\
        );

    \I__2574\ : InMux
    port map (
            O => \N__20838\,
            I => \pid_alt.un1_pid_prereg_0_cry_4\
        );

    \I__2573\ : InMux
    port map (
            O => \N__20835\,
            I => \pid_alt.un1_pid_prereg_0_cry_5\
        );

    \I__2572\ : InMux
    port map (
            O => \N__20832\,
            I => \bfn_7_14_0_\
        );

    \I__2571\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20826\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__20820\,
            I => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\
        );

    \I__2567\ : InMux
    port map (
            O => \N__20817\,
            I => \pid_alt.un1_pid_prereg_0_cry_7\
        );

    \I__2566\ : InMux
    port map (
            O => \N__20814\,
            I => \pid_alt.un1_pid_prereg_0_cry_8\
        );

    \I__2565\ : InMux
    port map (
            O => \N__20811\,
            I => \pid_alt.un1_pid_prereg_0_cry_9\
        );

    \I__2564\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__20802\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10\
        );

    \I__2561\ : InMux
    port map (
            O => \N__20799\,
            I => \pid_alt.un1_pid_prereg_0_cry_10\
        );

    \I__2560\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__2558\ : Odrv12
    port map (
            O => \N__20790\,
            I => \pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1\
        );

    \I__2557\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20784\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__20784\,
            I => \N__20779\
        );

    \I__2555\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20774\
        );

    \I__2554\ : InMux
    port map (
            O => \N__20782\,
            I => \N__20771\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__20779\,
            I => \N__20768\
        );

    \I__2552\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20765\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20762\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20757\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__20771\,
            I => \N__20757\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__20768\,
            I => \N__20754\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20749\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20749\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__20757\,
            I => \N__20746\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__20754\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__20749\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__20746\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__2541\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20735\
        );

    \I__2540\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20731\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20728\
        );

    \I__2538\ : InMux
    port map (
            O => \N__20734\,
            I => \N__20725\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20719\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__20728\,
            I => \N__20714\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__20725\,
            I => \N__20714\
        );

    \I__2534\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20711\
        );

    \I__2533\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20708\
        );

    \I__2532\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20705\
        );

    \I__2531\ : Span4Mux_h
    port map (
            O => \N__20719\,
            I => \N__20702\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__20714\,
            I => \N__20699\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20694\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__20708\,
            I => \N__20694\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20691\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__20702\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__20699\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__20694\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__20691\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__2522\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20678\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__20681\,
            I => \N__20674\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20671\
        );

    \I__2519\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20668\
        );

    \I__2518\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20665\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__20671\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__20668\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__20665\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__2514\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20652\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__20652\,
            I => \dron_frame_decoder_1.state_RNO_1Z0Z_0\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__20649\,
            I => \N__20646\
        );

    \I__2510\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20643\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20639\
        );

    \I__2508\ : InMux
    port map (
            O => \N__20642\,
            I => \N__20636\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__20639\,
            I => \N__20631\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__20636\,
            I => \N__20631\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__20631\,
            I => \N__20628\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__20628\,
            I => \N__20625\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__20625\,
            I => \pid_alt.error_d_reg_prev_i_0\
        );

    \I__2502\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20616\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__20616\,
            I => \N__20613\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__20613\,
            I => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\
        );

    \I__2498\ : InMux
    port map (
            O => \N__20610\,
            I => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\
        );

    \I__2497\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__20604\,
            I => \pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0\
        );

    \I__2495\ : InMux
    port map (
            O => \N__20601\,
            I => \pid_alt.un1_pid_prereg_0_cry_0\
        );

    \I__2494\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__20595\,
            I => \N__20592\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__20592\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2\
        );

    \I__2491\ : InMux
    port map (
            O => \N__20589\,
            I => \pid_alt.un1_pid_prereg_0_cry_1\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__20586\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__20583\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_\
        );

    \I__2488\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__20577\,
            I => \dron_frame_decoder_1.N_188_4\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__20574\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__20571\,
            I => \dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__20568\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\
        );

    \I__2483\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20562\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20562\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_1\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__20559\,
            I => \N__20556\
        );

    \I__2480\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20552\
        );

    \I__2479\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20549\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__20552\,
            I => \N__20546\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__20549\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__20546\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__20541\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_\
        );

    \I__2474\ : InMux
    port map (
            O => \N__20538\,
            I => \dron_frame_decoder_1.un1_WDT_cry_11\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__20535\,
            I => \N__20532\
        );

    \I__2472\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20528\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__20531\,
            I => \N__20524\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20520\
        );

    \I__2469\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20515\
        );

    \I__2468\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20515\
        );

    \I__2467\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20512\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20507\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20507\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__20512\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__20507\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__2462\ : InMux
    port map (
            O => \N__20502\,
            I => \dron_frame_decoder_1.un1_WDT_cry_12\
        );

    \I__2461\ : InMux
    port map (
            O => \N__20499\,
            I => \N__20496\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20491\
        );

    \I__2459\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20488\
        );

    \I__2458\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20485\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__20491\,
            I => \N__20480\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20480\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__20485\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__20480\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__2453\ : InMux
    port map (
            O => \N__20475\,
            I => \dron_frame_decoder_1.un1_WDT_cry_13\
        );

    \I__2452\ : InMux
    port map (
            O => \N__20472\,
            I => \dron_frame_decoder_1.un1_WDT_cry_14\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__20469\,
            I => \N__20466\
        );

    \I__2450\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20462\
        );

    \I__2449\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20459\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__20462\,
            I => \N__20455\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__20459\,
            I => \N__20452\
        );

    \I__2446\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20449\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__20455\,
            I => \N__20444\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__20452\,
            I => \N__20444\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__20449\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__20444\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__20439\,
            I => \N__20435\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20430\
        );

    \I__2439\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20430\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20430\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__20427\,
            I => \N__20424\
        );

    \I__2436\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20418\
        );

    \I__2435\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20418\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__20418\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__20415\,
            I => \dron_frame_decoder_1.N_188_4_cascade_\
        );

    \I__2432\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20409\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__20409\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20399\
        );

    \I__2428\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20396\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__20399\,
            I => \N__20393\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__20396\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__20393\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20388\,
            I => \dron_frame_decoder_1.un1_WDT_cry_3\
        );

    \I__2423\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20378\
        );

    \I__2421\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20375\
        );

    \I__2420\ : Span4Mux_v
    port map (
            O => \N__20378\,
            I => \N__20372\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__20375\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__20372\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20367\,
            I => \dron_frame_decoder_1.un1_WDT_cry_4\
        );

    \I__2416\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20361\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__20361\,
            I => \N__20357\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20354\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__20357\,
            I => \N__20351\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20354\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__20351\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__2410\ : InMux
    port map (
            O => \N__20346\,
            I => \dron_frame_decoder_1.un1_WDT_cry_5\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20340\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20336\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20333\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__20336\,
            I => \N__20330\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__20333\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__20330\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20325\,
            I => \dron_frame_decoder_1.un1_WDT_cry_6\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20318\
        );

    \I__2401\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20315\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20318\,
            I => \N__20312\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__20315\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__20312\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20307\,
            I => \bfn_7_8_0_\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20297\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20294\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20297\,
            I => \N__20291\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__20294\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__20291\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20286\,
            I => \dron_frame_decoder_1.un1_WDT_cry_8\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20279\
        );

    \I__2388\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20276\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20273\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20276\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__20273\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20268\,
            I => \dron_frame_decoder_1.un1_WDT_cry_9\
        );

    \I__2383\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20258\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20258\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20255\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20252\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__20255\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__20252\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__2377\ : InMux
    port map (
            O => \N__20247\,
            I => \dron_frame_decoder_1.un1_WDT_cry_10\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20244\,
            I => \N__20237\
        );

    \I__2375\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__2374\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20234\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20231\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__20234\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__20231\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__20223\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20217\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__20217\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__20214\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_\
        );

    \I__2365\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20208\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__20208\,
            I => \N__20203\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20198\
        );

    \I__2362\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20198\
        );

    \I__2361\ : Span12Mux_s5_h
    port map (
            O => \N__20203\,
            I => \N__20193\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__20198\,
            I => \N__20193\
        );

    \I__2359\ : Span12Mux_v
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2358\ : Odrv12
    port map (
            O => \N__20190\,
            I => \pid_alt.error_d_regZ0Z_23\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20183\
        );

    \I__2356\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20180\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__20183\,
            I => \pid_alt.error_d_reg_prevZ0Z_23\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__20180\,
            I => \pid_alt.error_d_reg_prevZ0Z_23\
        );

    \I__2353\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20169\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__20169\,
            I => \N__20166\
        );

    \I__2350\ : Span4Mux_h
    port map (
            O => \N__20166\,
            I => \N__20163\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__20163\,
            I => \pid_alt.O_1_8\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__20160\,
            I => \N__20156\
        );

    \I__2347\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20153\
        );

    \I__2346\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20150\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__20153\,
            I => \N__20145\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20145\
        );

    \I__2343\ : Span4Mux_h
    port map (
            O => \N__20145\,
            I => \N__20142\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__20142\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__2341\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20136\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__20136\,
            I => \dron_frame_decoder_1.WDTZ0Z_0\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__20130\,
            I => \dron_frame_decoder_1.WDTZ0Z_1\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20127\,
            I => \dron_frame_decoder_1.un1_WDT_cry_0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__20121\,
            I => \dron_frame_decoder_1.WDTZ0Z_2\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20118\,
            I => \dron_frame_decoder_1.un1_WDT_cry_1\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20115\,
            I => \N__20112\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__20112\,
            I => \dron_frame_decoder_1.WDTZ0Z_3\
        );

    \I__2331\ : InMux
    port map (
            O => \N__20109\,
            I => \dron_frame_decoder_1.un1_WDT_cry_2\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__20106\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20097\
        );

    \I__2328\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20097\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20097\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20088\
        );

    \I__2325\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20088\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20085\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__20085\,
            I => \N__20082\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__20082\,
            I => \N__20079\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__20079\,
            I => \pid_alt.error_p_regZ0Z_14\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\
        );

    \I__2319\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20064\
        );

    \I__2318\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20064\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20064\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20061\
        );

    \I__2315\ : Span12Mux_s6_h
    port map (
            O => \N__20061\,
            I => \N__20058\
        );

    \I__2314\ : Span12Mux_v
    port map (
            O => \N__20058\,
            I => \N__20055\
        );

    \I__2313\ : Odrv12
    port map (
            O => \N__20055\,
            I => \pid_alt.error_d_regZ0Z_14\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__2311\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20043\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20048\,
            I => \N__20043\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__20043\,
            I => \pid_alt.error_d_reg_prevZ0Z_14\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20034\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20034\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__2305\ : Span4Mux_h
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__20028\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__20022\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__20019\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20012\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20015\,
            I => \N__20009\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__20012\,
            I => \pid_alt.error_d_reg_prevZ0Z_22\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__20009\,
            I => \pid_alt.error_d_reg_prevZ0Z_22\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19998\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19998\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19994\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19991\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__19994\,
            I => \N__19986\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19986\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__19977\,
            I => \pid_alt.error_d_regZ0Z_22\
        );

    \I__2286\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19968\
        );

    \I__2285\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19968\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__19968\,
            I => \N__19965\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__19962\,
            I => \pid_alt.error_p_regZ0Z_7\
        );

    \I__2281\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19953\
        );

    \I__2280\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19953\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__19953\,
            I => \pid_alt.error_d_reg_prevZ0Z_7\
        );

    \I__2278\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19941\
        );

    \I__2277\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19941\
        );

    \I__2276\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19941\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__19932\,
            I => \pid_alt.error_d_regZ0Z_7\
        );

    \I__2271\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19925\
        );

    \I__2270\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19922\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19919\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19916\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__19919\,
            I => \N__19913\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__19916\,
            I => \N__19910\
        );

    \I__2265\ : Odrv4
    port map (
            O => \N__19913\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__19910\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__2263\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19898\
        );

    \I__2262\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19898\
        );

    \I__2261\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19895\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19890\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__19895\,
            I => \N__19890\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__19890\,
            I => \N__19887\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__19884\,
            I => \pid_alt.error_d_regZ0Z_8\
        );

    \I__2255\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19877\
        );

    \I__2254\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19874\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__19877\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__19874\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19863\
        );

    \I__2250\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19863\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19860\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__19860\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\
        );

    \I__2247\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__19854\,
            I => \pid_alt.error_d_reg_prevZ0Z_0\
        );

    \I__2245\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19847\
        );

    \I__2244\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19844\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__19847\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__19844\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__2241\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19835\
        );

    \I__2240\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19832\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19827\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19827\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__19821\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__2234\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19813\
        );

    \I__2233\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19810\
        );

    \I__2232\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19807\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__19813\,
            I => \N__19800\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19800\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19800\
        );

    \I__2228\ : Span12Mux_v
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__19797\,
            I => \pid_alt.error_d_regZ0Z_15\
        );

    \I__2226\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19791\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19791\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__19788\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_\
        );

    \I__2223\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19779\
        );

    \I__2222\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19779\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__19779\,
            I => \N__19776\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__19770\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__2216\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19758\
        );

    \I__2215\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19758\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__19758\,
            I => \pid_alt.error_d_reg_prevZ0Z_16\
        );

    \I__2213\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19746\
        );

    \I__2212\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19746\
        );

    \I__2211\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19746\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__2207\ : Span4Mux_h
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__19734\,
            I => \pid_alt.error_d_regZ0Z_16\
        );

    \I__2205\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19728\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__19728\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__19725\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_\
        );

    \I__2201\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__19716\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\
        );

    \I__2199\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__19710\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__19707\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\
        );

    \I__2196\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19698\
        );

    \I__2195\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19698\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__19695\,
            I => \N__19692\
        );

    \I__2192\ : Span4Mux_v
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__19689\,
            I => \pid_alt.error_p_regZ0Z_11\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__2189\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19677\
        );

    \I__2188\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19677\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__19677\,
            I => \pid_alt.error_d_reg_prevZ0Z_11\
        );

    \I__2186\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19665\
        );

    \I__2185\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19665\
        );

    \I__2184\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19665\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__19665\,
            I => \N__19661\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__19664\,
            I => \N__19658\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__2180\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19652\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__19655\,
            I => \N__19649\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__19652\,
            I => \pid_alt.error_d_regZ0Z_11\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__19649\,
            I => \pid_alt.error_d_regZ0Z_11\
        );

    \I__2176\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19641\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__19641\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11\
        );

    \I__2174\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19632\
        );

    \I__2173\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19632\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__19632\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__19620\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\
        );

    \I__2167\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__19614\,
            I => \N__19610\
        );

    \I__2165\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19607\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__19610\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__19607\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__19602\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_\
        );

    \I__2161\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__19596\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\
        );

    \I__2159\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19587\
        );

    \I__2158\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19587\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__2156\ : Span12Mux_h
    port map (
            O => \N__19584\,
            I => \N__19581\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__19581\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__19578\,
            I => \dron_frame_decoder_1.WDT10lto9_3_cascade_\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__19575\,
            I => \dron_frame_decoder_1.WDT10lt12_0_cascade_\
        );

    \I__2152\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19569\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__19569\,
            I => \dron_frame_decoder_1.WDT10_0_i_1\
        );

    \I__2150\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__19563\,
            I => \dron_frame_decoder_1.WDT10lt12_0\
        );

    \I__2148\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__19557\,
            I => \dron_frame_decoder_1.WDT10lt14_0\
        );

    \I__2146\ : CEMux
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__19551\,
            I => \pid_alt.state_1_0_0\
        );

    \I__2144\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19542\
        );

    \I__2143\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19542\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__19536\,
            I => \pid_alt.error_p_regZ0Z_12\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19527\
        );

    \I__2138\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19527\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__19527\,
            I => \pid_alt.error_d_reg_prevZ0Z_12\
        );

    \I__2136\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19515\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19515\
        );

    \I__2134\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19515\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__2131\ : Sp12to4
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__2130\ : Odrv12
    port map (
            O => \N__19506\,
            I => \pid_alt.error_d_regZ0Z_12\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\
        );

    \I__2128\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19495\
        );

    \I__2127\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19490\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19490\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19495\,
            I => \N__19485\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__19490\,
            I => \N__19485\
        );

    \I__2123\ : Span4Mux_h
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__2122\ : Sp12to4
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__19479\,
            I => \pid_alt.error_d_regZ0Z_13\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19476\,
            I => \N__19472\
        );

    \I__2119\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19469\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__19472\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19469\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2116\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__19458\,
            I => \N__19455\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__19455\,
            I => \pid_alt.O_0_15\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19446\
        );

    \I__2111\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19446\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__19446\,
            I => \N__19443\
        );

    \I__2109\ : Span4Mux_h
    port map (
            O => \N__19443\,
            I => \N__19440\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__19440\,
            I => \N__19437\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__19437\,
            I => \pid_alt.error_p_regZ0Z_18\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__19434\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\
        );

    \I__2105\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19422\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19422\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19422\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__19422\,
            I => \N__19419\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__19413\,
            I => \N__19410\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__19410\,
            I => \pid_alt.error_d_regZ0Z_18\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__2096\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19398\
        );

    \I__2095\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19398\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__19398\,
            I => \pid_alt.error_d_reg_prevZ0Z_18\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__19392\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19383\
        );

    \I__2090\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19383\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19380\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__19374\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19367\
        );

    \I__2084\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19364\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__19367\,
            I => \N__19359\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19359\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__19359\,
            I => \N__19356\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__19356\,
            I => \N__19353\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__19353\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__19350\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_\
        );

    \I__2077\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19344\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\
        );

    \I__2075\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__19338\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\
        );

    \I__2072\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__19329\,
            I => \pid_alt.g0_4_0\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19321\
        );

    \I__2069\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19318\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__19324\,
            I => \N__19314\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19308\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__19318\,
            I => \N__19308\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19305\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19300\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19300\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__19308\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__19305\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19300\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19293\,
            I => \N__19289\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19286\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19278\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19278\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19275\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19270\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19270\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__19278\,
            I => \N__19267\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19262\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19262\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__19267\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__2048\ : Odrv12
    port map (
            O => \N__19262\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19253\
        );

    \I__2046\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19250\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19242\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19242\
        );

    \I__2043\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19238\
        );

    \I__2042\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19233\
        );

    \I__2041\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19233\
        );

    \I__2040\ : Span4Mux_h
    port map (
            O => \N__19242\,
            I => \N__19230\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19227\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__19238\,
            I => \N__19222\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19222\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__19230\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19227\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__19222\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__2033\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__19212\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__19209\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__19203\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19193\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19193\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19190\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19193\,
            I => \N__19187\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19184\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__19187\,
            I => \N__19181\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__19184\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__19181\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__2020\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19169\
        );

    \I__2019\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19169\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19166\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19169\,
            I => \N__19163\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__19166\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__19163\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19152\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19149\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19144\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19144\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__19152\,
            I => \N__19141\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19149\,
            I => \N__19138\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__19144\,
            I => \N__19135\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__19141\,
            I => \N__19130\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__19138\,
            I => \N__19130\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__19135\,
            I => \N__19127\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__19130\,
            I => \pid_alt.error_d_regZ0Z_3\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__19127\,
            I => \pid_alt.error_d_regZ0Z_3\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19119\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19119\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\
        );

    \I__2000\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19110\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19110\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__19107\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__19104\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19097\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19094\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__19097\,
            I => \pid_alt.error_d_reg_prevZ0Z_20\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__19094\,
            I => \pid_alt.error_d_reg_prevZ0Z_20\
        );

    \I__1991\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19083\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19083\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__19083\,
            I => \N__19079\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19076\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__19079\,
            I => \N__19073\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19070\
        );

    \I__1985\ : Sp12to4
    port map (
            O => \N__19073\,
            I => \N__19065\
        );

    \I__1984\ : Span12Mux_h
    port map (
            O => \N__19070\,
            I => \N__19065\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__19065\,
            I => \pid_alt.error_d_regZ0Z_20\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__19059\,
            I => \N__19056\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__19056\,
            I => \N__19053\
        );

    \I__1979\ : Span4Mux_v
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__19050\,
            I => \pid_alt.O_1_7\
        );

    \I__1977\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19041\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__19041\,
            I => \N__19038\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__19038\,
            I => \N__19035\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__19035\,
            I => alt_kp_0
        );

    \I__1972\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19029\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__19029\,
            I => \N__19026\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__19026\,
            I => \N__19023\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__19023\,
            I => alt_kp_6
        );

    \I__1968\ : InMux
    port map (
            O => \N__19020\,
            I => \N__19017\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1966\ : Span4Mux_s3_h
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__19011\,
            I => alt_kp_5
        );

    \I__1964\ : InMux
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__19002\,
            I => \N__18999\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__18999\,
            I => \pid_alt.O_0_16\
        );

    \I__1960\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18993\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__18993\,
            I => \N__18989\
        );

    \I__1958\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18986\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__18989\,
            I => \N__18983\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18980\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__18983\,
            I => \N__18975\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__18980\,
            I => \N__18975\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__18975\,
            I => alt_kd_4
        );

    \I__1952\ : CEMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__18969\,
            I => \N__18966\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__18966\,
            I => \N__18961\
        );

    \I__1949\ : CEMux
    port map (
            O => \N__18965\,
            I => \N__18958\
        );

    \I__1948\ : CEMux
    port map (
            O => \N__18964\,
            I => \N__18955\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__18961\,
            I => \Commands_frame_decoder.source_alt_kd_1_sqmuxa\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__18958\,
            I => \Commands_frame_decoder.source_alt_kd_1_sqmuxa\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__18955\,
            I => \Commands_frame_decoder.source_alt_kd_1_sqmuxa\
        );

    \I__1944\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__18945\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__18942\,
            I => \pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_\
        );

    \I__1941\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18936\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__18936\,
            I => \pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0\
        );

    \I__1939\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__18930\,
            I => \pid_alt.N_1078_0\
        );

    \I__1937\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18924\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__18924\,
            I => \N__18915\
        );

    \I__1935\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18910\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18910\
        );

    \I__1933\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18907\
        );

    \I__1932\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18900\
        );

    \I__1931\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18900\
        );

    \I__1930\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18900\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__18915\,
            I => \N__18895\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__18910\,
            I => \N__18895\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18890\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18890\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__18895\,
            I => \N__18887\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__18890\,
            I => \N__18884\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__18887\,
            I => \pid_alt.error_p_regZ0Z_1\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__18884\,
            I => \pid_alt.error_p_regZ0Z_1\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__18879\,
            I => \N__18875\
        );

    \I__1920\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18869\
        );

    \I__1919\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18864\
        );

    \I__1918\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18864\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18861\
        );

    \I__1916\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18856\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18851\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__18864\,
            I => \N__18851\
        );

    \I__1913\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18844\
        );

    \I__1912\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18844\
        );

    \I__1911\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18844\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__18856\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__18851\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__18844\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1907\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18830\
        );

    \I__1906\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18830\
        );

    \I__1905\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18826\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__18830\,
            I => \N__18823\
        );

    \I__1903\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18818\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__18826\,
            I => \N__18813\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__18823\,
            I => \N__18813\
        );

    \I__1900\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18808\
        );

    \I__1899\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18808\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18818\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__18813\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__18808\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__1895\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18798\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__18798\,
            I => \pid_alt.N_1074_1\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__18795\,
            I => \pid_alt.N_3_1_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__18789\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2\
        );

    \I__1890\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__18780\,
            I => \pid_alt.g1_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__18774\,
            I => \N__18771\
        );

    \I__1885\ : Span4Mux_s3_h
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__18768\,
            I => alt_kp_2
        );

    \I__1883\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18762\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__18762\,
            I => \N__18759\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__18759\,
            I => \N__18756\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__18756\,
            I => \pid_alt.O_0_22\
        );

    \I__1879\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18749\
        );

    \I__1878\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18746\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__18749\,
            I => \N__18743\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__18746\,
            I => \N__18740\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__18743\,
            I => \N__18735\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__18740\,
            I => \N__18735\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__18735\,
            I => alt_kd_6
        );

    \I__1872\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18728\
        );

    \I__1871\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18725\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__18728\,
            I => \N__18722\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__18725\,
            I => \N__18719\
        );

    \I__1868\ : Span4Mux_s3_h
    port map (
            O => \N__18722\,
            I => \N__18716\
        );

    \I__1867\ : Span4Mux_s3_h
    port map (
            O => \N__18719\,
            I => \N__18713\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__18716\,
            I => alt_kd_5
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__18713\,
            I => alt_kd_5
        );

    \I__1864\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__18702\,
            I => \pid_alt.O_4\
        );

    \I__1861\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__18696\,
            I => \pid_alt.N_1074_0\
        );

    \I__1859\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18690\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__18690\,
            I => \pid_alt.N_5_0\
        );

    \I__1857\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18684\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__18684\,
            I => \pid_alt.g1_1\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__18681\,
            I => \pid_alt.N_1080_0_cascade_\
        );

    \I__1854\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18674\
        );

    \I__1853\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18671\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18666\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18666\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__18663\,
            I => \pid_alt.error_d_reg_fastZ0Z_1\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__1847\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18654\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__18654\,
            I => \pid_alt.N_3_0\
        );

    \I__1845\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18646\
        );

    \I__1844\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18641\
        );

    \I__1843\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18641\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18636\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18636\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__18636\,
            I => \N__18633\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__18630\,
            I => \pid_alt.error_d_regZ0Z_19\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__18627\,
            I => \N__18624\
        );

    \I__1836\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18618\
        );

    \I__1835\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18618\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__18618\,
            I => \pid_alt.error_d_reg_prevZ0Z_19\
        );

    \I__1833\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18609\
        );

    \I__1832\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18609\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__18609\,
            I => \N__18606\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__18606\,
            I => \N__18603\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__18603\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__1828\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18597\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__18597\,
            I => \N__18594\
        );

    \I__1826\ : Span12Mux_v
    port map (
            O => \N__18594\,
            I => \N__18591\
        );

    \I__1825\ : Odrv12
    port map (
            O => \N__18591\,
            I => \pid_alt.O_1_6\
        );

    \I__1824\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__18582\,
            I => \N__18579\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__18579\,
            I => \N__18576\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__18576\,
            I => \pid_alt.O_1_5\
        );

    \I__1819\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__1817\ : Span12Mux_v
    port map (
            O => \N__18567\,
            I => \N__18564\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__18564\,
            I => \pid_alt.O_1_14\
        );

    \I__1815\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__1813\ : Span4Mux_s2_h
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__18549\,
            I => alt_kp_3
        );

    \I__1810\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18543\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__18543\,
            I => \N__18540\
        );

    \I__1808\ : Span4Mux_s2_h
    port map (
            O => \N__18540\,
            I => \N__18537\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__18537\,
            I => alt_kp_1
        );

    \I__1806\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__18531\,
            I => \N__18528\
        );

    \I__1804\ : Span4Mux_s2_h
    port map (
            O => \N__18528\,
            I => \N__18525\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__18525\,
            I => alt_kp_7
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__18522\,
            I => \pid_alt.g0_0_0_cascade_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__18519\,
            I => \N__18516\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18513\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__18513\,
            I => \pid_alt.O_0_18\
        );

    \I__1798\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__18507\,
            I => \pid_alt.O_0_19\
        );

    \I__1796\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18497\
        );

    \I__1794\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18494\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__18497\,
            I => \N__18491\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__18494\,
            I => \N__18488\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__18491\,
            I => \N__18485\
        );

    \I__1790\ : Span12Mux_s11_v
    port map (
            O => \N__18488\,
            I => \N__18482\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__18485\,
            I => \N__18479\
        );

    \I__1788\ : Odrv12
    port map (
            O => \N__18482\,
            I => \pid_alt.error_p_regZ0Z_17\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__18479\,
            I => \pid_alt.error_p_regZ0Z_17\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18474\,
            I => \N__18470\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18467\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__18470\,
            I => \pid_alt.error_d_reg_prevZ0Z_17\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__18467\,
            I => \pid_alt.error_d_reg_prevZ0Z_17\
        );

    \I__1782\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18457\
        );

    \I__1781\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18454\
        );

    \I__1780\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18451\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__18457\,
            I => \N__18444\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__18454\,
            I => \N__18444\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18444\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__18444\,
            I => \pid_alt.error_d_regZ0Z_17\
        );

    \I__1775\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18437\
        );

    \I__1774\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18434\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__18437\,
            I => \N__18431\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__18434\,
            I => \N__18428\
        );

    \I__1771\ : Span4Mux_s2_h
    port map (
            O => \N__18431\,
            I => \N__18425\
        );

    \I__1770\ : Span4Mux_s2_h
    port map (
            O => \N__18428\,
            I => \N__18422\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__18425\,
            I => alt_kd_2
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__18422\,
            I => alt_kd_2
        );

    \I__1767\ : InMux
    port map (
            O => \N__18417\,
            I => \N__18413\
        );

    \I__1766\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18410\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18407\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__18410\,
            I => \N__18404\
        );

    \I__1763\ : Span4Mux_s3_h
    port map (
            O => \N__18407\,
            I => \N__18401\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__18404\,
            I => \N__18398\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__18401\,
            I => alt_kd_3
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__18398\,
            I => alt_kd_3
        );

    \I__1759\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18389\
        );

    \I__1758\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18386\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__18389\,
            I => \N__18383\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__18386\,
            I => \N__18380\
        );

    \I__1755\ : Span4Mux_s2_h
    port map (
            O => \N__18383\,
            I => \N__18377\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__18380\,
            I => \N__18374\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__18377\,
            I => alt_kd_7
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__18374\,
            I => alt_kd_7
        );

    \I__1751\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18365\
        );

    \I__1750\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18362\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18359\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__18362\,
            I => \N__18356\
        );

    \I__1747\ : Span12Mux_s9_v
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__1746\ : Span4Mux_s2_h
    port map (
            O => \N__18356\,
            I => \N__18350\
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__18353\,
            I => alt_kd_1
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__18350\,
            I => alt_kd_1
        );

    \I__1743\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18338\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18335\
        );

    \I__1740\ : Span4Mux_s1_h
    port map (
            O => \N__18338\,
            I => \N__18332\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__18335\,
            I => \N__18329\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__18332\,
            I => \N__18326\
        );

    \I__1737\ : Span4Mux_s2_h
    port map (
            O => \N__18329\,
            I => \N__18323\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__18326\,
            I => alt_kd_0
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__18323\,
            I => alt_kd_0
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__18318\,
            I => \N__18311\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18307\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__18316\,
            I => \N__18303\
        );

    \I__1731\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18288\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18288\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18288\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18288\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18288\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18288\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18288\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18288\,
            I => \pid_alt.O_1_21\
        );

    \I__1723\ : InMux
    port map (
            O => \N__18285\,
            I => \pid_alt.error_filt_cry_21\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18279\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__18279\,
            I => \N__18276\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__18273\,
            I => \pid_alt.O_1_11\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18267\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__18267\,
            I => \N__18264\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__18264\,
            I => \N__18261\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__18261\,
            I => \pid_alt.O_1_12\
        );

    \I__1714\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18255\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__18252\,
            I => \pid_alt.O_1_10\
        );

    \I__1711\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18246\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__1709\ : Span4Mux_h
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18240\,
            I => \pid_alt.O_0_17\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18234\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18231\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__18231\,
            I => \pid_alt.O_0_20\
        );

    \I__1704\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__18222\,
            I => \N__18219\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__18219\,
            I => \pid_alt.O_0_23\
        );

    \I__1700\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18213\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__18210\,
            I => \pid_alt.O_1_13\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18207\,
            I => \N__18204\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__18204\,
            I => \N__18201\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__18201\,
            I => \pid_alt.O_0_21\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18192\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__18192\,
            I => \pid_alt.O_0_24\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18186\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__18186\,
            I => \pid_alt.O_1_19\
        );

    \I__1689\ : InMux
    port map (
            O => \N__18183\,
            I => \pid_alt.error_filt_cry_13\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__18180\,
            I => \N__18177\
        );

    \I__1687\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18174\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18174\,
            I => \pid_alt.O_1_20\
        );

    \I__1685\ : InMux
    port map (
            O => \N__18171\,
            I => \pid_alt.error_filt_cry_14\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18168\,
            I => \bfn_1_18_0_\
        );

    \I__1683\ : InMux
    port map (
            O => \N__18165\,
            I => \pid_alt.error_filt_cry_16\
        );

    \I__1682\ : InMux
    port map (
            O => \N__18162\,
            I => \pid_alt.error_filt_cry_17\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18159\,
            I => \pid_alt.error_filt_cry_18\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18156\,
            I => \pid_alt.error_filt_cry_19\
        );

    \I__1679\ : InMux
    port map (
            O => \N__18153\,
            I => \pid_alt.error_filt_cry_20\
        );

    \I__1678\ : InMux
    port map (
            O => \N__18150\,
            I => \pid_alt.error_filt_cry_4\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__1675\ : Span4Mux_s2_h
    port map (
            O => \N__18141\,
            I => \N__18138\
        );

    \I__1674\ : Span4Mux_h
    port map (
            O => \N__18138\,
            I => \N__18135\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__18135\,
            I => \N__18132\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__18129\,
            I => \N__18126\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__18126\,
            I => \N__18123\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__18123\,
            I => \pid_alt.O_3_11\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__18120\,
            I => \N__18117\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__18114\,
            I => \pid_alt.O_2_11\
        );

    \I__1665\ : InMux
    port map (
            O => \N__18111\,
            I => \pid_alt.error_filt_cry_5\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__18105\,
            I => \pid_alt.O_2_12\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__18102\,
            I => \N__18099\
        );

    \I__1661\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18096\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18093\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__1658\ : Sp12to4
    port map (
            O => \N__18090\,
            I => \N__18087\
        );

    \I__1657\ : Span12Mux_h
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__1656\ : Odrv12
    port map (
            O => \N__18084\,
            I => \pid_alt.O_3_12\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18081\,
            I => \pid_alt.error_filt_cry_6\
        );

    \I__1654\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18075\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__1652\ : Span12Mux_v
    port map (
            O => \N__18072\,
            I => \N__18069\
        );

    \I__1651\ : Span12Mux_h
    port map (
            O => \N__18069\,
            I => \N__18066\
        );

    \I__1650\ : Span12Mux_h
    port map (
            O => \N__18066\,
            I => \N__18063\
        );

    \I__1649\ : Odrv12
    port map (
            O => \N__18063\,
            I => \pid_alt.O_3_13\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__18060\,
            I => \N__18057\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18054\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__18054\,
            I => \pid_alt.O_2_13\
        );

    \I__1645\ : InMux
    port map (
            O => \N__18051\,
            I => \bfn_1_17_0_\
        );

    \I__1644\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18045\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__18042\,
            I => \N__18039\
        );

    \I__1641\ : Sp12to4
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__1640\ : Span12Mux_h
    port map (
            O => \N__18036\,
            I => \N__18033\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__18033\,
            I => \pid_alt.O_3_14\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__18030\,
            I => \N__18027\
        );

    \I__1637\ : InMux
    port map (
            O => \N__18027\,
            I => \N__18024\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__18024\,
            I => \pid_alt.O_2_14\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18021\,
            I => \pid_alt.error_filt_cry_8\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__18018\,
            I => \N__18015\
        );

    \I__1633\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18012\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__18012\,
            I => \pid_alt.O_1_15\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18009\,
            I => \pid_alt.error_filt_cry_9\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__18006\,
            I => \N__18003\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18003\,
            I => \N__18000\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__18000\,
            I => \pid_alt.O_1_16\
        );

    \I__1627\ : InMux
    port map (
            O => \N__17997\,
            I => \pid_alt.error_filt_cry_10\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__17994\,
            I => \N__17991\
        );

    \I__1625\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17988\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__17988\,
            I => \pid_alt.O_1_17\
        );

    \I__1623\ : InMux
    port map (
            O => \N__17985\,
            I => \pid_alt.error_filt_cry_11\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__1621\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17976\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__17976\,
            I => \pid_alt.O_1_18\
        );

    \I__1619\ : InMux
    port map (
            O => \N__17973\,
            I => \pid_alt.error_filt_cry_12\
        );

    \I__1618\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__1616\ : Span12Mux_h
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__1615\ : Odrv12
    port map (
            O => \N__17961\,
            I => \pid_alt.O_1_4\
        );

    \I__1614\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17955\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__17955\,
            I => \N__17952\
        );

    \I__1612\ : Span4Mux_s3_h
    port map (
            O => \N__17952\,
            I => \N__17949\
        );

    \I__1611\ : Span4Mux_h
    port map (
            O => \N__17949\,
            I => \N__17946\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__17946\,
            I => \N__17943\
        );

    \I__1609\ : Span4Mux_h
    port map (
            O => \N__17943\,
            I => \N__17940\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__17940\,
            I => \N__17937\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__17937\,
            I => \N__17934\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__17934\,
            I => \pid_alt.error_filt_prevZ0Z_0\
        );

    \I__1605\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17927\
        );

    \I__1604\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17924\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__17927\,
            I => \N__17921\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__17924\,
            I => \N__17918\
        );

    \I__1601\ : Span12Mux_v
    port map (
            O => \N__17921\,
            I => \N__17915\
        );

    \I__1600\ : Span12Mux_s4_h
    port map (
            O => \N__17918\,
            I => \N__17912\
        );

    \I__1599\ : Span12Mux_h
    port map (
            O => \N__17915\,
            I => \N__17909\
        );

    \I__1598\ : Span12Mux_h
    port map (
            O => \N__17912\,
            I => \N__17906\
        );

    \I__1597\ : Span12Mux_h
    port map (
            O => \N__17909\,
            I => \N__17903\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__17906\,
            I => \pid_alt.error_filt\
        );

    \I__1595\ : Odrv12
    port map (
            O => \N__17903\,
            I => \pid_alt.error_filt\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__17898\,
            I => \N__17894\
        );

    \I__1593\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17891\
        );

    \I__1592\ : InMux
    port map (
            O => \N__17894\,
            I => \N__17888\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__17891\,
            I => \pid_alt.O_2_5\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__17888\,
            I => \pid_alt.O_2_5\
        );

    \I__1589\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17880\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__17880\,
            I => \N__17877\
        );

    \I__1587\ : Span4Mux_s2_h
    port map (
            O => \N__17877\,
            I => \N__17874\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__17874\,
            I => \pid_alt.error_filt_0\
        );

    \I__1585\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__17868\,
            I => \N__17865\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__1582\ : Sp12to4
    port map (
            O => \N__17862\,
            I => \N__17859\
        );

    \I__1581\ : Span12Mux_h
    port map (
            O => \N__17859\,
            I => \N__17856\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__17856\,
            I => \pid_alt.O_3_6\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__17853\,
            I => \N__17850\
        );

    \I__1578\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17847\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17847\,
            I => \pid_alt.O_2_6\
        );

    \I__1576\ : InMux
    port map (
            O => \N__17844\,
            I => \pid_alt.error_filt_cry_0\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17838\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17835\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__17835\,
            I => \N__17832\
        );

    \I__1572\ : Sp12to4
    port map (
            O => \N__17832\,
            I => \N__17829\
        );

    \I__1571\ : Span12Mux_h
    port map (
            O => \N__17829\,
            I => \N__17826\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__17826\,
            I => \pid_alt.O_3_7\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__17823\,
            I => \N__17820\
        );

    \I__1568\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17817\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__17817\,
            I => \pid_alt.O_2_7\
        );

    \I__1566\ : InMux
    port map (
            O => \N__17814\,
            I => \pid_alt.error_filt_cry_1\
        );

    \I__1565\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17808\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__17808\,
            I => \N__17805\
        );

    \I__1563\ : Span12Mux_s9_h
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__1562\ : Span12Mux_h
    port map (
            O => \N__17802\,
            I => \N__17799\
        );

    \I__1561\ : Odrv12
    port map (
            O => \N__17799\,
            I => \pid_alt.O_3_8\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__17796\,
            I => \N__17793\
        );

    \I__1559\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17790\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__17790\,
            I => \pid_alt.O_2_8\
        );

    \I__1557\ : InMux
    port map (
            O => \N__17787\,
            I => \pid_alt.error_filt_cry_2\
        );

    \I__1556\ : InMux
    port map (
            O => \N__17784\,
            I => \N__17781\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__17781\,
            I => \N__17778\
        );

    \I__1554\ : Span12Mux_v
    port map (
            O => \N__17778\,
            I => \N__17775\
        );

    \I__1553\ : Span12Mux_h
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__17769\,
            I => \pid_alt.O_3_9\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__17766\,
            I => \N__17763\
        );

    \I__1549\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17760\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__17760\,
            I => \pid_alt.O_2_9\
        );

    \I__1547\ : InMux
    port map (
            O => \N__17757\,
            I => \pid_alt.error_filt_cry_3\
        );

    \I__1546\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17751\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__17751\,
            I => \pid_alt.O_2_10\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__17748\,
            I => \N__17745\
        );

    \I__1543\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17742\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__17742\,
            I => \N__17739\
        );

    \I__1541\ : Span12Mux_s7_h
    port map (
            O => \N__17739\,
            I => \N__17736\
        );

    \I__1540\ : Span12Mux_h
    port map (
            O => \N__17736\,
            I => \N__17733\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__17733\,
            I => \pid_alt.O_3_10\
        );

    \I__1538\ : InMux
    port map (
            O => \N__17730\,
            I => \N__17727\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__17727\,
            I => \pid_alt.O_13\
        );

    \I__1536\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__17721\,
            I => \pid_alt.O_11\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__17718\,
            I => \N__17715\
        );

    \I__1533\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17709\
        );

    \I__1532\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17709\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__17709\,
            I => \pid_alt.O_5\
        );

    \I__1530\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17703\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__17703\,
            I => \pid_alt.O_14\
        );

    \I__1528\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17697\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__17697\,
            I => \pid_alt.O_6\
        );

    \I__1526\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17691\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__17691\,
            I => \pid_alt.O_12\
        );

    \I__1524\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17685\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__17685\,
            I => \pid_alt.O_9\
        );

    \I__1522\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17679\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__17679\,
            I => \N__17676\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__17676\,
            I => \pid_alt.O_7\
        );

    \I__1519\ : InMux
    port map (
            O => \N__17673\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_10\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__17670\,
            I => \N__17667\
        );

    \I__1517\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17664\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__17664\,
            I => \pid_alt.un1_error_d_reg_2_12\
        );

    \I__1515\ : InMux
    port map (
            O => \N__17661\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_11\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__17658\,
            I => \N__17655\
        );

    \I__1513\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17652\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__17652\,
            I => \pid_alt.un1_error_d_reg_2_13\
        );

    \I__1511\ : InMux
    port map (
            O => \N__17649\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_12\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__17646\,
            I => \N__17643\
        );

    \I__1509\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17640\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__17640\,
            I => \pid_alt.un1_error_d_reg_2_14\
        );

    \I__1507\ : InMux
    port map (
            O => \N__17637\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_13\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__17634\,
            I => \N__17631\
        );

    \I__1505\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17628\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__17628\,
            I => \pid_alt.un1_error_d_reg_2_15\
        );

    \I__1503\ : InMux
    port map (
            O => \N__17625\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_14\
        );

    \I__1502\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17612\
        );

    \I__1501\ : InMux
    port map (
            O => \N__17621\,
            I => \N__17605\
        );

    \I__1500\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17605\
        );

    \I__1499\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17605\
        );

    \I__1498\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17596\
        );

    \I__1497\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17596\
        );

    \I__1496\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17596\
        );

    \I__1495\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17596\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17591\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__17605\,
            I => \N__17591\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__17596\,
            I => \N__17588\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__17591\,
            I => \N__17585\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__17588\,
            I => \N__17582\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__17585\,
            I => \pid_alt.un1_error_d_reg_1_24\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__17582\,
            I => \pid_alt.un1_error_d_reg_1_24\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__1486\ : InMux
    port map (
            O => \N__17574\,
            I => \N__17571\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__17571\,
            I => \pid_alt.un1_error_d_reg_2_16\
        );

    \I__1484\ : InMux
    port map (
            O => \N__17568\,
            I => \bfn_1_8_0_\
        );

    \I__1483\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17562\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__17562\,
            I => \N__17559\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__17559\,
            I => \pid_alt.O_10\
        );

    \I__1480\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17553\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__17553\,
            I => \N__17550\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__17550\,
            I => \N__17546\
        );

    \I__1477\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17543\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__17546\,
            I => \pid_alt.un1_error_d_reg_2_0\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__17543\,
            I => \pid_alt.un1_error_d_reg_2_0\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__17538\,
            I => \N__17535\
        );

    \I__1473\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17531\
        );

    \I__1472\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17528\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__17531\,
            I => \N__17525\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17520\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__17525\,
            I => \N__17520\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__17520\,
            I => \pid_alt.un1_error_d_reg_1_15\
        );

    \I__1467\ : InMux
    port map (
            O => \N__17517\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_2\
        );

    \I__1466\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17511\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17508\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__17508\,
            I => \pid_alt.un1_error_d_reg_2_4\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__17505\,
            I => \N__17502\
        );

    \I__1462\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17499\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__17499\,
            I => \N__17496\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__17496\,
            I => \N__17493\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__17493\,
            I => \pid_alt.un1_error_d_reg_1_19\
        );

    \I__1458\ : InMux
    port map (
            O => \N__17490\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_3\
        );

    \I__1457\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17484\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__17484\,
            I => \pid_alt.un1_error_d_reg_2_5\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__1454\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17472\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__17469\,
            I => \pid_alt.un1_error_d_reg_1_20\
        );

    \I__1450\ : InMux
    port map (
            O => \N__17466\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_4\
        );

    \I__1449\ : InMux
    port map (
            O => \N__17463\,
            I => \N__17460\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__17460\,
            I => \pid_alt.un1_error_d_reg_2_6\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__1446\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17451\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__17451\,
            I => \N__17448\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__17448\,
            I => \N__17445\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__17445\,
            I => \pid_alt.un1_error_d_reg_1_21\
        );

    \I__1442\ : InMux
    port map (
            O => \N__17442\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_5\
        );

    \I__1441\ : InMux
    port map (
            O => \N__17439\,
            I => \N__17436\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__17436\,
            I => \N__17433\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__17430\,
            I => \pid_alt.un1_error_d_reg_1_22\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__1436\ : InMux
    port map (
            O => \N__17424\,
            I => \N__17421\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__17421\,
            I => \pid_alt.un1_error_d_reg_2_7\
        );

    \I__1434\ : InMux
    port map (
            O => \N__17418\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_6\
        );

    \I__1433\ : InMux
    port map (
            O => \N__17415\,
            I => \N__17412\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__17412\,
            I => \N__17409\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__17409\,
            I => \N__17406\
        );

    \I__1430\ : Span4Mux_s1_h
    port map (
            O => \N__17406\,
            I => \N__17403\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__17403\,
            I => \pid_alt.un1_error_d_reg_1_23\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__17400\,
            I => \N__17397\
        );

    \I__1427\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17394\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__17394\,
            I => \pid_alt.un1_error_d_reg_2_8\
        );

    \I__1425\ : InMux
    port map (
            O => \N__17391\,
            I => \bfn_1_7_0_\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__17388\,
            I => \N__17385\
        );

    \I__1423\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17382\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__17382\,
            I => \pid_alt.un1_error_d_reg_2_9\
        );

    \I__1421\ : InMux
    port map (
            O => \N__17379\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_8\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__17376\,
            I => \N__17373\
        );

    \I__1419\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17370\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__17370\,
            I => \pid_alt.un1_error_d_reg_2_10\
        );

    \I__1417\ : InMux
    port map (
            O => \N__17367\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_9\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__17364\,
            I => \N__17361\
        );

    \I__1415\ : InMux
    port map (
            O => \N__17361\,
            I => \N__17358\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__17358\,
            I => \pid_alt.un1_error_d_reg_2_11\
        );

    \I__1413\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17352\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__17352\,
            I => \pid_alt.un1_error_d_reg_2_1\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__17349\,
            I => \N__17346\
        );

    \I__1410\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17340\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__17340\,
            I => \N__17337\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__17337\,
            I => \pid_alt.un1_error_d_reg_1_16\
        );

    \I__1406\ : InMux
    port map (
            O => \N__17334\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_0\
        );

    \I__1405\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17328\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__17328\,
            I => \pid_alt.un1_error_d_reg_2_2\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__17325\,
            I => \N__17322\
        );

    \I__1402\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17316\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__17313\,
            I => \pid_alt.un1_error_d_reg_1_17\
        );

    \I__1398\ : InMux
    port map (
            O => \N__17310\,
            I => \pid_alt.un1_error_d_reg_add_1_cry_1\
        );

    \I__1397\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17304\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__17301\,
            I => \pid_alt.un1_error_d_reg_2_3\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__17298\,
            I => \N__17295\
        );

    \I__1393\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17292\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__17292\,
            I => \N__17289\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__17286\,
            I => \pid_alt.un1_error_d_reg_1_18\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_6\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_14\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_22\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un3_source_data_0_cry_7\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un2_source_data_0_cry_8\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un3_source_data_0_cry_7\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un2_source_data_0_cry_8\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_13\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_13\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un9lto29_i_a2_6\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_d_reg_add_1_cry_7\,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_d_reg_add_1_cry_15\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_cry_7\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un9_error_filt_add_1_cry_7\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_filt_cry_7\,
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_filt_cry_15\,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \dron_frame_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Commands_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_9_6_0_\
        );

    \reset_module_System.reset_RNITC69_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__43371\,
            GLOBALBUFFEROUTPUT => \N_411_g\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32938\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pid_alt.state_RNICP2N1_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22293\,
            GLOBALBUFFEROUTPUT => \pid_alt.N_410_0_g\
        );

    \debug_CH3_20A_c_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30507\,
            GLOBALBUFFEROUTPUT => \debug_CH3_20A_c_0_g\
        );

    \pid_alt.state_RNIH1EN_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24912\,
            GLOBALBUFFEROUTPUT => \pid_alt.state_0_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32886\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_322_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pid_alt.un1_error_d_reg_add_1_cry_0_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17549\,
            in2 => \N__17538\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_12_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17355\,
            in2 => \N__17349\,
            in3 => \N__17334\,
            lcout => \pid_alt.error_d_regZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_0\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_1\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_13_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17331\,
            in2 => \N__17325\,
            in3 => \N__17310\,
            lcout => \pid_alt.error_d_regZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_1\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_2\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_14_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17307\,
            in2 => \N__17298\,
            in3 => \N__17517\,
            lcout => \pid_alt.error_d_regZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_2\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_3\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_15_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17514\,
            in2 => \N__17505\,
            in3 => \N__17490\,
            lcout => \pid_alt.error_d_regZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_3\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_4\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_16_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17487\,
            in2 => \N__17481\,
            in3 => \N__17466\,
            lcout => \pid_alt.error_d_regZ0Z_16\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_4\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_5\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_17_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17463\,
            in2 => \N__17457\,
            in3 => \N__17442\,
            lcout => \pid_alt.error_d_regZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_5\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_6\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_18_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17439\,
            in2 => \N__17427\,
            in3 => \N__17418\,
            lcout => \pid_alt.error_d_regZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_6\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_7\,
            clk => \N__47478\,
            ce => \N__46815\,
            sr => \N__46628\
        );

    \pid_alt.error_d_reg_esr_19_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17415\,
            in2 => \N__17400\,
            in3 => \N__17391\,
            lcout => \pid_alt.error_d_regZ0Z_19\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_8\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_20_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17615\,
            in2 => \N__17388\,
            in3 => \N__17379\,
            lcout => \pid_alt.error_d_regZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_8\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_9\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_21_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17619\,
            in2 => \N__17376\,
            in3 => \N__17367\,
            lcout => \pid_alt.error_d_regZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_9\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_10\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_22_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17616\,
            in2 => \N__17364\,
            in3 => \N__17673\,
            lcout => \pid_alt.error_d_regZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_10\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_11\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_23_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17620\,
            in2 => \N__17670\,
            in3 => \N__17661\,
            lcout => \pid_alt.error_d_regZ0Z_23\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_11\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_12\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_24_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17617\,
            in2 => \N__17658\,
            in3 => \N__17649\,
            lcout => \pid_alt.error_d_regZ0Z_24\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_12\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_13\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_25_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17621\,
            in2 => \N__17646\,
            in3 => \N__17637\,
            lcout => \pid_alt.error_d_regZ0Z_25\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_13\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_14\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_26_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17618\,
            in2 => \N__17634\,
            in3 => \N__17625\,
            lcout => \pid_alt.error_d_regZ0Z_26\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_d_reg_add_1_cry_14\,
            carryout => \pid_alt.un1_error_d_reg_add_1_cry_15\,
            clk => \N__47477\,
            ce => \N__46814\,
            sr => \N__46627\
        );

    \pid_alt.error_d_reg_esr_27_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17622\,
            in2 => \N__17577\,
            in3 => \N__17568\,
            lcout => \pid_alt.error_d_regZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47476\,
            ce => \N__46812\,
            sr => \N__46626\
        );

    \pid_alt.error_d_reg_esr_6_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17565\,
            lcout => \pid_alt.error_d_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47476\,
            ce => \N__46812\,
            sr => \N__46626\
        );

    \pid_alt.error_d_reg_11_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__24128\,
            in1 => \N__17556\,
            in2 => \N__19664\,
            in3 => \N__17534\,
            lcout => \pid_alt.error_d_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47472\,
            ce => 'H',
            sr => \N__46625\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18474\,
            in2 => \_gnd_net_\,
            in3 => \N__18461\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17730\,
            lcout => \pid_alt.error_d_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__46809\,
            sr => \N__46624\
        );

    \pid_alt.error_d_reg_esr_7_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17724\,
            lcout => \pid_alt.error_d_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__46809\,
            sr => \N__46624\
        );

    \pid_alt.error_d_reg_esr_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17714\,
            lcout => \pid_alt.error_d_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_fast_esr_1_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17718\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_esr_10_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17706\,
            lcout => \pid_alt.error_d_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_esr_2_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17700\,
            lcout => \pid_alt.error_d_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_esr_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17694\,
            lcout => \pid_alt.error_d_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_esr_5_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17688\,
            lcout => \pid_alt.error_d_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47464\,
            ce => \N__46805\,
            sr => \N__46623\
        );

    \pid_alt.error_d_reg_esr_3_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17682\,
            lcout => \pid_alt.error_d_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47459\,
            ce => \N__46801\,
            sr => \N__46621\
        );

    \pid_alt.error_d_reg_prev_esr_2_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19249\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => \N__33622\,
            sr => \N__43831\
        );

    \pid_alt.error_p_reg_esr_0_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17970\,
            lcout => \pid_alt.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47438\,
            ce => \N__46800\,
            sr => \N__46620\
        );

    \pid_alt.error_filt_prev_esr_0_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17930\,
            in2 => \_gnd_net_\,
            in3 => \N__17897\,
            lcout => \pid_alt.error_filt_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47438\,
            ce => \N__46800\,
            sr => \N__46620\
        );

    \pid_alt.error_filt_error_filt_axb_0_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17931\,
            in2 => \N__17898\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_filt_0\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \pid_alt.error_filt_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_0_c_RNIBLFT_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17871\,
            in2 => \N__17853\,
            in3 => \N__17844\,
            lcout => \pid_alt.error_filt_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_0\,
            carryout => \pid_alt.error_filt_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_1_c_RNICNGT_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17841\,
            in2 => \N__17823\,
            in3 => \N__17814\,
            lcout => \pid_alt.error_filt_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_1\,
            carryout => \pid_alt.error_filt_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_2_c_RNIDPHT_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17811\,
            in2 => \N__17796\,
            in3 => \N__17787\,
            lcout => \pid_alt.error_filt_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_2\,
            carryout => \pid_alt.error_filt_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_3_c_RNIERIT_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17784\,
            in2 => \N__17766\,
            in3 => \N__17757\,
            lcout => \pid_alt.error_filt_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_3\,
            carryout => \pid_alt.error_filt_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_4_c_RNIFTJT_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17754\,
            in2 => \N__17748\,
            in3 => \N__18150\,
            lcout => \pid_alt.error_filt_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_4\,
            carryout => \pid_alt.error_filt_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_5_c_RNIGVKT_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18147\,
            in2 => \N__18120\,
            in3 => \N__18111\,
            lcout => \pid_alt.error_filt_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_5\,
            carryout => \pid_alt.error_filt_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_6_c_RNIH1MT_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18108\,
            in2 => \N__18102\,
            in3 => \N__18081\,
            lcout => \pid_alt.error_filt_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_6\,
            carryout => \pid_alt.error_filt_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_7_c_RNII3NT_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18078\,
            in2 => \N__18060\,
            in3 => \N__18051\,
            lcout => \pid_alt.error_filt_8\,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => \pid_alt.error_filt_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_8_c_RNIJ5OT_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18048\,
            in2 => \N__18030\,
            in3 => \N__18021\,
            lcout => \pid_alt.error_filt_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_8\,
            carryout => \pid_alt.error_filt_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_axb_0_RNIRHEM_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38310\,
            in2 => \N__18018\,
            in3 => \N__18009\,
            lcout => \pid_alt.error_filt_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_9\,
            carryout => \pid_alt.error_filt_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_1_s_RNI9PB01_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38250\,
            in2 => \N__18006\,
            in3 => \N__17997\,
            lcout => \pid_alt.error_filt_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_10\,
            carryout => \pid_alt.error_filt_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_2_s_RNIBTD01_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38739\,
            in2 => \N__17994\,
            in3 => \N__17985\,
            lcout => \pid_alt.error_filt_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_11\,
            carryout => \pid_alt.error_filt_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_3_s_RNID1G01_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38679\,
            in2 => \N__17982\,
            in3 => \N__17973\,
            lcout => \pid_alt.error_filt_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_12\,
            carryout => \pid_alt.error_filt_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_4_s_RNIF5I01_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18189\,
            in2 => \N__38640\,
            in3 => \N__18183\,
            lcout => \pid_alt.error_filt_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_13\,
            carryout => \pid_alt.error_filt_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_5_s_RNIH9K01_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38604\,
            in2 => \N__18180\,
            in3 => \N__18171\,
            lcout => \pid_alt.error_filt_15\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_14\,
            carryout => \pid_alt.error_filt_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_6_s_RNIJDM01_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38568\,
            in2 => \N__18316\,
            in3 => \N__18168\,
            lcout => \pid_alt.error_filt_16\,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \pid_alt.error_filt_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_7_s_RNILHO01_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18306\,
            in2 => \N__38526\,
            in3 => \N__18165\,
            lcout => \pid_alt.error_filt_17\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_16\,
            carryout => \pid_alt.error_filt_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_8_s_RNINLQ01_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38475\,
            in2 => \N__18317\,
            in3 => \N__18162\,
            lcout => \pid_alt.error_filt_18\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_17\,
            carryout => \pid_alt.error_filt_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_9_s_RNIPPS01_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18310\,
            in2 => \N__39195\,
            in3 => \N__18159\,
            lcout => \pid_alt.error_filt_19\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_18\,
            carryout => \pid_alt.error_filt_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_10_s_RNI20BR_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39156\,
            in2 => \N__18318\,
            in3 => \N__18156\,
            lcout => \pid_alt.error_filt_20\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_19\,
            carryout => \pid_alt.error_filt_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_20_c_RNIEB1O_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18314\,
            in2 => \N__39060\,
            in3 => \N__18153\,
            lcout => \pid_alt.error_filt_21\,
            ltout => OPEN,
            carryin => \pid_alt.error_filt_cry_20\,
            carryout => \pid_alt.error_filt_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_error_filt_cry_21_c_RNIFD2O_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18315\,
            in1 => \N__39059\,
            in2 => \_gnd_net_\,
            in3 => \N__18285\,
            lcout => \pid_alt.error_filt_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_7_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18282\,
            lcout => \pid_alt.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47393\,
            ce => \N__46793\,
            sr => \N__46616\
        );

    \pid_alt.error_p_reg_esr_8_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18270\,
            lcout => \pid_alt.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => \N__46791\,
            sr => \N__46614\
        );

    \pid_alt.error_p_reg_esr_6_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18258\,
            lcout => \pid_alt.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47366\,
            ce => \N__46790\,
            sr => \N__46613\
        );

    \pid_alt.error_p_reg_esr_13_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18249\,
            lcout => \pid_alt.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47366\,
            ce => \N__46790\,
            sr => \N__46613\
        );

    \pid_alt.error_p_reg_esr_16_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18237\,
            lcout => \pid_alt.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => \N__46789\,
            sr => \N__46612\
        );

    \pid_alt.error_p_reg_esr_19_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18228\,
            lcout => \pid_alt.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => \N__46789\,
            sr => \N__46612\
        );

    \pid_alt.error_p_reg_esr_9_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18216\,
            lcout => \pid_alt.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => \N__46789\,
            sr => \N__46612\
        );

    \pid_alt.error_p_reg_esr_17_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18207\,
            lcout => \pid_alt.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__46788\,
            sr => \N__46610\
        );

    \pid_alt.error_p_reg_esr_20_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18198\,
            lcout => \pid_alt.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__46788\,
            sr => \N__46610\
        );

    \pid_alt.error_p_reg_esr_14_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18519\,
            lcout => \pid_alt.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__46788\,
            sr => \N__46610\
        );

    \pid_alt.error_p_reg_esr_15_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18510\,
            lcout => \pid_alt.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47323\,
            ce => \N__46785\,
            sr => \N__46606\
        );

    \pid_alt.error_d_reg_prev_esr_17_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18462\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47474\,
            ce => \N__33599\,
            sr => \N__43803\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18504\,
            in1 => \N__18473\,
            in2 => \_gnd_net_\,
            in3 => \N__18460\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => alt_kd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => \N__18972\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_3_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43353\,
            lcout => alt_kd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => \N__18972\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_7_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45012\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => alt_kd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => \N__18972\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45200\,
            lcout => alt_kd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => \N__18972\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27677\,
            lcout => alt_kd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => \N__18972\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18829\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47461\,
            ce => \N__33610\,
            sr => \N__43814\
        );

    \pid_alt.error_d_reg_esr_RNITF511_1_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__18918\,
            in1 => \N__18859\,
            in2 => \_gnd_net_\,
            in3 => \N__18821\,
            lcout => \pid_alt.N_1074_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20777\,
            lcout => \pid_alt.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_RNITF511_2_1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__18822\,
            in1 => \_gnd_net_\,
            in2 => \N__18873\,
            in3 => \N__18920\,
            lcout => \pid_alt.error_d_reg_esr_RNITF511_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_fast_esr_RNIA7JS_1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__18860\,
            in1 => \N__18678\,
            in2 => \_gnd_net_\,
            in3 => \N__18919\,
            lcout => \pid_alt.N_1074_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19285\,
            in1 => \N__19317\,
            in2 => \_gnd_net_\,
            in3 => \N__19241\,
            lcout => \pid_alt.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__19248\,
            in1 => \_gnd_net_\,
            in2 => \N__19324\,
            in3 => \N__19284\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19283\,
            in1 => \N__19247\,
            in2 => \_gnd_net_\,
            in3 => \N__19313\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_RNIA37K_1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18835\,
            lcout => OPEN,
            ltout => \pid_alt.g0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIL2AQ1_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000001110"
        )
    port map (
            in0 => \N__20724\,
            in1 => \N__20778\,
            in2 => \N__18522\,
            in3 => \N__18921\,
            lcout => \pid_alt.error_p_reg_esr_RNIL2AQ1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_19_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__33623\,
            sr => \N__43832\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__18614\,
            in1 => \N__18623\,
            in2 => \_gnd_net_\,
            in3 => \N__18649\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__18650\,
            in1 => \_gnd_net_\,
            in2 => \N__18627\,
            in3 => \N__18615\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_2_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18600\,
            lcout => \pid_alt.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47418\,
            ce => \N__46799\,
            sr => \N__46619\
        );

    \pid_alt.error_p_reg_esr_1_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18588\,
            lcout => \pid_alt.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47408\,
            ce => \N__46796\,
            sr => \N__46618\
        );

    \pid_alt.error_p_reg_esr_10_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18573\,
            lcout => \pid_alt.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47380\,
            ce => \N__46792\,
            sr => \N__46615\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43365\,
            in2 => \_gnd_net_\,
            in3 => \N__46689\,
            lcout => alt_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => \N__22472\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_1_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45225\,
            in2 => \_gnd_net_\,
            in3 => \N__46688\,
            lcout => alt_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47355\,
            ce => \N__22474\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_6_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45015\,
            in2 => \_gnd_net_\,
            in3 => \N__46687\,
            lcout => alt_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => \N__22482\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36880\,
            in2 => \_gnd_net_\,
            in3 => \N__46686\,
            lcout => alt_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => \N__22482\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_18_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18765\,
            lcout => \pid_alt.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47326\,
            ce => \N__46786\,
            sr => \N__46608\
        );

    \Commands_frame_decoder.source_alt_kd_6_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33439\,
            lcout => alt_kd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47468\,
            ce => \N__18964\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_5_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44240\,
            lcout => alt_kd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47468\,
            ce => \N__18964\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18708\,
            lcout => \pid_alt.error_d_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47462\,
            ce => \N__46804\,
            sr => \N__46622\
        );

    \pid_alt.error_d_reg_fast_esr_RNICKGJ3_1_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100010"
        )
    port map (
            in0 => \N__18699\,
            in1 => \N__18693\,
            in2 => \N__18660\,
            in3 => \N__18687\,
            lcout => OPEN,
            ltout => \pid_alt.N_1080_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIFTRL5_3_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011010100"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__18933\,
            in2 => \N__18681\,
            in3 => \N__19198\,
            lcout => \pid_alt.error_p_reg_esr_RNIFTRL5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_fast_esr_RNIA7JS_0_1_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18677\,
            in1 => \N__18927\,
            in2 => \_gnd_net_\,
            in3 => \N__18872\,
            lcout => \pid_alt.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_RNITF511_0_1_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__18837\,
            in1 => \_gnd_net_\,
            in2 => \N__18879\,
            in3 => \N__18923\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_esr_RNITF511_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF0465_2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__30039\,
            in1 => \N__18948\,
            in2 => \N__18942\,
            in3 => \N__18939\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF0465Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19292\,
            in1 => \N__19325\,
            in2 => \_gnd_net_\,
            in3 => \N__19256\,
            lcout => \pid_alt.N_1078_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_RNITF511_1_1_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18922\,
            in1 => \N__18874\,
            in2 => \_gnd_net_\,
            in3 => \N__18836\,
            lcout => OPEN,
            ltout => \pid_alt.N_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5LS3_2_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__18786\,
            in1 => \N__18801\,
            in2 => \N__18795\,
            in3 => \N__18792\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20782\,
            in2 => \_gnd_net_\,
            in3 => \N__20722\,
            lcout => \pid_alt.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__23174\,
            in2 => \N__21227\,
            in3 => \N__30771\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_20_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => \N__33624\,
            sr => \N__43833\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24634\,
            in1 => \N__19101\,
            in2 => \_gnd_net_\,
            in3 => \N__19088\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19371\,
            in1 => \N__19476\,
            in2 => \_gnd_net_\,
            in3 => \N__19500\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19100\,
            in1 => \N__24608\,
            in2 => \_gnd_net_\,
            in3 => \N__19082\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGGKM_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_3_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19062\,
            lcout => \pid_alt.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__46794\,
            sr => \N__46617\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27681\,
            in2 => \_gnd_net_\,
            in3 => \N__46684\,
            lcout => alt_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47342\,
            ce => \N__22473\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33435\,
            lcout => alt_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47342\,
            ce => \N__22473\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44291\,
            in2 => \_gnd_net_\,
            in3 => \N__46683\,
            lcout => alt_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47327\,
            ce => \N__22481\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_12_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19008\,
            lcout => \pid_alt.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => \N__46783\,
            sr => \N__46605\
        );

    \Commands_frame_decoder.state_RNIRSI31_11_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23709\,
            in1 => \N__27040\,
            in2 => \_gnd_net_\,
            in3 => \N__44092\,
            lcout => \Commands_frame_decoder.source_alt_kd_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_4_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45350\,
            lcout => alt_kd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47455\,
            ce => \N__18965\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_3_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19158\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47447\,
            ce => \N__33602\,
            sr => \N__43808\
        );

    \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19157\,
            lcout => \pid_alt.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19199\,
            in1 => \N__19175\,
            in2 => \_gnd_net_\,
            in3 => \N__19156\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__19326\,
            in1 => \N__19293\,
            in2 => \_gnd_net_\,
            in3 => \N__19257\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__29997\,
            in1 => \N__19215\,
            in2 => \N__19209\,
            in3 => \N__19206\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19200\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__19155\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30138\,
            in1 => \N__20783\,
            in2 => \_gnd_net_\,
            in3 => \N__20734\,
            lcout => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19115\,
            in1 => \N__19122\,
            in2 => \N__20888\,
            in3 => \N__30809\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__19430\,
            in1 => \_gnd_net_\,
            in2 => \N__19407\,
            in3 => \N__19452\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19116\,
            in1 => \_gnd_net_\,
            in2 => \N__19104\,
            in3 => \N__30810\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19451\,
            in1 => \N__19403\,
            in2 => \_gnd_net_\,
            in3 => \N__19429\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19389\,
            in2 => \N__19434\,
            in3 => \N__30846\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_18_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19431\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47409\,
            ce => \N__33620\,
            sr => \N__43824\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19395\,
            in1 => \N__19388\,
            in2 => \N__20930\,
            in3 => \N__30845\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_12_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => \N__33625\,
            sr => \N__43834\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19370\,
            in1 => \N__19475\,
            in2 => \_gnd_net_\,
            in3 => \N__19498\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19347\,
            in2 => \N__19350\,
            in3 => \N__30215\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19548\,
            in1 => \N__19533\,
            in2 => \_gnd_net_\,
            in3 => \N__19523\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIT4AF4_12_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__21119\,
            in1 => \N__19341\,
            in2 => \N__19335\,
            in3 => \N__30214\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIT4AF4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19547\,
            in1 => \N__19532\,
            in2 => \_gnd_net_\,
            in3 => \N__19522\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI1QHB2_11_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19617\,
            in1 => \_gnd_net_\,
            in2 => \N__19503\,
            in3 => \N__30255\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI1QHB2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_13_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19499\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => \N__33625\,
            sr => \N__43834\
        );

    \pid_alt.error_d_reg_prev_esr_0_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20739\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__33628\,
            sr => \N__43840\
        );

    \pid_alt.error_d_reg_prev_esr_RNIKKKM_0_22_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20015\,
            in1 => \N__19997\,
            in2 => \_gnd_net_\,
            in3 => \N__24622\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIKKKM_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMMKM_23_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__20187\,
            in1 => \N__24614\,
            in2 => \_gnd_net_\,
            in3 => \N__20211\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMMKMZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_esr_5_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44292\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => \N__26400\,
            sr => \N__43863\
        );

    \pid_alt.error_p_reg_esr_11_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19464\,
            lcout => \pid_alt.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__46787\,
            sr => \N__46609\
        );

    \dron_frame_decoder_1.WDT_RNIA9RK1_11_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__20243\,
            in1 => \N__20495\,
            in2 => \N__20531\,
            in3 => \N__20264\,
            lcout => \dron_frame_decoder_1.WDT10_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20322\,
            in1 => \N__20385\,
            in2 => \N__20304\,
            in3 => \N__20406\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.WDT10lto9_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI9TKF_6_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__20283\,
            in1 => \N__20343\,
            in2 => \N__19578\,
            in3 => \N__20364\,
            lcout => \dron_frame_decoder_1.WDT10lt12_0\,
            ltout => \dron_frame_decoder_1.WDT10lt12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIBUTU2_15_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101010101"
        )
    port map (
            in0 => \N__20465\,
            in1 => \N__20527\,
            in2 => \N__19575\,
            in3 => \N__19572\,
            lcout => \dron_frame_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNINA9N1_11_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__20265\,
            in1 => \N__20244\,
            in2 => \N__20535\,
            in3 => \N__19566\,
            lcout => \dron_frame_decoder_1.WDT10lt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIPI9R2_15_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__29672\,
            in1 => \N__20499\,
            in2 => \N__20469\,
            in3 => \N__19560\,
            lcout => \dron_frame_decoder_1.WDT_RNIPI9R2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_RNO_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24961\,
            in2 => \_gnd_net_\,
            in3 => \N__44100\,
            lcout => \pid_alt.state_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33229\,
            lcout => pid_altitude_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47430\,
            ce => \N__19554\,
            sr => \N__43809\
        );

    \pid_alt.source_pid_1_4_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__33204\,
            in1 => \N__25914\,
            in2 => \N__29396\,
            in3 => \N__24165\,
            lcout => throttle_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47420\,
            ce => 'H',
            sr => \N__27875\
        );

    \pid_alt.error_d_reg_prev_esr_RNIKQBI4_10_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19637\,
            in1 => \N__19644\,
            in2 => \N__23082\,
            in3 => \N__30299\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIKQBI4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__22946\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI7E8R_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__19673\,
            in1 => \_gnd_net_\,
            in2 => \N__19686\,
            in3 => \N__19704\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI7E8RZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_11_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19674\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47410\,
            ce => \N__33611\,
            sr => \N__43815\
        );

    \pid_alt.error_d_reg_prev_esr_10_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47410\,
            ce => \N__33611\,
            sr => \N__43815\
        );

    \pid_alt.error_d_reg_prev_esr_RNI7E8R_0_11_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19703\,
            in1 => \N__19682\,
            in2 => \_gnd_net_\,
            in3 => \N__19672\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI7E8R_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOFGB2_10_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19638\,
            in1 => \_gnd_net_\,
            in2 => \N__19629\,
            in3 => \N__30300\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIOFGB2Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIP92N4_11_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19626\,
            in1 => \N__19613\,
            in2 => \N__19602\,
            in3 => \N__30250\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIP92N4Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19599\,
            in1 => \N__19593\,
            in2 => \_gnd_net_\,
            in3 => \N__30882\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__19754\,
            in1 => \_gnd_net_\,
            in2 => \N__19767\,
            in3 => \N__19785\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__19592\,
            in2 => \N__19788\,
            in3 => \N__30881\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_16_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19755\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => \N__33615\,
            sr => \N__43819\
        );

    \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19731\,
            in1 => \N__19869\,
            in2 => \_gnd_net_\,
            in3 => \N__30915\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19784\,
            in1 => \N__19763\,
            in2 => \_gnd_net_\,
            in3 => \N__19753\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__21011\,
            in1 => \N__19868\,
            in2 => \N__19725\,
            in3 => \N__30914\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_7_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47382\,
            ce => \N__33621\,
            sr => \N__43825\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__19880\,
            in2 => \_gnd_net_\,
            in3 => \N__19903\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19719\,
            in2 => \N__19722\,
            in3 => \N__30432\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19974\,
            in1 => \N__19959\,
            in2 => \_gnd_net_\,
            in3 => \N__19949\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26316\,
            in1 => \N__19713\,
            in2 => \N__19707\,
            in3 => \N__30431\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19973\,
            in1 => \N__19958\,
            in2 => \_gnd_net_\,
            in3 => \N__19948\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19929\,
            in1 => \N__19881\,
            in2 => \_gnd_net_\,
            in3 => \N__19904\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_8_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47369\,
            ce => \N__33626\,
            sr => \N__43835\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19839\,
            in1 => \N__19851\,
            in2 => \_gnd_net_\,
            in3 => \N__19817\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_15_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19818\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47369\,
            ce => \N__33626\,
            sr => \N__43835\
        );

    \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19857\,
            lcout => \pid_alt.error_d_reg_prev_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19794\,
            in1 => \N__20102\,
            in2 => \N__21047\,
            in3 => \N__30950\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19850\,
            in1 => \N__19838\,
            in2 => \_gnd_net_\,
            in3 => \N__19816\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20103\,
            in2 => \N__20106\,
            in3 => \N__30951\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__20072\,
            in1 => \_gnd_net_\,
            in2 => \N__20052\,
            in3 => \N__20094\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20093\,
            in1 => \N__20048\,
            in2 => \_gnd_net_\,
            in3 => \N__20071\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__20039\,
            in1 => \N__21086\,
            in2 => \N__20076\,
            in3 => \N__30185\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_14_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20073\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47356\,
            ce => \N__33629\,
            sr => \N__43841\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__20040\,
            in1 => \N__20025\,
            in2 => \_gnd_net_\,
            in3 => \N__30186\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_22_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__33630\,
            sr => \N__43849\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMMKM_0_23_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20186\,
            in1 => \N__20206\,
            in2 => \_gnd_net_\,
            in3 => \N__24612\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIMMKM_0Z0Z_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6BU12_22_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20226\,
            in2 => \N__20019\,
            in3 => \N__30703\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6BU12Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIKKKM_22_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__20016\,
            in1 => \N__20003\,
            in2 => \_gnd_net_\,
            in3 => \N__24613\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIKKKMZ0Z_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8IS34_22_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__20220\,
            in1 => \N__23052\,
            in2 => \N__20214\,
            in3 => \N__30704\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8IS34Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_23_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20207\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__33630\,
            sr => \N__43849\
        );

    \pid_alt.error_p_reg_esr_4_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20175\,
            lcout => \pid_alt.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47293\,
            ce => \N__46782\,
            sr => \N__46602\
        );

    \uart_drone_sync.Q_0__0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22329\,
            lcout => \debug_CH0_16A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20139\,
            in2 => \N__20160\,
            in3 => \N__20159\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_0\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20133\,
            in2 => \_gnd_net_\,
            in3 => \N__20127\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_0\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_1\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20124\,
            in2 => \_gnd_net_\,
            in3 => \N__20118\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_1\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_2\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20115\,
            in2 => \_gnd_net_\,
            in3 => \N__20109\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_2\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_3\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20402\,
            in2 => \_gnd_net_\,
            in3 => \N__20388\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_3\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_4\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20381\,
            in2 => \_gnd_net_\,
            in3 => \N__20367\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_4\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_5\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20360\,
            in2 => \_gnd_net_\,
            in3 => \N__20346\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_5\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_6\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20339\,
            in2 => \_gnd_net_\,
            in3 => \N__20325\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_6\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_7\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__22323\
        );

    \dron_frame_decoder_1.WDT_8_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20321\,
            in2 => \_gnd_net_\,
            in3 => \N__20307\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_8\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_9_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20300\,
            in2 => \_gnd_net_\,
            in3 => \N__20286\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_8\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_9\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_10_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20282\,
            in2 => \_gnd_net_\,
            in3 => \N__20268\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_9\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_10\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_11_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20263\,
            in2 => \_gnd_net_\,
            in3 => \N__20247\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_10\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_11\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_12_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20242\,
            in2 => \_gnd_net_\,
            in3 => \N__20538\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_11\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_12\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_13_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20523\,
            in2 => \_gnd_net_\,
            in3 => \N__20502\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_12\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_13\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_14_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20494\,
            in2 => \_gnd_net_\,
            in3 => \N__20475\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_13\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_14\,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.WDT_15_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20458\,
            in2 => \_gnd_net_\,
            in3 => \N__20472\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__22322\
        );

    \dron_frame_decoder_1.state_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__22515\,
            in1 => \N__20412\,
            in2 => \N__20559\,
            in3 => \N__20438\,
            lcout => \dron_frame_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => 'H',
            sr => \N__43800\
        );

    \dron_frame_decoder_1.state_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22516\,
            in1 => \N__22392\,
            in2 => \N__20427\,
            in3 => \N__29662\,
            lcout => \dron_frame_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => 'H',
            sr => \N__43800\
        );

    \dron_frame_decoder_1.state_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__29661\,
            in1 => \N__20423\,
            in2 => \N__20439\,
            in3 => \N__22514\,
            lcout => \dron_frame_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => 'H',
            sr => \N__43800\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26190\,
            in1 => \N__25209\,
            in2 => \N__25137\,
            in3 => \N__25002\,
            lcout => \dron_frame_decoder_1.N_188_4\,
            ltout => \dron_frame_decoder_1.N_188_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20677\,
            in1 => \_gnd_net_\,
            in2 => \N__20415\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23757\,
            in2 => \_gnd_net_\,
            in3 => \N__27039\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIC08S_3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20586\,
            in3 => \N__44088\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25090\,
            in2 => \_gnd_net_\,
            in3 => \N__25174\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24732\,
            in1 => \N__25042\,
            in2 => \N__20583\,
            in3 => \N__29657\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__22629\,
            in1 => \N__20580\,
            in2 => \N__20574\,
            in3 => \N__20565\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__22530\,
            in1 => \N__20658\,
            in2 => \N__20571\,
            in3 => \N__22648\,
            lcout => \dron_frame_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__43804\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25216\,
            in2 => \_gnd_net_\,
            in3 => \N__25009\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25138\,
            in1 => \N__22647\,
            in2 => \N__20568\,
            in3 => \N__26200\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_0_1\,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_1_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__20682\,
            in1 => \N__20555\,
            in2 => \N__20541\,
            in3 => \N__22529\,
            lcout => \dron_frame_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__43804\
        );

    \pid_alt.un9lto29_i_a2_7_c_RNO_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22739\,
            in2 => \_gnd_net_\,
            in3 => \N__22566\,
            lcout => \pid_alt.N_232_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIFPN33_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__20796\,
            in1 => \N__20787\,
            in2 => \N__30102\,
            in3 => \N__20738\,
            lcout => \pid_alt.error_p_reg_esr_RNIFPN33Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_12_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23708\,
            in2 => \_gnd_net_\,
            in3 => \N__27045\,
            lcout => \Commands_frame_decoder.N_354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIM4TM_16_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20910\,
            in1 => \N__20952\,
            in2 => \N__20868\,
            in3 => \N__20991\,
            lcout => \pid_alt.un9lto29_i_a2_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_1_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__22650\,
            in1 => \N__29713\,
            in2 => \N__20681\,
            in3 => \N__29667\,
            lcout => \dron_frame_decoder_1.state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20642\,
            in2 => \N__20649\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20622\,
            in2 => \N__30137\,
            in3 => \N__20610\,
            lcout => \pid_alt.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_0\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20607\,
            in2 => \N__30101\,
            in3 => \N__20601\,
            lcout => \pid_alt.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_0\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_1\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20598\,
            in2 => \N__30035\,
            in3 => \N__20589\,
            lcout => \pid_alt.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_1\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_2\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20853\,
            in2 => \N__29996\,
            in3 => \N__20844\,
            lcout => \pid_alt.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_2\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_3\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_4_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26114\,
            in2 => \N__26091\,
            in3 => \N__20841\,
            lcout => \pid_alt.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_3\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_4\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_5_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22668\,
            in2 => \N__26049\,
            in3 => \N__20838\,
            lcout => \pid_alt.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_4\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_5\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_6_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22698\,
            in2 => \N__22692\,
            in3 => \N__20835\,
            lcout => \pid_alt.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_5\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_6\,
            clk => \N__47397\,
            ce => \N__33600\,
            sr => \N__43810\
        );

    \pid_alt.pid_prereg_esr_7_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22752\,
            in2 => \N__22772\,
            in3 => \N__20832\,
            lcout => \pid_alt.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_7\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_8_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20829\,
            in2 => \N__26315\,
            in3 => \N__20817\,
            lcout => \pid_alt.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_7\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_8\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_9_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22779\,
            in2 => \N__22808\,
            in3 => \N__20814\,
            lcout => \pid_alt.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_8\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_9\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_10_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22980\,
            in2 => \N__22902\,
            in3 => \N__20811\,
            lcout => \pid_alt.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_9\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_10\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_11_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20808\,
            in2 => \N__23081\,
            in3 => \N__20799\,
            lcout => \pid_alt.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_10\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_11\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_12_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21165\,
            in2 => \N__21156\,
            in3 => \N__21144\,
            lcout => \pid_alt.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_11\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_12\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_13_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21141\,
            in2 => \N__21126\,
            in3 => \N__21105\,
            lcout => \pid_alt.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_12\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_13\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_14_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21102\,
            in2 => \N__21090\,
            in3 => \N__21066\,
            lcout => \pid_alt.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_13\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_14\,
            clk => \N__47383\,
            ce => \N__33603\,
            sr => \N__43816\
        );

    \pid_alt.pid_prereg_esr_15_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21063\,
            in2 => \N__21051\,
            in3 => \N__21027\,
            lcout => \pid_alt.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_15\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_16_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21024\,
            in2 => \N__21015\,
            in3 => \N__20982\,
            lcout => \pid_alt.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_15\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_16\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_17_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20979\,
            in2 => \N__20970\,
            in3 => \N__20943\,
            lcout => \pid_alt.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_16\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_17\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_18_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20940\,
            in2 => \N__20931\,
            in3 => \N__20901\,
            lcout => \pid_alt.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_17\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_18\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_19_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20898\,
            in2 => \N__20889\,
            in3 => \N__20856\,
            lcout => \pid_alt.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_18\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_19\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_20_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21237\,
            in2 => \N__21228\,
            in3 => \N__21207\,
            lcout => \pid_alt.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_19\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_20\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_21_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23256\,
            in2 => \N__23292\,
            in3 => \N__21204\,
            lcout => \pid_alt.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_20\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_21\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_22_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22998\,
            in2 => \N__23010\,
            in3 => \N__21201\,
            lcout => \pid_alt.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_21\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_22\,
            clk => \N__47370\,
            ce => \N__33607\,
            sr => \N__43820\
        );

    \pid_alt.pid_prereg_esr_23_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23045\,
            in2 => \N__21198\,
            in3 => \N__21183\,
            lcout => \pid_alt.pid_preregZ0Z_23\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_23\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_24_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26243\,
            in2 => \N__26220\,
            in3 => \N__21180\,
            lcout => \pid_alt.pid_preregZ0Z_24\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_23\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_24\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_25_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24239\,
            in2 => \N__24324\,
            in3 => \N__21177\,
            lcout => \pid_alt.pid_preregZ0Z_25\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_24\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_25\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_26_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24260\,
            in2 => \N__24384\,
            in3 => \N__21174\,
            lcout => \pid_alt.pid_preregZ0Z_26\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_25\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_26\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_27_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21279\,
            in2 => \N__24347\,
            in3 => \N__21171\,
            lcout => \pid_alt.pid_preregZ0Z_27\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_26\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_27\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_28_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21270\,
            in2 => \N__21246\,
            in3 => \N__21168\,
            lcout => \pid_alt.pid_preregZ0Z_28\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_27\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_28\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_29_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21990\,
            in2 => \N__22068\,
            in3 => \N__21285\,
            lcout => \pid_alt.pid_preregZ0Z_29\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_28\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_29\,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.pid_prereg_esr_30_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000101111110"
        )
    port map (
            in0 => \N__22015\,
            in1 => \N__30720\,
            in2 => \N__22053\,
            in3 => \N__21282\,
            lcout => \pid_alt.pid_preregZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47357\,
            ce => \N__33612\,
            sr => \N__43826\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8JT34_26_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22008\,
            in1 => \N__21260\,
            in2 => \N__24351\,
            in3 => \N__30718\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8JT34Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISSKM_26_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__23153\,
            in1 => \N__23138\,
            in2 => \_gnd_net_\,
            in3 => \N__24635\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNISSKMZ0Z_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMRU12_26_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__22009\,
            in1 => \_gnd_net_\,
            in2 => \N__21273\,
            in3 => \N__30717\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMRU12Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_26_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23139\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47345\,
            ce => \N__33616\,
            sr => \N__43836\
        );

    \pid_alt.error_d_reg_prev_esr_RNIUUKM_0_27_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24636\,
            in1 => \N__21494\,
            in2 => \_gnd_net_\,
            in3 => \N__21523\,
            lcout => \pid_alt.un1_pid_prereg_296_1\,
            ltout => \pid_alt.un1_pid_prereg_296_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIKQJO2_26_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__30719\,
            in1 => \N__21261\,
            in2 => \N__21249\,
            in3 => \N__22047\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIKQJO2Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_27_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21525\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47345\,
            ce => \N__33616\,
            sr => \N__43836\
        );

    \pid_alt.error_d_reg_prev_esr_RNIUUKM_27_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__21524\,
            in1 => \_gnd_net_\,
            in2 => \N__21498\,
            in3 => \N__24637\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIUUKMZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_1_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__45186\,
            in2 => \N__31849\,
            in3 => \N__21977\,
            lcout => alt_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__43842\
        );

    \Commands_frame_decoder.source_CH1data_2_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__36888\,
            in1 => \N__24100\,
            in2 => \N__21909\,
            in3 => \N__31842\,
            lcout => alt_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__43842\
        );

    \Commands_frame_decoder.source_CH1data_3_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__24101\,
            in1 => \N__43354\,
            in2 => \N__31850\,
            in3 => \N__21849\,
            lcout => alt_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__43842\
        );

    \pid_alt.error_cry_0_c_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23244\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \pid_alt.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_RNI1N2F_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23436\,
            in3 => \N__21438\,
            lcout => \pid_alt.error_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_0\,
            carryout => \pid_alt.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_1_c_RNI3Q3F_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23400\,
            in3 => \N__21393\,
            lcout => \pid_alt.error_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_1\,
            carryout => \pid_alt.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_2_c_RNI5T4F_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23229\,
            in3 => \N__21342\,
            lcout => \pid_alt.error_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_2\,
            carryout => \pid_alt.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_3_c_RNIKE1T_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23364\,
            in2 => \N__24810\,
            in3 => \N__21288\,
            lcout => \pid_alt.error_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_3\,
            carryout => \pid_alt.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_4_c_RNINI2T_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21978\,
            in2 => \N__24792\,
            in3 => \N__21912\,
            lcout => \pid_alt.error_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_4\,
            carryout => \pid_alt.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_5_c_RNIQM3T_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24774\,
            in2 => \N__21908\,
            in3 => \N__21852\,
            lcout => \pid_alt.error_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_5\,
            carryout => \pid_alt.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_6_c_RNITQ4T_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21848\,
            in2 => \N__24759\,
            in3 => \N__21783\,
            lcout => \pid_alt.error_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_6\,
            carryout => \pid_alt.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_7_c_RNI9LEM_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22098\,
            in2 => \N__24747\,
            in3 => \N__21729\,
            lcout => \pid_alt.error_8\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \pid_alt.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_8_c_RNICPFM_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22092\,
            in2 => \N__23373\,
            in3 => \N__21675\,
            lcout => \pid_alt.error_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_8\,
            carryout => \pid_alt.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_9_c_RNIMMUJ_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22083\,
            in2 => \N__23220\,
            in3 => \N__21630\,
            lcout => \pid_alt.error_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_9\,
            carryout => \pid_alt.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_10_c_RNI0SDO_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22074\,
            in2 => \N__23211\,
            in3 => \N__21582\,
            lcout => \pid_alt.error_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_10\,
            carryout => \pid_alt.error_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_11_c_RNI5JAH_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23427\,
            in3 => \N__21528\,
            lcout => \pid_alt.error_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_11\,
            carryout => \pid_alt.error_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_12_c_RNI7MBH_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23418\,
            in3 => \N__22209\,
            lcout => \pid_alt.error_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_12\,
            carryout => \pid_alt.error_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_13_c_RNI9PCH_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23409\,
            in3 => \N__22155\,
            lcout => \pid_alt.error_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_13\,
            carryout => \pid_alt.error_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_14_c_RNIBSDH_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25062\,
            in2 => \_gnd_net_\,
            in3 => \N__22152\,
            lcout => \pid_alt.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_esr_4_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45362\,
            lcout => alt_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47294\,
            ce => \N__31791\,
            sr => \N__43864\
        );

    \Commands_frame_decoder.source_CH1data_esr_5_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44290\,
            lcout => alt_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47294\,
            ce => \N__31791\,
            sr => \N__43864\
        );

    \Commands_frame_decoder.source_CH1data_esr_6_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33441\,
            lcout => alt_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47294\,
            ce => \N__31791\,
            sr => \N__43864\
        );

    \Commands_frame_decoder.source_CH1data_esr_7_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45014\,
            lcout => alt_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47294\,
            ce => \N__31791\,
            sr => \N__43864\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOTU12_27_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22052\,
            in1 => \N__22023\,
            in2 => \_gnd_net_\,
            in3 => \N__30706\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOTU12Z0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOTU12_0_27_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22051\,
            in1 => \N__22022\,
            in2 => \_gnd_net_\,
            in3 => \N__30651\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOTU12_0Z0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNICP2N1_0_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24135\,
            in2 => \_gnd_net_\,
            in3 => \N__46674\,
            lcout => \pid_alt.N_410_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_2__0__0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22281\,
            lcout => \uart_drone_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => \uart_drone_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_0__0__0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNID7P31_6_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23476\,
            in1 => \N__25406\,
            in2 => \_gnd_net_\,
            in3 => \N__25382\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__23456\,
            in1 => \N__22257\,
            in2 => \N__22260\,
            in3 => \N__22344\,
            lcout => \Commands_frame_decoder.WDT8lt14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__25427\,
            in1 => \N__25405\,
            in2 => \N__23607\,
            in3 => \N__25381\,
            lcout => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNII19A1_0_4_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23647\,
            in1 => \N__23494\,
            in2 => \N__23630\,
            in3 => \N__23512\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lto9_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNII01C2_6_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__23455\,
            in1 => \N__23477\,
            in2 => \N__22251\,
            in3 => \N__23605\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lt12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPJEG6_6_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22350\,
            in2 => \N__22353\,
            in3 => \N__25284\,
            lcout => \Commands_frame_decoder.state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIR9JL1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__25347\,
            in1 => \N__25308\,
            in2 => \N__25275\,
            in3 => \N__25426\,
            lcout => \Commands_frame_decoder.state_0_sqmuxacf1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNII19A1_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23648\,
            in1 => \N__23495\,
            in2 => \N__23631\,
            in3 => \N__23513\,
            lcout => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22338\,
            lcout => \uart_drone_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29668\,
            in2 => \_gnd_net_\,
            in3 => \N__44086\,
            lcout => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIJN1J_7_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23678\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIG48S_7_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22299\,
            in3 => \N__44087\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_2_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__25359\,
            in1 => \N__25316\,
            in2 => \N__27044\,
            in3 => \N__23663\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_322_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25238\,
            in2 => \N__22296\,
            in3 => \N__25616\,
            lcout => \Commands_frame_decoder.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIF38S_6_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__27009\,
            in1 => \N__25524\,
            in2 => \_gnd_net_\,
            in3 => \N__44068\,
            lcout => \Commands_frame_decoder.state_RNIF38SZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIQRI31_10_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__27010\,
            in1 => \_gnd_net_\,
            in2 => \N__23777\,
            in3 => \N__44067\,
            lcout => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_12_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__24863\,
            in1 => \N__26448\,
            in2 => \N__22431\,
            in3 => \N__26466\,
            lcout => \Commands_frame_decoder.stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47431\,
            ce => 'H',
            sr => \N__43801\
        );

    \Commands_frame_decoder.state_8_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__22413\,
            in1 => \N__22419\,
            in2 => \_gnd_net_\,
            in3 => \N__24862\,
            lcout => \Commands_frame_decoder.stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47431\,
            ce => 'H',
            sr => \N__43801\
        );

    \Commands_frame_decoder.state_RNIKO1J_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22412\,
            in2 => \_gnd_net_\,
            in3 => \N__27008\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0TLI1_5_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__22391\,
            in1 => \N__29705\,
            in2 => \N__22404\,
            in3 => \N__44082\,
            lcout => \dron_frame_decoder_1.N_392_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29642\,
            in2 => \_gnd_net_\,
            in3 => \N__22366\,
            lcout => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\,
            ltout => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__22389\,
            in2 => \N__22395\,
            in3 => \N__29704\,
            lcout => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__22367\,
            in1 => \N__22390\,
            in2 => \N__29663\,
            in3 => \N__22531\,
            lcout => \dron_frame_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47422\,
            ce => 'H',
            sr => \N__43805\
        );

    \dron_frame_decoder_1.state_7_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__22533\,
            in1 => \N__29643\,
            in2 => \N__22371\,
            in3 => \N__22494\,
            lcout => \dron_frame_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47422\,
            ce => 'H',
            sr => \N__43805\
        );

    \uart_drone.data_rdy_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31647\,
            lcout => uart_drone_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47422\,
            ce => 'H',
            sr => \N__43805\
        );

    \dron_frame_decoder_1.state_6_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__22532\,
            in1 => \N__22493\,
            in2 => \N__29714\,
            in3 => \N__29647\,
            lcout => \dron_frame_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47422\,
            ce => 'H',
            sr => \N__43805\
        );

    \pid_alt.un9lto29_i_a2_0_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22584\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \pid_alt.un9lto29_i_a2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_1_c_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24216\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2\,
            carryout => \pid_alt.un9lto29_i_a2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_2_c_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23904\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_0\,
            carryout => \pid_alt.un9lto29_i_a2_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_3_c_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22575\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_1\,
            carryout => \pid_alt.un9lto29_i_a2_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_4_c_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23891\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_2\,
            carryout => \pid_alt.un9lto29_i_a2_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_5_c_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23865\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_3\,
            carryout => \pid_alt.un9lto29_i_a2_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_6_c_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23994\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_4\,
            carryout => \pid_alt.un9lto29_i_a2_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_7_c_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22662\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pid_alt.un9lto29_i_a2_5\,
            carryout => \pid_alt.un9lto29_i_a2_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_7_c_RNIOG6V_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__33173\,
            in1 => \N__28043\,
            in2 => \_gnd_net_\,
            in3 => \N__22653\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24950\,
            in1 => \N__29601\,
            in2 => \_gnd_net_\,
            in3 => \N__33174\,
            lcout => \pid_alt.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__43811\
        );

    \dron_frame_decoder_1.state_RNO_2_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29712\,
            in2 => \_gnd_net_\,
            in3 => \N__22649\,
            lcout => \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI2K0N_20_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22623\,
            in1 => \N__22614\,
            in2 => \N__22605\,
            in3 => \N__22593\,
            lcout => \pid_alt.un9lto29_i_a2_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIDJJA1_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25951\,
            in1 => \N__23830\,
            in2 => \N__25886\,
            in3 => \N__25928\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_0_c_RNO_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25927\,
            in1 => \N__25975\,
            in2 => \N__25958\,
            in3 => \N__25879\,
            lcout => \pid_alt.source_pid10lt4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_3_c_RNO_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22716\,
            in1 => \N__23973\,
            in2 => \N__22548\,
            in3 => \N__23829\,
            lcout => \pid_alt.un9lto29_i_a2_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIK4VM_14_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22565\,
            in1 => \N__22544\,
            in2 => \N__22740\,
            in3 => \N__22715\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_12_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__23831\,
            in1 => \N__23972\,
            in2 => \N__28067\,
            in3 => \N__23813\,
            lcout => throttle_command_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47384\,
            ce => \N__27913\,
            sr => \N__27865\
        );

    \pid_alt.source_pid_1_esr_13_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__23814\,
            in1 => \N__28047\,
            in2 => \_gnd_net_\,
            in3 => \N__23974\,
            lcout => throttle_command_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47384\,
            ce => \N__27913\,
            sr => \N__27865\
        );

    \pid_alt.error_d_reg_prev_esr_5_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25809\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47371\,
            ce => \N__33601\,
            sr => \N__43821\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__25782\,
            in2 => \_gnd_net_\,
            in3 => \N__29880\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24539\,
            in1 => \N__24510\,
            in2 => \_gnd_net_\,
            in3 => \N__24487\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI171A6_5_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__22691\,
            in1 => \N__25781\,
            in2 => \N__22701\,
            in3 => \N__29879\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI171A6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICUVC3_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__24072\,
            in1 => \N__22677\,
            in2 => \_gnd_net_\,
            in3 => \N__29906\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICUVC3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__25848\,
            in1 => \N__25824\,
            in2 => \_gnd_net_\,
            in3 => \N__25808\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOGSO6_4_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24071\,
            in1 => \N__26048\,
            in2 => \N__22671\,
            in3 => \N__29905\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOGSO6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__22853\,
            in1 => \_gnd_net_\,
            in2 => \N__22866\,
            in3 => \N__22887\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__22901\,
            in1 => \N__23093\,
            in2 => \N__22983\,
            in3 => \N__30339\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__22970\,
            in1 => \N__22950\,
            in2 => \_gnd_net_\,
            in3 => \N__22932\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_9_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22854\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => \N__33604\,
            sr => \N__43827\
        );

    \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22824\,
            in1 => \N__22830\,
            in2 => \_gnd_net_\,
            in3 => \N__30378\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__22886\,
            in1 => \N__22862\,
            in2 => \_gnd_net_\,
            in3 => \N__22852\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22823\,
            in1 => \N__22809\,
            in2 => \N__22782\,
            in3 => \N__30377\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26345\,
            in1 => \N__26327\,
            in2 => \N__22773\,
            in3 => \N__30480\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__23202\,
            in1 => \N__23184\,
            in2 => \_gnd_net_\,
            in3 => \N__30770\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0AAT1_7_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23163\,
            in2 => \_gnd_net_\,
            in3 => \N__44083\,
            lcout => \dron_frame_decoder_1.N_384_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISSKM_0_26_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__23154\,
            in1 => \N__23132\,
            in2 => \_gnd_net_\,
            in3 => \N__24663\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISSKM_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__23100\,
            in1 => \N__23094\,
            in2 => \_gnd_net_\,
            in3 => \N__30338\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_21_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23322\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__33613\,
            sr => \N__43843\
        );

    \pid_alt.error_d_reg_prev_esr_RNI27U12_21_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__30697\,
            in1 => \N__23034\,
            in2 => \_gnd_net_\,
            in3 => \N__23028\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI27U12Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIIIKM_21_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__23321\,
            in1 => \_gnd_net_\,
            in2 => \N__23334\,
            in3 => \N__24658\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIIIKMZ0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0AS34_21_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__30696\,
            in1 => \N__23027\,
            in2 => \N__23013\,
            in3 => \N__22997\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0AS34Z0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIU2U12_20_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__23298\,
            in1 => \N__23277\,
            in2 => \_gnd_net_\,
            in3 => \N__30695\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIU2U12Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIIIKM_0_21_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24657\,
            in1 => \N__23330\,
            in2 => \_gnd_net_\,
            in3 => \N__23320\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIIIKM_0Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIQ8034_20_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__23291\,
            in1 => \N__23276\,
            in2 => \N__23259\,
            in3 => \N__30694\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIQ8034Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_inv_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23243\,
            in1 => \N__42886\,
            in2 => \_gnd_net_\,
            in3 => \N__24418\,
            lcout => \pid_alt.drone_altitude_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_3_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24390\,
            lcout => \pid_alt.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_6_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47314\,
            ce => \N__33617\,
            sr => \N__43850\
        );

    \pid_alt.error_i_acumm_prereg_esr_3_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29989\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47314\,
            ce => \N__33617\,
            sr => \N__43850\
        );

    \pid_alt.error_i_acumm_prereg_esr_13_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30219\,
            lcout => \pid_alt.error_i_acumm7lto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47314\,
            ce => \N__33617\,
            sr => \N__43850\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24705\,
            lcout => drone_altitude_i_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26157\,
            lcout => drone_altitude_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_1_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24402\,
            lcout => \pid_alt.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_12_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25182\,
            lcout => \pid_alt.error_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_13_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25146\,
            lcout => \pid_alt.error_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_14_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25098\,
            lcout => \pid_alt.error_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_2_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24396\,
            lcout => \pid_alt.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_0_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27662\,
            in2 => \_gnd_net_\,
            in3 => \N__46682\,
            lcout => alt_ki_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__44821\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24972\,
            lcout => drone_altitude_i_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_0_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__24102\,
            in1 => \N__27673\,
            in2 => \N__31851\,
            in3 => \N__23363\,
            lcout => alt_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__43873\
        );

    \pid_alt.error_p_reg_esr_5_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23349\,
            lcout => \pid_alt.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__46784\,
            sr => \N__46598\
        );

    \uart_pc_sync.aux_0__0__0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23571\,
            lcout => \uart_pc_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47475\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23547\,
            in2 => \N__23564\,
            in3 => \N__23565\,
            lcout => \Commands_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_0\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23541\,
            in2 => \_gnd_net_\,
            in3 => \N__23535\,
            lcout => \Commands_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_0\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_1\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23532\,
            in2 => \_gnd_net_\,
            in3 => \N__23526\,
            lcout => \Commands_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_1\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_2\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23523\,
            in2 => \_gnd_net_\,
            in3 => \N__23517\,
            lcout => \Commands_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_2\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_3\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23514\,
            in2 => \_gnd_net_\,
            in3 => \N__23499\,
            lcout => \Commands_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_3\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_4\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23496\,
            in2 => \_gnd_net_\,
            in3 => \N__23481\,
            lcout => \Commands_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_4\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_5\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23478\,
            in2 => \_gnd_net_\,
            in3 => \N__23460\,
            lcout => \Commands_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_5\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_6\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23457\,
            in2 => \_gnd_net_\,
            in3 => \N__23439\,
            lcout => \Commands_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_6\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_7\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__25439\
        );

    \Commands_frame_decoder.WDT_8_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23649\,
            in2 => \_gnd_net_\,
            in3 => \N__23634\,
            lcout => \Commands_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_8\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_9_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23629\,
            in2 => \_gnd_net_\,
            in3 => \N__23610\,
            lcout => \Commands_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_8\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_9\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_10_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23606\,
            in2 => \_gnd_net_\,
            in3 => \N__23589\,
            lcout => \Commands_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_9\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_10\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_11_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25383\,
            in2 => \_gnd_net_\,
            in3 => \N__23586\,
            lcout => \Commands_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_10\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_11\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_12_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25407\,
            in2 => \_gnd_net_\,
            in3 => \N__23583\,
            lcout => \Commands_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_11\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_12\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_13_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25428\,
            in2 => \_gnd_net_\,
            in3 => \N__23580\,
            lcout => \Commands_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_12\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_13\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_14_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25315\,
            in2 => \_gnd_net_\,
            in3 => \N__23577\,
            lcout => \Commands_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_13\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_14\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.WDT_15_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25354\,
            in2 => \_gnd_net_\,
            in3 => \N__23574\,
            lcout => \Commands_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__25440\
        );

    \Commands_frame_decoder.state_RNI4OPK_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26476\,
            in2 => \_gnd_net_\,
            in3 => \N__25581\,
            lcout => \Commands_frame_decoder.N_320_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27041\,
            in1 => \N__43286\,
            in2 => \N__33404\,
            in3 => \N__25599\,
            lcout => \Commands_frame_decoder.N_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__25617\,
            in1 => \N__24861\,
            in2 => \N__25539\,
            in3 => \N__23727\,
            lcout => \Commands_frame_decoder.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47432\,
            ce => 'H',
            sr => \N__43802\
        );

    \Commands_frame_decoder.state_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__25562\,
            in1 => \N__25584\,
            in2 => \N__25227\,
            in3 => \N__24859\,
            lcout => \Commands_frame_decoder.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47432\,
            ce => 'H',
            sr => \N__43802\
        );

    \Commands_frame_decoder.state_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25563\,
            in1 => \N__25590\,
            in2 => \N__23721\,
            in3 => \N__24860\,
            lcout => \Commands_frame_decoder.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47432\,
            ce => 'H',
            sr => \N__43802\
        );

    \Commands_frame_decoder.state_RNIEI1J_2_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23717\,
            in2 => \_gnd_net_\,
            in3 => \N__26972\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_11_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__23701\,
            in1 => \N__26989\,
            in2 => \N__23778\,
            in3 => \N__24853\,
            lcout => \Commands_frame_decoder.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.state_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__24858\,
            in1 => \N__25528\,
            in2 => \N__23682\,
            in3 => \N__26998\,
            lcout => \Commands_frame_decoder.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.state_6_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__25529\,
            in1 => \N__25716\,
            in2 => \_gnd_net_\,
            in3 => \N__24857\,
            lcout => \Commands_frame_decoder.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__25358\,
            in1 => \N__25317\,
            in2 => \N__27026\,
            in3 => \N__23667\,
            lcout => \Commands_frame_decoder.N_358\,
            ltout => \Commands_frame_decoder.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_10_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__23776\,
            in1 => \_gnd_net_\,
            in2 => \N__23781\,
            in3 => \N__27348\,
            lcout => \Commands_frame_decoder.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.state_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__24854\,
            in1 => \N__23753\,
            in2 => \_gnd_net_\,
            in3 => \N__31810\,
            lcout => \Commands_frame_decoder.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.state_4_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__23739\,
            in1 => \N__25479\,
            in2 => \_gnd_net_\,
            in3 => \N__24855\,
            lcout => \Commands_frame_decoder.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \Commands_frame_decoder.state_5_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__24856\,
            in1 => \N__25467\,
            in2 => \_gnd_net_\,
            in3 => \N__25728\,
            lcout => \Commands_frame_decoder.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__43806\
        );

    \uart_drone.data_esr_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25703\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25688\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25673\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_3_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25644\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_5_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_6_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25769\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \uart_drone.data_esr_7_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25754\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__26601\,
            sr => \N__26619\
        );

    \Commands_frame_decoder.source_offset3data_ess_7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44984\,
            lcout => \frame_decoder_OFF3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47399\,
            ce => \N__26744\,
            sr => \N__43812\
        );

    \pid_alt.pid_prereg_esr_RNIU1UR2_14_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23990\,
            in1 => \N__23892\,
            in2 => \N__23877\,
            in3 => \N__23864\,
            lcout => \pid_alt.N_123\,
            ltout => \pid_alt.N_123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI0T1S7_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23850\,
            in1 => \N__24144\,
            in2 => \N__23841\,
            in3 => \N__23942\,
            lcout => \pid_alt.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIH58S_8_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24881\,
            in2 => \_gnd_net_\,
            in3 => \N__44085\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIV9C73_12_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__23979\,
            in1 => \N__23838\,
            in2 => \_gnd_net_\,
            in3 => \N__23812\,
            lcout => \pid_alt.N_106\,
            ltout => \pid_alt.N_106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIIJ486_30_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000011"
        )
    port map (
            in0 => \N__23943\,
            in1 => \N__28068\,
            in2 => \N__23799\,
            in3 => \N__24207\,
            lcout => \pid_alt.N_91_1\,
            ltout => \pid_alt.N_91_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_7_c_RNI7EJCF_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__23796\,
            in1 => \N__23790\,
            in2 => \N__23784\,
            in3 => \N__32928\,
            lcout => \pid_alt.un1_reset_0_i\,
            ltout => \pid_alt.un1_reset_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIS3RQF_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24048\,
            in3 => \N__33181\,
            lcout => \pid_alt.N_96_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNII41N_24_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24045\,
            in1 => \N__24033\,
            in2 => \N__24021\,
            in3 => \N__24006\,
            lcout => \pid_alt.un9lto29_i_a2_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_5_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__27977\,
            in1 => \N__23941\,
            in2 => \N__24198\,
            in3 => \N__28065\,
            lcout => throttle_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__27912\,
            sr => \N__27863\
        );

    \pid_alt.source_pid_1_esr_10_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__27105\,
            in1 => \_gnd_net_\,
            in2 => \N__28072\,
            in3 => \N__27975\,
            lcout => throttle_command_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__27912\,
            sr => \N__27863\
        );

    \pid_alt.source_pid_1_esr_11_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__27976\,
            in1 => \N__28057\,
            in2 => \_gnd_net_\,
            in3 => \N__27140\,
            lcout => throttle_command_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__27912\,
            sr => \N__27863\
        );

    \pid_alt.source_pid_1_esr_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__27978\,
            in1 => \_gnd_net_\,
            in2 => \N__27177\,
            in3 => \N__28058\,
            lcout => throttle_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__27912\,
            sr => \N__27863\
        );

    \pid_alt.source_pid_1_esr_8_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__23925\,
            in1 => \_gnd_net_\,
            in2 => \N__28073\,
            in3 => \N__27979\,
            lcout => throttle_command_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__27912\,
            sr => \N__27863\
        );

    \pid_alt.pid_prereg_esr_RNI0VB22_6_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26006\,
            in1 => \N__23975\,
            in2 => \N__27078\,
            in3 => \N__23921\,
            lcout => \pid_alt.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_2_c_RNO_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__27097\,
            in2 => \N__27136\,
            in3 => \N__23920\,
            lcout => \pid_alt.N_12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9lto29_i_a2_1_c_RNO_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24195\,
            in1 => \N__26005\,
            in2 => \N__27170\,
            in3 => \N__24166\,
            lcout => \pid_alt.un9lto29_i_a2_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI35JO_4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__24168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24197\,
            lcout => \pid_alt.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIL84J1_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24196\,
            in1 => \N__24167\,
            in2 => \N__33172\,
            in3 => \N__25986\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24957\,
            lcout => \pid_alt.N_96_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => 'H',
            sr => \N__43828\
        );

    \pid_alt.state_RNIFCSD1_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__33146\,
            in1 => \N__29590\,
            in2 => \N__24962\,
            in3 => \N__44066\,
            lcout => \pid_alt.state_RNIFCSD1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto7_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26361\,
            in1 => \N__25862\,
            in2 => \N__45351\,
            in3 => \N__33405\,
            lcout => \Commands_frame_decoder.source_CH1data8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__45494\,
            in1 => \_gnd_net_\,
            in2 => \N__26022\,
            in3 => \N__24063\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24062\,
            in1 => \N__26018\,
            in2 => \_gnd_net_\,
            in3 => \N__45493\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIQQKM_25_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24300\,
            in1 => \N__24312\,
            in2 => \_gnd_net_\,
            in3 => \N__24662\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIQQKMZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0BT34_25_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30699\,
            in1 => \N__24359\,
            in2 => \N__24261\,
            in3 => \N__24368\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0BT34Z0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIINU12_25_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__30702\,
            in1 => \N__24369\,
            in2 => \_gnd_net_\,
            in3 => \N__24360\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIINU12Z0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_25_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24299\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47331\,
            ce => \N__33605\,
            sr => \N__43844\
        );

    \pid_alt.error_d_reg_prev_esr_RNIO2T34_24_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24548\,
            in1 => \N__24270\,
            in2 => \N__24240\,
            in3 => \N__30701\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIO2T34Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIQQKM_0_25_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24311\,
            in1 => \N__24298\,
            in2 => \_gnd_net_\,
            in3 => \N__24661\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIQQKM_0Z0Z_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIEJU12_24_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__24549\,
            in1 => \_gnd_net_\,
            in2 => \N__24264\,
            in3 => \N__30700\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIEJU12Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_24_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47315\,
            ce => \N__33608\,
            sr => \N__43851\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOOKM_0_24_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24698\,
            in1 => \N__24688\,
            in2 => \_gnd_net_\,
            in3 => \N__24659\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIOOKM_0Z0Z_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIAFU12_23_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26280\,
            in2 => \N__24243\,
            in3 => \N__30698\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIAFU12Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOOKM_24_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__24699\,
            in1 => \N__24689\,
            in2 => \_gnd_net_\,
            in3 => \N__24660\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOOKMZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24540\,
            in1 => \N__24509\,
            in2 => \_gnd_net_\,
            in3 => \N__24494\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_0_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25049\,
            lcout => drone_altitude_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25010\,
            lcout => drone_altitude_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_2_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_3_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_4_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25217\,
            lcout => \dron_frame_decoder_1.drone_altitude_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_5_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.drone_altitude_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_6_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25139\,
            lcout => \dron_frame_decoder_1.drone_altitude_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \dron_frame_decoder_1.source_Altitude_esr_7_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25091\,
            lcout => \dron_frame_decoder_1.drone_altitude_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__24900\,
            sr => \N__43857\
        );

    \Commands_frame_decoder.state_9_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__27059\,
            in1 => \N__24888\,
            in2 => \_gnd_net_\,
            in3 => \N__24867\,
            lcout => \Commands_frame_decoder.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47296\,
            ce => 'H',
            sr => \N__43865\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24816\,
            lcout => drone_altitude_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24798\,
            lcout => drone_altitude_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24780\,
            lcout => drone_altitude_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24765\,
            lcout => drone_altitude_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25020\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_10_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.drone_altitude_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_12_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25218\,
            lcout => drone_altitude_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_13_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_14_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25140\,
            lcout => drone_altitude_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_15_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25092\,
            lcout => drone_altitude_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_8_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25053\,
            lcout => \dron_frame_decoder_1.drone_altitude_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \dron_frame_decoder_1.source_Altitude_esr_9_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25011\,
            lcout => \dron_frame_decoder_1.drone_altitude_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__26148\,
            sr => \N__43874\
        );

    \Commands_frame_decoder.source_CH4data_esr_4_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45358\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => \N__26396\,
            sr => \N__43879\
        );

    \pid_alt.state_RNIH1EN_0_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24966\,
            in2 => \_gnd_net_\,
            in3 => \N__44069\,
            lcout => \pid_alt.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25461\,
            lcout => \uart_pc_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25446\,
            lcout => \uart_pc_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_1__0__0_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25455\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.un1_state53_i_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27027\,
            in2 => \_gnd_net_\,
            in3 => \N__44099\,
            lcout => \Commands_frame_decoder.un1_state53_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIRGQ51_11_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__25425\,
            in1 => \N__25404\,
            in2 => \_gnd_net_\,
            in3 => \N__25380\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_0_sqmuxacf0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIC9QE2_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__25266\,
            in1 => \N__25346\,
            in2 => \N__25320\,
            in3 => \N__25307\,
            lcout => \Commands_frame_decoder.state_0_sqmuxacf0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27028\,
            in2 => \_gnd_net_\,
            in3 => \N__25267\,
            lcout => \Commands_frame_decoder.preinitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__43799\
        );

    \Commands_frame_decoder.source_data_valid_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__25268\,
            in1 => \N__25251\,
            in2 => \N__27043\,
            in3 => \N__30528\,
            lcout => \debug_CH3_20A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__43799\
        );

    \Commands_frame_decoder.source_data_valid_RNO_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__26654\,
            in1 => \N__26634\,
            in2 => \_gnd_net_\,
            in3 => \N__26482\,
            lcout => \Commands_frame_decoder.count_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26499\,
            in1 => \N__25242\,
            in2 => \N__44271\,
            in3 => \N__36839\,
            lcout => \Commands_frame_decoder.state_ns_0_a4_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_3_0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25615\,
            in1 => \N__44254\,
            in2 => \N__36866\,
            in3 => \N__26498\,
            lcout => \Commands_frame_decoder.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45274\,
            in2 => \_gnd_net_\,
            in3 => \N__45176\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_2_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44954\,
            in2 => \_gnd_net_\,
            in3 => \N__27615\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a4_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_2_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__44258\,
            in1 => \N__36838\,
            in2 => \N__25593\,
            in3 => \N__25583\,
            lcout => \Commands_frame_decoder.state_ns_0_a4_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_4_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__27616\,
            in1 => \N__25866\,
            in2 => \N__36867\,
            in3 => \N__25582\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010101"
        )
    port map (
            in0 => \N__26444\,
            in1 => \N__25561\,
            in2 => \N__25548\,
            in3 => \N__25545\,
            lcout => \Commands_frame_decoder.state_ns_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_4_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__25493\,
            in1 => \N__27022\,
            in2 => \N__25530\,
            in3 => \N__45296\,
            lcout => alt_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47401\,
            ce => 'H',
            sr => \N__43807\
        );

    \uart_pc.data_rdy_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31228\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47401\,
            ce => 'H',
            sr => \N__43807\
        );

    \Commands_frame_decoder.state_RNIGK1J_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25478\,
            in2 => \_gnd_net_\,
            in3 => \N__27020\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNID18S_4_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25731\,
            in3 => \N__44073\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIHL1J_5_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25727\,
            in2 => \_gnd_net_\,
            in3 => \N__27021\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIE28S_5_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25707\,
            in3 => \N__44072\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__26556\,
            in1 => \N__31382\,
            in2 => \N__25704\,
            in3 => \N__31430\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31431\,
            in1 => \N__26550\,
            in2 => \N__25689\,
            in3 => \N__31389\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__34089\,
            in1 => \N__31383\,
            in2 => \N__25674\,
            in3 => \N__31432\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31433\,
            in1 => \N__27507\,
            in2 => \N__25659\,
            in3 => \N__31390\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_4_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__27519\,
            in1 => \N__25643\,
            in2 => \N__31397\,
            in3 => \N__31434\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_5_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31435\,
            in1 => \N__27693\,
            in2 => \N__25632\,
            in3 => \N__31391\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__34077\,
            in1 => \N__31384\,
            in2 => \N__25770\,
            in3 => \N__31436\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \uart_drone.data_Aux_7_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__31437\,
            in1 => \N__31388\,
            in2 => \N__25755\,
            in3 => \N__44468\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => 'H',
            sr => \N__31869\
        );

    \Commands_frame_decoder.source_CH3data_esr_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27652\,
            lcout => \frame_decoder_CH3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45211\,
            lcout => \frame_decoder_CH3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_2_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_3_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43339\,
            lcout => \frame_decoder_CH3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45314\,
            lcout => \frame_decoder_CH3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44262\,
            lcout => \frame_decoder_CH3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_esr_6_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33389\,
            lcout => \frame_decoder_CH3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \Commands_frame_decoder.source_CH3data_ess_7_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44983\,
            lcout => \frame_decoder_CH3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__25740\,
            sr => \N__43813\
        );

    \pid_alt.source_pid_1_esr_6_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__28074\,
            in1 => \N__27980\,
            in2 => \_gnd_net_\,
            in3 => \N__26010\,
            lcout => throttle_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => \N__27917\,
            sr => \N__27862\
        );

    \pid_alt.source_pid_1_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33163\,
            in1 => \N__25904\,
            in2 => \N__36992\,
            in3 => \N__25985\,
            lcout => throttle_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__27864\
        );

    \pid_alt.source_pid_1_1_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__25905\,
            in1 => \N__33164\,
            in2 => \N__29300\,
            in3 => \N__25959\,
            lcout => throttle_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__27864\
        );

    \pid_alt.source_pid_1_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33165\,
            in1 => \N__25906\,
            in2 => \N__29345\,
            in3 => \N__25932\,
            lcout => throttle_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__27864\
        );

    \pid_alt.source_pid_1_3_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__25907\,
            in1 => \N__33166\,
            in2 => \N__35477\,
            in3 => \N__25887\,
            lcout => throttle_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__27864\
        );

    \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__29014\,
            in1 => \N__28981\,
            in2 => \_gnd_net_\,
            in3 => \N__28945\,
            lcout => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_1_1_0_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44263\,
            in2 => \_gnd_net_\,
            in3 => \N__45001\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_1_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__25847\,
            in1 => \N__25823\,
            in2 => \_gnd_net_\,
            in3 => \N__25802\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIRFO19_3_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26075\,
            in1 => \N__29947\,
            in2 => \N__26118\,
            in3 => \N__26058\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIRFO19Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26076\,
            in1 => \N__26057\,
            in2 => \_gnd_net_\,
            in3 => \N__29948\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_4_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45495\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47317\,
            ce => \N__33598\,
            sr => \N__43837\
        );

    \pid_alt.error_i_acumm_prereg_esr_4_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm7lto4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47317\,
            ce => \N__33598\,
            sr => \N__43837\
        );

    \pid_alt.error_i_acumm_prereg_esr_5_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29910\,
            lcout => \pid_alt.error_i_acumm7lto5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47317\,
            ce => \N__33598\,
            sr => \N__43837\
        );

    \Commands_frame_decoder.source_CH4data_esr_1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45214\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \Commands_frame_decoder.source_CH4data_esr_2_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36865\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \Commands_frame_decoder.source_CH4data_esr_3_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43349\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \Commands_frame_decoder.source_CH4data_esr_0_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27669\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \Commands_frame_decoder.source_CH4data_esr_6_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33409\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \Commands_frame_decoder.source_CH4data_ess_7_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45005\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => \N__26383\,
            sr => \N__43845\
        );

    \CONSTANT_ONE_LUT4_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__43342\,
            in1 => \N__36857\,
            in2 => \_gnd_net_\,
            in3 => \N__45204\,
            lcout => \Commands_frame_decoder.source_CH1data8lt7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__26352\,
            in1 => \N__26328\,
            in2 => \_gnd_net_\,
            in3 => \N__30479\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGQS34_23_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26286\,
            in1 => \N__26279\,
            in2 => \N__26250\,
            in3 => \N__30705\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGQS34Z0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_11_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26205\,
            lcout => \dron_frame_decoder_1.drone_altitude_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47283\,
            ce => \N__26147\,
            sr => \N__43866\
        );

    \pid_alt.error_i_acumm_prereg_esr_7_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47270\,
            ce => \N__33618\,
            sr => \N__43880\
        );

    \pid_alt.error_i_acumm_prereg_esr_15_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30944\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47270\,
            ce => \N__33618\,
            sr => \N__43880\
        );

    \pid_alt.error_i_acumm_prereg_esr_6_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29870\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47270\,
            ce => \N__33618\,
            sr => \N__43880\
        );

    \uart_pc_sync.Q_0__0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26421\,
            lcout => \debug_CH2_18A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__26535\,
            in1 => \N__26510\,
            in2 => \N__26538\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27495\,
            in3 => \N__26415\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31615\,
            in3 => \N__26412\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31489\,
            in2 => \_gnd_net_\,
            in3 => \N__26409\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__44104\,
            in1 => \N__27462\,
            in2 => \N__27555\,
            in3 => \N__26406\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__26537\,
            in1 => \N__27547\,
            in2 => \N__27467\,
            in3 => \N__44105\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__31601\,
            in1 => \N__27490\,
            in2 => \N__31505\,
            in3 => \N__31546\,
            lcout => \uart_pc.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__31547\,
            in1 => \N__31271\,
            in2 => \N__44135\,
            in3 => \N__31490\,
            lcout => \uart_pc.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIMQ8T1_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26574\,
            in2 => \_gnd_net_\,
            in3 => \N__44079\,
            lcout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__27553\,
            in1 => \N__26544\,
            in2 => \N__27468\,
            in3 => \N__44081\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26536\,
            in2 => \_gnd_net_\,
            in3 => \N__26511\,
            lcout => OPEN,
            ltout => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__44080\,
            in1 => \N__27463\,
            in2 => \N__26514\,
            in3 => \N__27552\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_0_a4_0_0_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44914\,
            in2 => \_gnd_net_\,
            in3 => \N__27613\,
            lcout => \Commands_frame_decoder.state_ns_0_a4_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIVGCQ_12_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26484\,
            lcout => \Commands_frame_decoder.state_ns_i_a4_2_0_0\,
            ltout => \Commands_frame_decoder.state_ns_i_a4_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26650\,
            in2 => \N__26487\,
            in3 => \N__44107\,
            lcout => \Commands_frame_decoder.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNI0V5H1_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__26649\,
            in1 => \N__26632\,
            in2 => \N__26999\,
            in3 => \N__26483\,
            lcout => \Commands_frame_decoder.N_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__33840\,
            in1 => \N__37320\,
            in2 => \_gnd_net_\,
            in3 => \N__33791\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__44106\,
            in1 => \N__26430\,
            in2 => \N__26655\,
            in3 => \N__26633\,
            lcout => \Commands_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__31060\,
            in1 => \N__30992\,
            in2 => \N__28878\,
            in3 => \N__27614\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26708\,
            in2 => \_gnd_net_\,
            in3 => \N__26685\,
            lcout => \scaler_3.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__37319\,
            in1 => \N__33786\,
            in2 => \N__33849\,
            in3 => \N__34818\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_4_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__26586\,
            in1 => \N__31043\,
            in2 => \N__28824\,
            in3 => \N__45297\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__31370\,
            in1 => \N__31642\,
            in2 => \_gnd_net_\,
            in3 => \N__44075\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__31643\,
            in1 => \_gnd_net_\,
            in2 => \N__26604\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.data_rdyc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__31178\,
            in1 => \N__26584\,
            in2 => \_gnd_net_\,
            in3 => \N__44078\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__44423\,
            in1 => \N__36691\,
            in2 => \_gnd_net_\,
            in3 => \N__39516\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__39517\,
            in1 => \N__36692\,
            in2 => \_gnd_net_\,
            in3 => \N__44424\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.N_1239_i_l_ofx_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26709\,
            in2 => \_gnd_net_\,
            in3 => \N__26684\,
            lcout => \scaler_3.N_1239_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28103\,
            in2 => \_gnd_net_\,
            in3 => \N__28091\,
            lcout => \scaler_2.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27651\,
            lcout => \frame_decoder_CH2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45190\,
            lcout => \frame_decoder_CH2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36856\,
            lcout => \frame_decoder_CH2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45313\,
            lcout => \frame_decoder_CH2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44249\,
            lcout => \frame_decoder_CH2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_esr_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33393\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_CH2data_ess_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47362\,
            ce => \N__26670\,
            sr => \N__43817\
        );

    \Commands_frame_decoder.source_offset3data_esr_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27654\,
            lcout => \frame_decoder_OFF3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45212\,
            lcout => \frame_decoder_OFF3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36872\,
            lcout => \frame_decoder_OFF3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43340\,
            lcout => \frame_decoder_OFF3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45330\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44250\,
            lcout => \frame_decoder_OFF3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \Commands_frame_decoder.source_offset3data_esr_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33394\,
            lcout => \frame_decoder_OFF3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__26751\,
            sr => \N__43822\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28944\,
            in2 => \N__28980\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26733\,
            in2 => \N__26727\,
            in3 => \N__26712\,
            lcout => \scaler_3.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_0\,
            carryout => \scaler_3.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26895\,
            in2 => \N__26886\,
            in3 => \N__26877\,
            lcout => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_1\,
            carryout => \scaler_3.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26874\,
            in2 => \N__26865\,
            in3 => \N__26856\,
            lcout => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_2\,
            carryout => \scaler_3.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26853\,
            in2 => \N__26841\,
            in3 => \N__26832\,
            lcout => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_3\,
            carryout => \scaler_3.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26829\,
            in2 => \N__26817\,
            in3 => \N__26805\,
            lcout => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_4\,
            carryout => \scaler_3.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26802\,
            in2 => \N__26790\,
            in3 => \N__26781\,
            lcout => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_5\,
            carryout => \scaler_3.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26778\,
            in2 => \_gnd_net_\,
            in3 => \N__26769\,
            lcout => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_6\,
            carryout => \scaler_3.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26766\,
            in2 => \N__42916\,
            in3 => \N__26757\,
            lcout => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26754\,
            lcout => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI7G141_10_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27166\,
            in1 => \N__27947\,
            in2 => \N__27141\,
            in3 => \N__27104\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNILP1J_9_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27066\,
            in2 => \_gnd_net_\,
            in3 => \N__27042\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27655\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45213\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36873\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43341\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45331\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_5_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44270\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_esr_6_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33413\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \Commands_frame_decoder.source_offset4data_ess_7_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44988\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => \N__27327\,
            sr => \N__43846\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29493\,
            in2 => \N__29550\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27309\,
            in2 => \N__27303\,
            in3 => \N__27294\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27291\,
            in2 => \N__27285\,
            in3 => \N__27273\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27270\,
            in2 => \N__27264\,
            in3 => \N__27255\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27252\,
            in2 => \N__27237\,
            in3 => \N__27228\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27225\,
            in2 => \N__27219\,
            in3 => \N__27201\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27198\,
            in2 => \N__27192\,
            in3 => \N__27183\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27384\,
            in2 => \_gnd_net_\,
            in3 => \N__27180\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27354\,
            in2 => \N__42841\,
            in3 => \N__27390\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27387\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27365\,
            in2 => \_gnd_net_\,
            in3 => \N__27377\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_1251_i_l_ofx_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27378\,
            in1 => \_gnd_net_\,
            in2 => \N__27369\,
            in3 => \_gnd_net_\,
            lcout => \scaler_4.N_1251_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNII68S_9_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27341\,
            in2 => \_gnd_net_\,
            in3 => \N__44091\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_1_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30085\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47275\,
            ce => \N__33606\,
            sr => \N__43875\
        );

    \pid_alt.error_i_acumm_prereg_esr_16_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30913\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47275\,
            ce => \N__33606\,
            sr => \N__43875\
        );

    \pid_alt.error_i_acumm_prereg_esr_11_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30298\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47275\,
            ce => \N__33606\,
            sr => \N__43875\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27423\,
            in1 => \N__27402\,
            in2 => \N__27417\,
            in3 => \N__27315\,
            lcout => OPEN,
            ltout => \pid_alt.m7_e_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27396\,
            in1 => \N__27435\,
            in2 => \N__27429\,
            in3 => \N__27408\,
            lcout => \pid_alt.N_238\,
            ltout => \pid_alt.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111010"
        )
    port map (
            in0 => \N__32845\,
            in1 => \N__28595\,
            in2 => \N__27426\,
            in3 => \N__32822\,
            lcout => \pid_alt.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_18_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30839\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47271\,
            ce => \N__33609\,
            sr => \N__43881\
        );

    \pid_alt.error_i_acumm_prereg_esr_19_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30800\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47271\,
            ce => \N__33609\,
            sr => \N__43881\
        );

    \pid_alt.error_i_acumm_prereg_esr_14_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30179\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47271\,
            ce => \N__33609\,
            sr => \N__43881\
        );

    \pid_alt.error_i_acumm_prereg_esr_2_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30028\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_17_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30875\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_20_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30766\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_12_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30254\,
            lcout => \pid_alt.error_i_acumm7lto12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_10_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30334\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_21_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__33614\,
            sr => \N__43885\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_0_6_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28732\,
            in1 => \N__28552\,
            in2 => \N__28718\,
            in3 => \N__33274\,
            lcout => \pid_alt.m21_e_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIE3BQ1_6_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28733\,
            in1 => \N__28553\,
            in2 => \N__28719\,
            in3 => \N__33275\,
            lcout => \pid_alt.m35_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_8_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47265\,
            ce => \N__33619\,
            sr => \N__43889\
        );

    \pid_alt.error_i_acumm_prereg_esr_9_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30376\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47265\,
            ce => \N__33619\,
            sr => \N__43889\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31605\,
            in2 => \_gnd_net_\,
            in3 => \N__27494\,
            lcout => \uart_pc.N_126_li\,
            ltout => \uart_pc.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__27477\,
            in1 => \N__31554\,
            in2 => \N__27471\,
            in3 => \N__31709\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__31710\,
            in1 => \N__31503\,
            in2 => \N__31113\,
            in3 => \N__31606\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => \uart_pc.timer_Count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__27444\,
            in1 => \N__27554\,
            in2 => \N__27438\,
            in3 => \N__44125\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__44102\,
            in1 => \N__31722\,
            in2 => \N__28539\,
            in3 => \N__27551\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__31504\,
            in1 => \N__31611\,
            in2 => \N__31112\,
            in3 => \N__31721\,
            lcout => OPEN,
            ltout => \uart_pc.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__31108\,
            in1 => \N__28535\,
            in2 => \N__27522\,
            in3 => \N__44103\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_5_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__33345\,
            in1 => \N__31068\,
            in2 => \N__31001\,
            in3 => \N__28781\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIEAGS_4_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__31711\,
            in1 => \N__31555\,
            in2 => \_gnd_net_\,
            in3 => \N__44089\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_6_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__30990\,
            in1 => \N__29123\,
            in2 => \N__31074\,
            in3 => \N__44946\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__36819\,
            in1 => \N__31067\,
            in2 => \N__28842\,
            in3 => \N__30991\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__39518\,
            in1 => \N__36679\,
            in2 => \_gnd_net_\,
            in3 => \N__44420\,
            lcout => \uart_drone.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__44421\,
            in1 => \N__36687\,
            in2 => \_gnd_net_\,
            in3 => \N__39502\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__39503\,
            in1 => \_gnd_net_\,
            in2 => \N__36693\,
            in3 => \N__44422\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_4_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__31052\,
            in1 => \N__31000\,
            in2 => \N__28800\,
            in3 => \N__44205\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset2data_esr_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27653\,
            lcout => \frame_decoder_OFF2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45161\,
            lcout => \frame_decoder_OFF2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36855\,
            lcout => \frame_decoder_OFF2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43308\,
            lcout => \frame_decoder_OFF2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45298\,
            lcout => \frame_decoder_OFF2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44206\,
            lcout => \frame_decoder_OFF2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_esr_6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33362\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \Commands_frame_decoder.source_offset2data_ess_7_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44953\,
            lcout => \frame_decoder_OFF2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__27567\,
            sr => \N__43818\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29035\,
            in2 => \N__29081\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27810\,
            in2 => \N__27804\,
            in3 => \N__27795\,
            lcout => \scaler_2.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_0\,
            carryout => \scaler_2.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27792\,
            in2 => \N__27786\,
            in3 => \N__27777\,
            lcout => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_1\,
            carryout => \scaler_2.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27774\,
            in2 => \N__27768\,
            in3 => \N__27759\,
            lcout => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_2\,
            carryout => \scaler_2.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27756\,
            in2 => \N__27750\,
            in3 => \N__27741\,
            lcout => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_3\,
            carryout => \scaler_2.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27738\,
            in2 => \N__27732\,
            in3 => \N__27723\,
            lcout => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_4\,
            carryout => \scaler_2.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27720\,
            in2 => \N__27714\,
            in3 => \N__27705\,
            lcout => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_5\,
            carryout => \scaler_2.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__27696\,
            lcout => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_6\,
            carryout => \scaler_2.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28080\,
            in2 => \N__43123\,
            in3 => \N__28113\,
            lcout => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28110\,
            lcout => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42274\,
            in2 => \_gnd_net_\,
            in3 => \N__42010\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.N_1227_i_l_ofx_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28107\,
            in2 => \_gnd_net_\,
            in3 => \N__28092\,
            lcout => \scaler_2.N_1227_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_9_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__28066\,
            in1 => \N__27987\,
            in2 => \_gnd_net_\,
            in3 => \N__27951\,
            lcout => throttle_command_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47316\,
            ce => \N__27918\,
            sr => \N__27876\
        );

    \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__32284\,
            in1 => \N__29044\,
            in2 => \_gnd_net_\,
            in3 => \N__29082\,
            lcout => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__28913\,
            in1 => \N__29551\,
            in2 => \_gnd_net_\,
            in3 => \N__29512\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29007\,
            in2 => \N__27825\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.source_data_1_esr_6_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28226\,
            in2 => \N__29015\,
            in3 => \N__27813\,
            lcout => scaler_3_data_6,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_1\,
            carryout => \scaler_3.un2_source_data_0_cry_2\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_7_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28211\,
            in2 => \N__28230\,
            in3 => \N__28218\,
            lcout => scaler_3_data_7,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_2\,
            carryout => \scaler_3.un2_source_data_0_cry_3\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_8_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28196\,
            in2 => \N__28215\,
            in3 => \N__28203\,
            lcout => scaler_3_data_8,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_3\,
            carryout => \scaler_3.un2_source_data_0_cry_4\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_9_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28181\,
            in2 => \N__28200\,
            in3 => \N__28188\,
            lcout => scaler_3_data_9,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_4\,
            carryout => \scaler_3.un2_source_data_0_cry_5\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_10_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28166\,
            in2 => \N__28185\,
            in3 => \N__28173\,
            lcout => scaler_3_data_10,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_5\,
            carryout => \scaler_3.un2_source_data_0_cry_6\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_11_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28151\,
            in2 => \N__28170\,
            in3 => \N__28158\,
            lcout => scaler_3_data_11,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_6\,
            carryout => \scaler_3.un2_source_data_0_cry_7\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_12_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28139\,
            in2 => \N__28155\,
            in3 => \N__28143\,
            lcout => scaler_3_data_12,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_7\,
            carryout => \scaler_3.un2_source_data_0_cry_8\,
            clk => \N__47305\,
            ce => \N__32403\,
            sr => \N__43847\
        );

    \scaler_3.source_data_1_esr_13_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28140\,
            in2 => \N__28128\,
            in3 => \N__28119\,
            lcout => scaler_3_data_13,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_9\,
            clk => \N__47297\,
            ce => \N__32402\,
            sr => \N__43852\
        );

    \scaler_3.source_data_1_esr_14_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28116\,
            lcout => scaler_3_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => \N__32402\,
            sr => \N__43852\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28899\,
            in2 => \N__28359\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28340\,
            in2 => \N__28909\,
            in3 => \N__28347\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_7_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28325\,
            in2 => \N__28344\,
            in3 => \N__28332\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_8_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28310\,
            in2 => \N__28329\,
            in3 => \N__28317\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_9_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28295\,
            in2 => \N__28314\,
            in3 => \N__28302\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_10_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28280\,
            in2 => \N__28299\,
            in3 => \N__28287\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_11_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28265\,
            in2 => \N__28284\,
            in3 => \N__28272\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_12_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28253\,
            in2 => \N__28269\,
            in3 => \N__28257\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__47290\,
            ce => \N__32401\,
            sr => \N__43858\
        );

    \scaler_4.source_data_1_esr_13_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28254\,
            in2 => \N__28242\,
            in3 => \N__28233\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__47282\,
            ce => \N__32400\,
            sr => \N__43867\
        );

    \scaler_4.source_data_1_esr_14_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28365\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47282\,
            ce => \N__32400\,
            sr => \N__43867\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__41922\,
            in1 => \N__40755\,
            in2 => \_gnd_net_\,
            in3 => \N__42275\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIHB5T_5_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28626\,
            in2 => \_gnd_net_\,
            in3 => \N__28507\,
            lcout => \pid_alt.m21_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIAAPN5_1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__33208\,
            in1 => \N__32942\,
            in2 => \_gnd_net_\,
            in3 => \N__28425\,
            lcout => \pid_alt.un1_reset_1_0_i\,
            ltout => \pid_alt.un1_reset_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIVV066_1_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28362\,
            in3 => \N__33209\,
            lcout => \pid_alt.N_96_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__28520\,
            in1 => \N__33654\,
            in2 => \N__28672\,
            in3 => \N__28401\,
            lcout => \pid_alt.error_i_acummZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__32771\,
            sr => \N__33693\
        );

    \pid_alt.error_i_acumm_esr_1_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__28521\,
            in1 => \N__28388\,
            in2 => \N__28673\,
            in3 => \N__28402\,
            lcout => \pid_alt.error_i_acummZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__32771\,
            sr => \N__33693\
        );

    \pid_alt.error_i_acumm_esr_2_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__28403\,
            in1 => \N__28667\,
            in2 => \N__28527\,
            in3 => \N__28487\,
            lcout => \pid_alt.error_i_acummZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__32771\,
            sr => \N__33693\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIAP1A_13_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__32844\,
            in1 => \N__32795\,
            in2 => \_gnd_net_\,
            in3 => \N__32821\,
            lcout => \pid_alt.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_4_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__28522\,
            in1 => \N__28637\,
            in2 => \N__28674\,
            in3 => \N__33076\,
            lcout => \pid_alt.error_i_acummZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__32771\,
            sr => \N__33693\
        );

    \pid_alt.error_i_acumm_esr_3_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__28404\,
            in1 => \N__28668\,
            in2 => \N__28467\,
            in3 => \N__28523\,
            lcout => \pid_alt.error_i_acummZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__32771\,
            sr => \N__33693\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNICMLK3_2_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28488\,
            in1 => \N__28473\,
            in2 => \N__28466\,
            in3 => \N__28437\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIO7B05_21_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__32852\,
            in1 => \N__28371\,
            in2 => \N__28428\,
            in3 => \N__28573\,
            lcout => \pid_alt.N_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI4SOH2_10_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__28574\,
            in1 => \N__28416\,
            in2 => \N__28683\,
            in3 => \N__33049\,
            lcout => \pid_alt.N_62_mux\,
            ltout => \pid_alt.N_62_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIEPGB3_5_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33050\,
            in1 => \_gnd_net_\,
            in2 => \N__28407\,
            in3 => \N__28636\,
            lcout => \pid_alt.N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI935T_0_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28389\,
            in2 => \_gnd_net_\,
            in3 => \N__33653\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIB9F01_10_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33097\,
            in1 => \N__28696\,
            in2 => \N__28374\,
            in3 => \N__28594\,
            lcout => \pid_alt.m21_e_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_10_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111010"
        )
    port map (
            in0 => \N__33230\,
            in1 => \N__28698\,
            in2 => \N__30354\,
            in3 => \N__33067\,
            lcout => \pid_alt.error_i_acummZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47264\,
            ce => 'H',
            sr => \N__33703\
        );

    \pid_alt.error_i_acumm_8_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__30444\,
            in1 => \N__28734\,
            in2 => \N__33244\,
            in3 => \N__33068\,
            lcout => \pid_alt.error_i_acummZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47264\,
            ce => 'H',
            sr => \N__33703\
        );

    \pid_alt.error_i_acumm_9_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__33069\,
            in1 => \N__33235\,
            in2 => \N__30399\,
            in3 => \N__28717\,
            lcout => \pid_alt.error_i_acummZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47264\,
            ce => 'H',
            sr => \N__33703\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIBO62_10_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28697\,
            lcout => \pid_alt.m35_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_5_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__28660\,
            in1 => \N__29924\,
            in2 => \N__28641\,
            in3 => \N__33231\,
            lcout => \pid_alt.error_i_acummZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47264\,
            ce => 'H',
            sr => \N__33703\
        );

    \pid_alt.error_i_acumm_12_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__33236\,
            in1 => \N__30267\,
            in2 => \N__28602\,
            in3 => \N__28578\,
            lcout => \pid_alt.error_i_acummZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__33718\
        );

    \pid_alt.error_i_acumm_7_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__30494\,
            in1 => \N__33070\,
            in2 => \N__33245\,
            in3 => \N__28560\,
            lcout => \pid_alt.error_i_acummZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__33718\
        );

    \uart_drone.state_RNO_0_0_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__31658\,
            in1 => \N__31372\,
            in2 => \_gnd_net_\,
            in3 => \N__44090\,
            lcout => \uart_drone.state_srsts_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31509\,
            in1 => \N__31773\,
            in2 => \_gnd_net_\,
            in3 => \N__31607\,
            lcout => \uart_pc.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30999\,
            in1 => \N__31072\,
            in2 => \N__28857\,
            in3 => \N__45130\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34832\,
            in2 => \_gnd_net_\,
            in3 => \N__34853\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__33842\,
            in1 => \N__37318\,
            in2 => \N__28881\,
            in3 => \N__33792\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29214\,
            in1 => \N__31220\,
            in2 => \N__28874\,
            in3 => \N__28760\,
            lcout => \uart_pc.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_1_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__28761\,
            in1 => \N__28853\,
            in2 => \N__29205\,
            in3 => \N__31224\,
            lcout => \uart_pc.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_2_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29094\,
            in1 => \N__31221\,
            in2 => \N__28841\,
            in3 => \N__28762\,
            lcout => \uart_pc.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_3_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__28763\,
            in1 => \N__29100\,
            in2 => \N__31019\,
            in3 => \N__31225\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29193\,
            in1 => \N__31222\,
            in2 => \N__28817\,
            in3 => \N__28764\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_5_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__28765\,
            in1 => \N__29088\,
            in2 => \N__28799\,
            in3 => \N__31226\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_6_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__31992\,
            in1 => \N__31223\,
            in2 => \N__28782\,
            in3 => \N__28766\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_7_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__28767\,
            in1 => \N__31227\,
            in2 => \N__29127\,
            in3 => \N__31772\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => 'H',
            sr => \N__29109\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__32031\,
            in1 => \N__32075\,
            in2 => \_gnd_net_\,
            in3 => \N__32123\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__32030\,
            in1 => \N__32074\,
            in2 => \_gnd_net_\,
            in3 => \N__32122\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__32032\,
            in1 => \N__32076\,
            in2 => \_gnd_net_\,
            in3 => \N__32124\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_5_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__29259\,
            in2 => \N__37261\,
            in3 => \N__35218\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__43823\
        );

    \scaler_2.source_data_1_4_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__30566\,
            in1 => \N__29079\,
            in2 => \N__29180\,
            in3 => \N__29051\,
            lcout => scaler_2_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__43823\
        );

    \scaler_3.source_data_1_4_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__30567\,
            in1 => \N__28989\,
            in2 => \N__29156\,
            in3 => \N__28952\,
            lcout => scaler_3_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__43823\
        );

    \scaler_2.source_data_1_esr_5_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32278\,
            in1 => \N__29080\,
            in2 => \_gnd_net_\,
            in3 => \N__29052\,
            lcout => scaler_2_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__32406\,
            sr => \N__43829\
        );

    \scaler_3.source_data_1_esr_5_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29019\,
            in1 => \N__28988\,
            in2 => \_gnd_net_\,
            in3 => \N__28953\,
            lcout => scaler_3_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__32406\,
            sr => \N__43829\
        );

    \scaler_4.source_data_1_esr_5_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28917\,
            in1 => \N__29556\,
            in2 => \_gnd_net_\,
            in3 => \N__29517\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__32406\,
            sr => \N__43829\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32071\,
            in1 => \N__32119\,
            in2 => \_gnd_net_\,
            in3 => \N__32025\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__32120\,
            in1 => \_gnd_net_\,
            in2 => \N__32034\,
            in3 => \N__32072\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32073\,
            in1 => \N__32121\,
            in2 => \_gnd_net_\,
            in3 => \N__32029\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_4_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29181\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.aileron_esr_5_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29163\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.elevator_esr_4_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29157\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.elevator_esr_5_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29139\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.rudder_esr_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29475\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.rudder_esr_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29133\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__36267\,
            sr => \N__43838\
        );

    \ppm_encoder_1.un1_throttle_cry_0_c_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36988\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29296\,
            in2 => \N__42994\,
            in3 => \N__29271\,
            lcout => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_0\,
            carryout => \ppm_encoder_1.un1_throttle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29341\,
            in2 => \_gnd_net_\,
            in3 => \N__29268\,
            lcout => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_1\,
            carryout => \ppm_encoder_1.un1_throttle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35473\,
            in2 => \N__42995\,
            in3 => \N__29265\,
            lcout => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_2\,
            carryout => \ppm_encoder_1.un1_throttle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29392\,
            in2 => \_gnd_net_\,
            in3 => \N__29262\,
            lcout => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_3\,
            carryout => \ppm_encoder_1.un1_throttle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29258\,
            in2 => \_gnd_net_\,
            in3 => \N__29226\,
            lcout => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_4\,
            carryout => \ppm_encoder_1.un1_throttle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42923\,
            in2 => \N__34307\,
            in3 => \N__29223\,
            lcout => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_5\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31892\,
            in2 => \_gnd_net_\,
            in3 => \N__29220\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34223\,
            in2 => \_gnd_net_\,
            in3 => \N__29217\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32588\,
            in2 => \_gnd_net_\,
            in3 => \N__29367\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29435\,
            in2 => \_gnd_net_\,
            in3 => \N__29364\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32723\,
            in2 => \_gnd_net_\,
            in3 => \N__29361\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32492\,
            in2 => \_gnd_net_\,
            in3 => \N__29358\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34460\,
            in2 => \N__43081\,
            in3 => \N__29355\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29352\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => \N__36262\,
            sr => \N__43853\
        );

    \ppm_encoder_1.throttle_2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__37091\,
            in1 => \N__29349\,
            in2 => \N__37631\,
            in3 => \N__29319\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \ppm_encoder_1.pulses2count_16_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__40809\,
            in1 => \N__39773\,
            in2 => \N__39738\,
            in3 => \N__41892\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \ppm_encoder_1.throttle_1_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__29310\,
            in1 => \N__29301\,
            in2 => \N__37148\,
            in3 => \N__34570\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \ppm_encoder_1.rudder_6_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__29790\,
            in1 => \N__37092\,
            in2 => \_gnd_net_\,
            in3 => \N__36205\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \dron_frame_decoder_1.source_data_valid_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__29721\,
            in1 => \N__29676\,
            in2 => \_gnd_net_\,
            in3 => \N__29577\,
            lcout => \debug_CH1_0A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \scaler_4.source_data_1_4_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__30577\,
            in1 => \N__29552\,
            in2 => \N__29474\,
            in3 => \N__29513\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \N__43859\
        );

    \ppm_encoder_1.ppm_output_reg_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001111010000"
        )
    port map (
            in0 => \N__34680\,
            in1 => \N__32868\,
            in2 => \N__29453\,
            in3 => \N__39042\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.rudder_7_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__29766\,
            in1 => \N__29778\,
            in2 => \N__40690\,
            in3 => \N__37102\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.rudder_9_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__29742\,
            in1 => \N__29754\,
            in2 => \N__37150\,
            in3 => \N__40535\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.throttle_10_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__29436\,
            in1 => \N__29418\,
            in2 => \N__32618\,
            in3 => \N__37103\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.elevator_8_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__29817\,
            in1 => \N__29834\,
            in2 => \N__37149\,
            in3 => \N__34241\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.throttle_4_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__29409\,
            in1 => \N__29400\,
            in2 => \N__35374\,
            in3 => \N__37104\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__43868\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29789\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29777\,
            in2 => \_gnd_net_\,
            in3 => \N__29760\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34520\,
            in2 => \_gnd_net_\,
            in3 => \N__29757\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29753\,
            in2 => \_gnd_net_\,
            in3 => \N__29736\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32960\,
            in2 => \_gnd_net_\,
            in3 => \N__29733\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32741\,
            in2 => \_gnd_net_\,
            in3 => \N__29730\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32654\,
            in2 => \_gnd_net_\,
            in3 => \N__29727\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36290\,
            in2 => \N__42885\,
            in3 => \N__29724\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29847\,
            in2 => \_gnd_net_\,
            in3 => \N__29841\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47284\,
            ce => \N__36244\,
            sr => \N__43882\
        );

    \ppm_encoder_1.un1_elevator_cry_6_c_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34356\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31943\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29835\,
            in2 => \_gnd_net_\,
            in3 => \N__29808\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32351\,
            in2 => \_gnd_net_\,
            in3 => \N__29805\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33011\,
            in2 => \_gnd_net_\,
            in3 => \N__29802\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32696\,
            in2 => \_gnd_net_\,
            in3 => \N__29799\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32528\,
            in2 => \_gnd_net_\,
            in3 => \N__29796\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34499\,
            in2 => \N__43020\,
            in3 => \N__29793\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30153\,
            in2 => \_gnd_net_\,
            in3 => \N__30141\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47272\,
            ce => \N__36266\,
            sr => \N__43890\
        );

    \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33665\,
            in2 => \N__39585\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.un1_pid_prereg_0\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30108\,
            in2 => \N__34866\,
            in3 => \N__30048\,
            lcout => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30045\,
            in2 => \N__36729\,
            in3 => \N__30006\,
            lcout => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30003\,
            in2 => \N__39552\,
            in3 => \N__29958\,
            lcout => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29955\,
            in2 => \N__43206\,
            in3 => \N__29928\,
            lcout => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNIT8KA1_5_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45408\,
            in2 => \N__29925\,
            in3 => \N__29883\,
            lcout => \pid_alt.error_i_reg_esr_RNIT8KA1Z0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46215\,
            in2 => \N__33261\,
            in3 => \N__29850\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30498\,
            in2 => \N__46239\,
            in3 => \N__30447\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30443\,
            in2 => \N__45384\,
            in3 => \N__30402\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47616\,
            in2 => \N__30395\,
            in3 => \N__30357\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30350\,
            in2 => \N__44760\,
            in3 => \N__30303\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33026\,
            in2 => \N__44727\,
            in3 => \N__30270\,
            lcout => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI7RNP_12_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30266\,
            in2 => \N__44694\,
            in3 => \N__30222\,
            lcout => \pid_alt.error_i_reg_esr_RNI7RNPZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32784\,
            in2 => \N__45819\,
            in3 => \N__30189\,
            lcout => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47595\,
            in2 => \_gnd_net_\,
            in3 => \N__30156\,
            lcout => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46194\,
            in2 => \_gnd_net_\,
            in3 => \N__30918\,
            lcout => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47511\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47553\,
            in2 => \_gnd_net_\,
            in3 => \N__30849\,
            lcout => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47532\,
            in2 => \_gnd_net_\,
            in3 => \N__30813\,
            lcout => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47496\,
            in2 => \_gnd_net_\,
            in3 => \N__30774\,
            lcout => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47576\,
            in2 => \_gnd_net_\,
            in3 => \N__30726\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30723\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_ctle_14_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30579\,
            in2 => \_gnd_net_\,
            in3 => \N__44071\,
            lcout => \debug_CH3_20A_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_0_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__31244\,
            in1 => \N__31216\,
            in2 => \_gnd_net_\,
            in3 => \N__44101\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__31520\,
            in1 => \N__31278\,
            in2 => \N__31260\,
            in3 => \N__31563\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__33489\,
            in1 => \N__33916\,
            in2 => \N__33885\,
            in3 => \N__44126\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101010101"
        )
    port map (
            in0 => \N__31257\,
            in1 => \N__36616\,
            in2 => \N__31452\,
            in3 => \N__36488\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_1_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__31130\,
            in1 => \N__31230\,
            in2 => \N__31251\,
            in3 => \N__44127\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33508\,
            in2 => \_gnd_net_\,
            in3 => \N__36531\,
            lcout => \uart_drone.N_126_li\,
            ltout => \uart_drone.N_126_li_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__36605\,
            in1 => \N__36483\,
            in2 => \N__31233\,
            in3 => \N__44096\,
            lcout => \uart_drone.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__44097\,
            in1 => \N__31101\,
            in2 => \N__31131\,
            in3 => \N__31212\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__31620\,
            in1 => \N__31519\,
            in2 => \N__31134\,
            in3 => \N__31129\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_3_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__43266\,
            in1 => \N__31073\,
            in2 => \N__31020\,
            in3 => \N__31002\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34755\,
            in2 => \_gnd_net_\,
            in3 => \N__34849\,
            lcout => \reset_module_System.reset6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__44098\,
            in1 => \N__31659\,
            in2 => \N__31301\,
            in3 => \N__31393\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__33480\,
            in1 => \N__33917\,
            in2 => \N__44138\,
            in3 => \N__33870\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__36525\,
            in1 => \N__33510\,
            in2 => \N__36608\,
            in3 => \N__36475\,
            lcout => \uart_drone.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__33462\,
            in1 => \N__33918\,
            in2 => \N__44139\,
            in3 => \N__33871\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110011"
        )
    port map (
            in0 => \N__31619\,
            in1 => \N__31562\,
            in2 => \N__31521\,
            in3 => \N__31723\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__36476\,
            in1 => \N__31448\,
            in2 => \N__33525\,
            in3 => \N__44539\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__33750\,
            in1 => \N__31392\,
            in2 => \N__31302\,
            in3 => \N__44077\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__36537\,
            in1 => \N__36607\,
            in2 => \N__31305\,
            in3 => \N__31300\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__44076\,
            in1 => \N__36484\,
            in2 => \_gnd_net_\,
            in3 => \N__44541\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001011110000"
        )
    port map (
            in0 => \N__31725\,
            in1 => \N__31768\,
            in2 => \N__32130\,
            in3 => \N__31748\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__43830\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32125\,
            lcout => OPEN,
            ltout => \uart_pc.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_2_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__31671\,
            in1 => \N__32033\,
            in2 => \N__31854\,
            in3 => \N__32080\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__43830\
        );

    \uart_pc.bit_Count_1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__31749\,
            in1 => \N__32129\,
            in2 => \N__32082\,
            in3 => \N__31670\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__43830\
        );

    \Commands_frame_decoder.state_RNIBV7S_2_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31828\,
            in2 => \_gnd_net_\,
            in3 => \N__44070\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__33998\,
            in1 => \N__40408\,
            in2 => \N__33981\,
            in3 => \N__41815\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32023\,
            in1 => \N__32117\,
            in2 => \_gnd_net_\,
            in3 => \N__32067\,
            lcout => \uart_pc.N_152\,
            ltout => \uart_pc.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31746\,
            in2 => \N__31728\,
            in3 => \N__31724\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37686\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__32118\,
            in1 => \_gnd_net_\,
            in2 => \N__32081\,
            in3 => \N__32024\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAIVN2_7_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31969\,
            in1 => \N__35784\,
            in2 => \N__31920\,
            in3 => \N__35697\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIJII96_7_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35319\,
            in2 => \N__31980\,
            in3 => \N__40251\,
            lcout => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40135\,
            in1 => \N__35338\,
            in2 => \_gnd_net_\,
            in3 => \N__31918\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31970\,
            in1 => \_gnd_net_\,
            in2 => \N__31977\,
            in3 => \N__38925\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__35568\,
            in1 => \N__35582\,
            in2 => \N__31974\,
            in3 => \N__37089\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47364\,
            ce => 'H',
            sr => \N__43848\
        );

    \ppm_encoder_1.elevator_7_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__31919\,
            in1 => \N__31956\,
            in2 => \N__37147\,
            in3 => \N__31944\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47364\,
            ce => 'H',
            sr => \N__43848\
        );

    \ppm_encoder_1.throttle_7_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__31905\,
            in1 => \N__35339\,
            in2 => \N__31899\,
            in3 => \N__37090\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47364\,
            ce => 'H',
            sr => \N__43848\
        );

    \scaler_2.un2_source_data_0_cry_1_c_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32285\,
            in2 => \N__32301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_6_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32252\,
            in2 => \N__32289\,
            in3 => \N__32259\,
            lcout => scaler_2_data_6,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_1\,
            carryout => \scaler_2.un2_source_data_0_cry_2\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_7_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32231\,
            in2 => \N__32256\,
            in3 => \N__32238\,
            lcout => scaler_2_data_7,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_2\,
            carryout => \scaler_2.un2_source_data_0_cry_3\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_8_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32210\,
            in2 => \N__32235\,
            in3 => \N__32217\,
            lcout => scaler_2_data_8,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_3\,
            carryout => \scaler_2.un2_source_data_0_cry_4\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_9_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32189\,
            in2 => \N__32214\,
            in3 => \N__32196\,
            lcout => scaler_2_data_9,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_4\,
            carryout => \scaler_2.un2_source_data_0_cry_5\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_10_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32168\,
            in2 => \N__32193\,
            in3 => \N__32175\,
            lcout => scaler_2_data_10,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_5\,
            carryout => \scaler_2.un2_source_data_0_cry_6\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_11_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32147\,
            in2 => \N__32172\,
            in3 => \N__32154\,
            lcout => scaler_2_data_11,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_6\,
            carryout => \scaler_2.un2_source_data_0_cry_7\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_12_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32450\,
            in2 => \N__32151\,
            in3 => \N__32133\,
            lcout => scaler_2_data_12,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_7\,
            carryout => \scaler_2.un2_source_data_0_cry_8\,
            clk => \N__47349\,
            ce => \N__32405\,
            sr => \N__43854\
        );

    \scaler_2.source_data_1_esr_13_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32451\,
            in2 => \N__32427\,
            in3 => \N__32412\,
            lcout => scaler_2_data_13,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_9\,
            clk => \N__47332\,
            ce => \N__32404\,
            sr => \N__43860\
        );

    \scaler_2.source_data_1_esr_14_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32409\,
            lcout => scaler_2_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47332\,
            ce => \N__32404\,
            sr => \N__43860\
        );

    \ppm_encoder_1.throttle_RNIU7KK2_9_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__40531\,
            in1 => \N__35286\,
            in2 => \N__32571\,
            in3 => \N__37581\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNITSI96_9_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__40574\,
            in1 => \_gnd_net_\,
            in2 => \N__32379\,
            in3 => \N__32376\,
            lcout => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIEMVN2_9_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__35801\,
            in1 => \N__32365\,
            in2 => \N__32316\,
            in3 => \N__35731\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40127\,
            in1 => \N__32569\,
            in2 => \_gnd_net_\,
            in3 => \N__32314\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__38945\,
            in1 => \_gnd_net_\,
            in2 => \N__32370\,
            in3 => \N__32366\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_9_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__32367\,
            in1 => \N__36014\,
            in2 => \N__37242\,
            in3 => \N__35997\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => 'H',
            sr => \N__43869\
        );

    \ppm_encoder_1.elevator_9_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__32315\,
            in1 => \N__37193\,
            in2 => \N__32355\,
            in3 => \N__32328\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => 'H',
            sr => \N__43869\
        );

    \ppm_encoder_1.throttle_9_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32595\,
            in1 => \N__32577\,
            in2 => \N__37243\,
            in3 => \N__32570\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => 'H',
            sr => \N__43869\
        );

    \ppm_encoder_1.throttle_RNII6JI2_12_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37582\,
            in1 => \N__32635\,
            in2 => \N__34064\,
            in3 => \N__35288\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFQRT5_12_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__38096\,
            in1 => \_gnd_net_\,
            in2 => \N__32556\,
            in3 => \N__32553\,
            lcout => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI25DH2_12_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__32542\,
            in1 => \N__35818\,
            in2 => \N__34040\,
            in3 => \N__35733\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32543\,
            in1 => \N__38983\,
            in2 => \_gnd_net_\,
            in3 => \N__34020\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__35946\,
            in1 => \N__35922\,
            in2 => \N__32547\,
            in3 => \N__37191\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47309\,
            ce => 'H',
            sr => \N__43876\
        );

    \ppm_encoder_1.elevator_12_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__34036\,
            in1 => \N__32529\,
            in2 => \N__37241\,
            in3 => \N__32505\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47309\,
            ce => 'H',
            sr => \N__43876\
        );

    \ppm_encoder_1.throttle_12_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__32493\,
            in1 => \N__37192\,
            in2 => \N__32463\,
            in3 => \N__34060\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47309\,
            ce => 'H',
            sr => \N__43876\
        );

    \ppm_encoder_1.throttle_RNIG4JI2_11_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__34600\,
            in1 => \N__35287\,
            in2 => \N__34632\,
            in3 => \N__37591\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_11_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__37233\,
            in1 => \N__32754\,
            in2 => \N__34605\,
            in3 => \N__32748\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47299\,
            ce => 'H',
            sr => \N__43883\
        );

    \ppm_encoder_1.throttle_11_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__34630\,
            in1 => \N__37232\,
            in2 => \N__32730\,
            in3 => \N__32706\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47299\,
            ce => 'H',
            sr => \N__43883\
        );

    \ppm_encoder_1.elevator_11_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__32697\,
            in1 => \N__32673\,
            in2 => \N__34928\,
            in3 => \N__37231\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47299\,
            ce => 'H',
            sr => \N__43883\
        );

    \ppm_encoder_1.rudder_12_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__32637\,
            in1 => \N__32661\,
            in2 => \N__37258\,
            in3 => \N__32643\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47299\,
            ce => 'H',
            sr => \N__43883\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40928\,
            in1 => \N__37740\,
            in2 => \_gnd_net_\,
            in3 => \N__32636\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__41141\,
            in1 => \_gnd_net_\,
            in2 => \N__32622\,
            in3 => \N__35532\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIU0DH2_10_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__34735\,
            in1 => \N__35814\,
            in2 => \N__32982\,
            in3 => \N__35732\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIE2JI2_10_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__35848\,
            in1 => \N__35285\,
            in2 => \N__32619\,
            in3 => \N__37590\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40128\,
            in1 => \N__32617\,
            in2 => \_gnd_net_\,
            in3 => \N__32980\,
            lcout => \ppm_encoder_1.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_10_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__32981\,
            in1 => \N__33015\,
            in2 => \N__37260\,
            in3 => \N__32988\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47291\,
            ce => 'H',
            sr => \N__43886\
        );

    \ppm_encoder_1.aileron_10_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__34736\,
            in1 => \N__35985\,
            in2 => \N__37259\,
            in3 => \N__35964\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47291\,
            ce => 'H',
            sr => \N__43886\
        );

    \ppm_encoder_1.rudder_10_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__32967\,
            in1 => \N__32949\,
            in2 => \N__35858\,
            in3 => \N__37240\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47291\,
            ce => 'H',
            sr => \N__43886\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__40300\,
            in1 => \N__34711\,
            in2 => \N__32943\,
            in3 => \N__44665\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34671\,
            in2 => \_gnd_net_\,
            in3 => \N__40299\,
            lcout => \ppm_encoder_1.PPM_STATE_59_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__40301\,
            in1 => \N__34712\,
            in2 => \N__34679\,
            in3 => \N__44666\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47285\,
            ce => 'H',
            sr => \N__43891\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__40302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34713\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47285\,
            ce => 'H',
            sr => \N__43891\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34893\,
            in1 => \N__34722\,
            in2 => \N__34701\,
            in3 => \N__39642\,
            lcout => \ppm_encoder_1.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_13_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__32856\,
            in1 => \N__32826\,
            in2 => \_gnd_net_\,
            in3 => \N__32799\,
            lcout => \pid_alt.error_i_acummZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => \N__32775\,
            sr => \N__33719\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__41771\,
            in1 => \N__42276\,
            in2 => \_gnd_net_\,
            in3 => \N__37764\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37763\,
            in1 => \_gnd_net_\,
            in2 => \N__42291\,
            in3 => \N__41775\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__41772\,
            in1 => \N__42277\,
            in2 => \_gnd_net_\,
            in3 => \N__37739\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_12_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37738\,
            in1 => \_gnd_net_\,
            in2 => \N__42290\,
            in3 => \N__41774\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.N_1330_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37712\,
            in2 => \_gnd_net_\,
            in3 => \N__41770\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_6_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33440\,
            in2 => \_gnd_net_\,
            in3 => \N__46681\,
            lcout => alt_ki_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47273\,
            ce => \N__44828\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_6_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__33260\,
            in1 => \N__33282\,
            in2 => \N__33246\,
            in3 => \N__33078\,
            lcout => \pid_alt.error_i_acummZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => 'H',
            sr => \N__33720\
        );

    \pid_alt.error_i_acumm_11_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__33240\,
            in1 => \N__33027\,
            in2 => \N__33105\,
            in3 => \N__33077\,
            lcout => \pid_alt.error_i_acummZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => 'H',
            sr => \N__33720\
        );

    \pid_alt.error_i_acumm_prereg_esr_0_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39581\,
            in2 => \_gnd_net_\,
            in3 => \N__33672\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47266\,
            ce => \N__33627\,
            sr => \N__43899\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__33954\,
            in1 => \N__33929\,
            in2 => \N__33957\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33509\,
            in2 => \_gnd_net_\,
            in3 => \N__33483\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36544\,
            in2 => \_gnd_net_\,
            in3 => \N__33468\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36615\,
            in2 => \_gnd_net_\,
            in3 => \N__33465\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__33956\,
            in1 => \N__33914\,
            in2 => \N__33884\,
            in3 => \N__44122\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__37317\,
            in1 => \N__34779\,
            in2 => \N__33841\,
            in3 => \N__33787\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34988\,
            in1 => \N__35003\,
            in2 => \N__34974\,
            in3 => \N__35033\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35105\,
            in1 => \N__35088\,
            in2 => \N__33450\,
            in3 => \N__33447\,
            lcout => \reset_module_System.reset6_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33955\,
            in2 => \_gnd_net_\,
            in3 => \N__33930\,
            lcout => OPEN,
            ltout => \uart_drone.timer_Count_RNO_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__33869\,
            in1 => \N__33915\,
            in2 => \N__33933\,
            in3 => \N__44128\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__44538\,
            in1 => \N__33913\,
            in2 => \N__36714\,
            in3 => \N__44123\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__44537\,
            in1 => \N__36604\,
            in2 => \N__33752\,
            in3 => \N__36535\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35019\,
            in1 => \N__34770\,
            in2 => \N__35067\,
            in3 => \N__34791\,
            lcout => \reset_module_System.reset6_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34831\,
            in1 => \N__34947\,
            in2 => \N__35145\,
            in3 => \N__33801\,
            lcout => \reset_module_System.reset6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36671\,
            in1 => \N__39496\,
            in2 => \_gnd_net_\,
            in3 => \N__44391\,
            lcout => \uart_drone.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__44540\,
            in1 => \N__36606\,
            in2 => \N__33753\,
            in3 => \N__36536\,
            lcout => OPEN,
            ltout => \uart_drone.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__33751\,
            in1 => \N__36710\,
            in2 => \N__33723\,
            in3 => \N__44124\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__36677\,
            in1 => \N__39512\,
            in2 => \_gnd_net_\,
            in3 => \N__44405\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__44406\,
            in1 => \_gnd_net_\,
            in2 => \N__39519\,
            in3 => \N__36678\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__34008\,
            in1 => \N__44110\,
            in2 => \N__40926\,
            in3 => \N__42009\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40131\,
            in1 => \N__34068\,
            in2 => \_gnd_net_\,
            in3 => \N__34044\,
            lcout => \ppm_encoder_1.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111010"
        )
    port map (
            in0 => \N__33999\,
            in1 => \N__42167\,
            in2 => \N__44136\,
            in3 => \N__41947\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__41945\,
            in1 => \N__38917\,
            in2 => \N__33980\,
            in3 => \N__44116\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__40134\,
            in1 => \N__40888\,
            in2 => \N__38946\,
            in3 => \N__42166\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__41946\,
            in1 => \N__44112\,
            in2 => \N__34002\,
            in3 => \N__35310\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33997\,
            in1 => \N__35129\,
            in2 => \N__33979\,
            in3 => \N__35309\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34113\,
            in3 => \N__41943\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__41944\,
            in1 => \N__44111\,
            in2 => \N__40377\,
            in3 => \N__38916\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIS5KK2_8_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__38401\,
            in1 => \N__35267\,
            in2 => \N__34188\,
            in3 => \N__37552\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35308\,
            lcout => \ppm_encoder_1.N_227\,
            ltout => \ppm_encoder_1.N_227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__34100\,
            in1 => \_gnd_net_\,
            in2 => \N__34110\,
            in3 => \N__42114\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__42008\,
            in1 => \_gnd_net_\,
            in2 => \N__34107\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__35780\,
            in1 => \N__34139\,
            in2 => \N__34166\,
            in3 => \N__35684\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110000000"
        )
    port map (
            in0 => \N__40136\,
            in1 => \N__40958\,
            in2 => \N__38971\,
            in3 => \N__39981\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__35683\,
            in2 => \N__34104\,
            in3 => \N__42007\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIALN65_1_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001111"
        )
    port map (
            in0 => \N__37553\,
            in1 => \N__34577\,
            in2 => \N__34092\,
            in3 => \N__37973\,
            lcout => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40472\,
            in1 => \N__40407\,
            in2 => \N__40378\,
            in3 => \N__41923\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__35378\,
            in2 => \_gnd_net_\,
            in3 => \N__40373\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38918\,
            in2 => \N__34146\,
            in3 => \N__34143\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__40471\,
            in1 => \N__40406\,
            in2 => \N__40379\,
            in3 => \N__41924\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIO1KK2_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__34276\,
            in1 => \N__36212\,
            in2 => \N__34125\,
            in3 => \N__35268\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__35269\,
            in1 => \N__41021\,
            in2 => \N__35649\,
            in3 => \N__37568\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8GVN2_6_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__34366\,
            in1 => \N__35783\,
            in2 => \N__34335\,
            in3 => \N__35730\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEDI96_6_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__37787\,
            in1 => \_gnd_net_\,
            in2 => \N__34122\,
            in3 => \N__34119\,
            lcout => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40114\,
            in1 => \N__34277\,
            in2 => \_gnd_net_\,
            in3 => \N__34333\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__34367\,
            in1 => \_gnd_net_\,
            in2 => \N__34371\,
            in3 => \N__38949\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__37250\,
            in1 => \N__35600\,
            in2 => \_gnd_net_\,
            in3 => \N__34368\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => 'H',
            sr => \N__43870\
        );

    \ppm_encoder_1.elevator_6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__34355\,
            in2 => \_gnd_net_\,
            in3 => \N__37254\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => 'H',
            sr => \N__43870\
        );

    \ppm_encoder_1.throttle_6_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__34320\,
            in1 => \N__34308\,
            in2 => \N__37263\,
            in3 => \N__34278\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => 'H',
            sr => \N__43870\
        );

    \ppm_encoder_1.elevator_RNICKVN2_8_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__35800\,
            in2 => \N__34251\,
            in3 => \N__35734\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIONI96_8_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__40623\,
            in1 => \_gnd_net_\,
            in2 => \N__34263\,
            in3 => \N__34260\,
            lcout => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__34183\,
            in2 => \_gnd_net_\,
            in3 => \N__34250\,
            lcout => \ppm_encoder_1.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_8_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__34227\,
            in1 => \N__34200\,
            in2 => \N__37256\,
            in3 => \N__34184\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47333\,
            ce => 'H',
            sr => \N__43877\
        );

    \ppm_encoder_1.aileron_8_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__38801\,
            in1 => \N__37214\,
            in2 => \N__36027\,
            in3 => \N__36047\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47333\,
            ce => 'H',
            sr => \N__43877\
        );

    \ppm_encoder_1.rudder_8_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__34542\,
            in1 => \N__34527\,
            in2 => \N__37255\,
            in3 => \N__38405\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47333\,
            ce => 'H',
            sr => \N__43877\
        );

    \ppm_encoder_1.throttle_RNIK8JI2_13_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__39001\,
            in1 => \N__35289\,
            in2 => \N__34425\,
            in3 => \N__37583\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKVRT5_13_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38045\,
            in2 => \N__34509\,
            in3 => \N__34506\,
            lcout => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI47DH2_13_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__34384\,
            in1 => \N__35819\,
            in2 => \N__34407\,
            in3 => \N__35744\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_13_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__35883\,
            in1 => \N__34385\,
            in2 => \N__35907\,
            in3 => \N__37224\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47320\,
            ce => 'H',
            sr => \N__43884\
        );

    \ppm_encoder_1.elevator_13_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__34405\,
            in1 => \N__34500\,
            in2 => \N__37257\,
            in3 => \N__34476\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47320\,
            ce => 'H',
            sr => \N__43884\
        );

    \ppm_encoder_1.throttle_13_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__34464\,
            in1 => \N__34423\,
            in2 => \N__34440\,
            in3 => \N__37225\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47320\,
            ce => 'H',
            sr => \N__43884\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40125\,
            in1 => \N__34424\,
            in2 => \_gnd_net_\,
            in3 => \N__34406\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38974\,
            in2 => \N__34389\,
            in3 => \N__34386\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40126\,
            in1 => \N__34631\,
            in2 => \_gnd_net_\,
            in3 => \N__34921\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38973\,
            in2 => \N__34614\,
            in3 => \N__36148\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNISFRP_13_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41332\,
            in1 => \N__42233\,
            in2 => \_gnd_net_\,
            in3 => \N__41840\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIALRT5_11_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__38144\,
            in1 => \N__34611\,
            in2 => \_gnd_net_\,
            in3 => \N__34902\,
            lcout => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34601\,
            in1 => \N__40927\,
            in2 => \_gnd_net_\,
            in3 => \N__37762\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41148\,
            in2 => \N__34584\,
            in3 => \N__35527\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111100"
        )
    port map (
            in0 => \N__42234\,
            in1 => \N__40454\,
            in2 => \N__44137\,
            in3 => \N__41777\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__40092\,
            in1 => \_gnd_net_\,
            in2 => \N__38984\,
            in3 => \N__37630\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__34581\,
            in1 => \N__40091\,
            in2 => \_gnd_net_\,
            in3 => \N__38976\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38975\,
            in1 => \N__34548\,
            in2 => \_gnd_net_\,
            in3 => \N__34737\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__34638\,
            in1 => \N__42445\,
            in2 => \N__34647\,
            in3 => \N__39263\,
            lcout => \ppm_encoder_1.N_145_17\,
            ltout => \ppm_encoder_1.N_145_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34892\,
            in1 => \N__39641\,
            in2 => \N__34716\,
            in3 => \N__34653\,
            lcout => \ppm_encoder_1.N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__36371\,
            in1 => \N__39356\,
            in2 => \N__40321\,
            in3 => \N__39385\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI5GRT5_10_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__39030\,
            in1 => \N__34692\,
            in2 => \_gnd_net_\,
            in3 => \N__34686\,
            lcout => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44084\,
            in2 => \_gnd_net_\,
            in3 => \N__41814\,
            lcout => \ppm_encoder_1.N_1330_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39355\,
            in1 => \N__36370\,
            in2 => \N__39387\,
            in3 => \N__34675\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42706\,
            in1 => \N__36320\,
            in2 => \N__42741\,
            in3 => \N__36341\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__36081\,
            in1 => \N__36369\,
            in2 => \N__36393\,
            in3 => \N__36057\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39245\,
            in2 => \_gnd_net_\,
            in3 => \N__42484\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__40055\,
            in1 => \N__44118\,
            in2 => \N__38985\,
            in3 => \N__41776\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI03DH2_11_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__36153\,
            in1 => \N__35820\,
            in2 => \N__34929\,
            in3 => \N__35745\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__36391\,
            in1 => \N__44620\,
            in2 => \N__39294\,
            in3 => \N__44584\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_1_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34881\,
            lcout => \pid_alt.error_i_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47277\,
            ce => \N__46797\,
            sr => \N__46593\
        );

    \reset_module_System.count_1_cry_1_c_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34854\,
            in2 => \N__34833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34790\,
            in2 => \_gnd_net_\,
            in3 => \N__34773\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34769\,
            in2 => \_gnd_net_\,
            in3 => \N__34758\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34754\,
            in2 => \_gnd_net_\,
            in3 => \N__34740\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35034\,
            in2 => \_gnd_net_\,
            in3 => \N__35022\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35018\,
            in2 => \_gnd_net_\,
            in3 => \N__35007\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35004\,
            in2 => \_gnd_net_\,
            in3 => \N__34992\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34989\,
            in2 => \_gnd_net_\,
            in3 => \N__34977\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34970\,
            in2 => \_gnd_net_\,
            in3 => \N__34956\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37331\,
            in2 => \_gnd_net_\,
            in3 => \N__34953\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37370\,
            in2 => \_gnd_net_\,
            in3 => \N__34950\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34946\,
            in2 => \_gnd_net_\,
            in3 => \N__34935\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35157\,
            in2 => \_gnd_net_\,
            in3 => \N__34932\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37358\,
            in2 => \_gnd_net_\,
            in3 => \N__35112\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35181\,
            in2 => \_gnd_net_\,
            in3 => \N__35109\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35106\,
            in2 => \_gnd_net_\,
            in3 => \N__35094\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__47437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37343\,
            in2 => \_gnd_net_\,
            in3 => \N__35091\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35087\,
            in2 => \_gnd_net_\,
            in3 => \N__35073\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35046\,
            in3 => \N__35070\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35066\,
            in2 => \_gnd_net_\,
            in3 => \N__35052\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35049\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35042\,
            in1 => \N__35180\,
            in2 => \N__35169\,
            in3 => \N__35156\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35222\,
            in1 => \N__35408\,
            in2 => \_gnd_net_\,
            in3 => \N__40362\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38860\,
            in2 => \N__35136\,
            in3 => \N__35430\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40363\,
            in1 => \N__40490\,
            in2 => \N__40929\,
            in3 => \N__39993\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_159_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__42038\,
            in1 => \_gnd_net_\,
            in2 => \N__35133\,
            in3 => \N__37704\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__41978\,
            in1 => \N__36941\,
            in2 => \N__37703\,
            in3 => \N__42337\,
            lcout => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__40132\,
            in1 => \N__38857\,
            in2 => \_gnd_net_\,
            in3 => \N__36965\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__44108\,
            in1 => \N__35130\,
            in2 => \N__35196\,
            in3 => \N__41977\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__38858\,
            in1 => \N__40133\,
            in2 => \_gnd_net_\,
            in3 => \N__35451\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001110"
        )
    port map (
            in0 => \N__41976\,
            in1 => \N__44109\,
            in2 => \N__42231\,
            in3 => \N__38859\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37687\,
            in2 => \_gnd_net_\,
            in3 => \N__41975\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__39975\,
            in1 => \N__40130\,
            in2 => \_gnd_net_\,
            in3 => \N__40485\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__41122\,
            in1 => \N__40909\,
            in2 => \N__35385\,
            in3 => \N__37386\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__37454\,
            in1 => \N__35249\,
            in2 => \N__35382\,
            in3 => \N__37550\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37865\,
            in2 => \N__35349\,
            in3 => \N__35346\,
            lcout => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__40691\,
            in1 => \N__35250\,
            in2 => \N__35340\,
            in3 => \N__37551\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35307\,
            in2 => \_gnd_net_\,
            in3 => \N__39974\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__37412\,
            in1 => \N__35248\,
            in2 => \N__35226\,
            in3 => \N__37549\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__42002\,
            in1 => \N__44117\,
            in2 => \N__39991\,
            in3 => \N__35192\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_3_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41611\,
            in1 => \N__39867\,
            in2 => \N__41444\,
            in3 => \N__37887\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47376\,
            ce => 'H',
            sr => \N__43871\
        );

    \ppm_encoder_1.throttle_RNIT9352_3_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010011001"
        )
    port map (
            in0 => \N__35549\,
            in1 => \N__42327\,
            in2 => \N__35450\,
            in3 => \N__37548\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI82223_3_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35553\,
            in3 => \N__37898\,
            lcout => \ppm_encoder_1.throttle_RNI82223Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__35547\,
            in1 => \N__42151\,
            in2 => \_gnd_net_\,
            in3 => \N__41995\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__41996\,
            in1 => \_gnd_net_\,
            in2 => \N__42228\,
            in3 => \N__35548\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__41124\,
            in1 => \N__35550\,
            in2 => \N__35531\,
            in3 => \N__40948\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__37653\,
            in1 => \N__41123\,
            in2 => \N__40977\,
            in3 => \N__35523\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_3_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__35446\,
            in1 => \N__35490\,
            in2 => \N__37262\,
            in3 => \N__35478\,
            lcout => \ppm_encoder_1.throttleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47376\,
            ce => 'H',
            sr => \N__43871\
        );

    \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__35429\,
            in1 => \N__35781\,
            in2 => \N__35409\,
            in3 => \N__35728\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__37833\,
            in1 => \_gnd_net_\,
            in2 => \N__35832\,
            in3 => \N__35829\,
            lcout => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38373\,
            in1 => \N__35782\,
            in2 => \N__35625\,
            in3 => \N__35729\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__41190\,
            in1 => \_gnd_net_\,
            in2 => \N__35658\,
            in3 => \N__35655\,
            lcout => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIANUS_2_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__37650\,
            in1 => \N__42172\,
            in2 => \_gnd_net_\,
            in3 => \N__41993\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35645\,
            in1 => \N__40121\,
            in2 => \_gnd_net_\,
            in3 => \N__35624\,
            lcout => \ppm_encoder_1.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42171\,
            in2 => \_gnd_net_\,
            in3 => \N__41992\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIERUS_6_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__41994\,
            in1 => \_gnd_net_\,
            in2 => \N__42232\,
            in3 => \N__37486\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_c_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35604\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35586\,
            in2 => \_gnd_net_\,
            in3 => \N__35556\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36048\,
            in2 => \_gnd_net_\,
            in3 => \N__36018\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36015\,
            in2 => \_gnd_net_\,
            in3 => \N__35988\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35984\,
            in2 => \_gnd_net_\,
            in3 => \N__35952\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36185\,
            in2 => \_gnd_net_\,
            in3 => \N__35949\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35945\,
            in2 => \_gnd_net_\,
            in3 => \N__35910\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35906\,
            in2 => \N__43050\,
            in3 => \N__35877\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35874\,
            in2 => \_gnd_net_\,
            in3 => \N__35862\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => \N__36227\,
            sr => \N__43887\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__41145\,
            in1 => \N__41247\,
            in2 => \N__40991\,
            in3 => \N__35859\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_13_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__36294\,
            in1 => \N__36279\,
            in2 => \N__37227\,
            in3 => \N__39005\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__43892\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37165\,
            in2 => \_gnd_net_\,
            in3 => \N__44074\,
            lcout => \ppm_encoder_1.pid_altitude_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__40982\,
            in1 => \N__37494\,
            in2 => \N__36216\,
            in3 => \N__41146\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_11_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__36186\,
            in1 => \N__36162\,
            in2 => \N__37226\,
            in3 => \N__36149\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__43892\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36117\,
            in1 => \N__36319\,
            in2 => \N__36099\,
            in3 => \N__36340\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__37440\,
            in1 => \_gnd_net_\,
            in2 => \N__42617\,
            in3 => \N__36129\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => \N__42540\,
            sr => \N__43894\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36111\,
            in1 => \N__42603\,
            in2 => \_gnd_net_\,
            in3 => \N__37398\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => \N__42540\,
            sr => \N__43894\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42598\,
            in1 => \N__36090\,
            in2 => \_gnd_net_\,
            in3 => \N__36921\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => \N__42540\,
            sr => \N__43894\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42599\,
            in1 => \N__36072\,
            in2 => \_gnd_net_\,
            in3 => \N__36066\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => \N__42540\,
            sr => \N__43894\
        );

    \ppm_encoder_1.counter_0_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36392\,
            in2 => \N__36417\,
            in3 => \N__36416\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_1_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36372\,
            in2 => \_gnd_net_\,
            in3 => \N__36351\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_2_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39357\,
            in2 => \_gnd_net_\,
            in3 => \N__36348\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_3_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39386\,
            in2 => \_gnd_net_\,
            in3 => \N__36345\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_4_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36342\,
            in2 => \_gnd_net_\,
            in3 => \N__36324\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_5_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36321\,
            in2 => \_gnd_net_\,
            in3 => \N__36303\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_6_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42708\,
            in2 => \_gnd_net_\,
            in3 => \N__36300\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_7_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42740\,
            in2 => \_gnd_net_\,
            in3 => \N__36297\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__47301\,
            ce => 'H',
            sr => \N__36903\
        );

    \ppm_encoder_1.counter_8_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39264\,
            in2 => \_gnd_net_\,
            in3 => \N__36447\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_9_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39293\,
            in2 => \_gnd_net_\,
            in3 => \N__36444\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_10_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44585\,
            in2 => \_gnd_net_\,
            in3 => \N__36441\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_11_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44621\,
            in2 => \_gnd_net_\,
            in3 => \N__36438\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_12_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42446\,
            in2 => \_gnd_net_\,
            in3 => \N__36435\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_13_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42485\,
            in2 => \_gnd_net_\,
            in3 => \N__36432\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_14_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39246\,
            in2 => \_gnd_net_\,
            in3 => \N__36429\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_15_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39699\,
            in2 => \_gnd_net_\,
            in3 => \N__36426\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__47292\,
            ce => 'H',
            sr => \N__36902\
        );

    \ppm_encoder_1.counter_16_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39659\,
            in2 => \_gnd_net_\,
            in3 => \N__36423\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__47287\,
            ce => 'H',
            sr => \N__36901\
        );

    \ppm_encoder_1.counter_17_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39682\,
            in2 => \_gnd_net_\,
            in3 => \N__36420\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__47287\,
            ce => 'H',
            sr => \N__36901\
        );

    \ppm_encoder_1.counter_18_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39612\,
            in2 => \_gnd_net_\,
            in3 => \N__36906\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => 'H',
            sr => \N__36901\
        );

    \Commands_frame_decoder.source_alt_ki_2_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36887\,
            in2 => \_gnd_net_\,
            in3 => \N__46678\,
            lcout => alt_ki_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47278\,
            ce => \N__44849\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_2_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36738\,
            lcout => \pid_alt.error_i_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47274\,
            ce => \N__46795\,
            sr => \N__46586\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__44461\,
            in1 => \N__36618\,
            in2 => \_gnd_net_\,
            in3 => \N__36549\,
            lcout => \uart_drone.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__39537\,
            in1 => \N__39495\,
            in2 => \N__36686\,
            in3 => \N__39531\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => 'H',
            sr => \N__43839\
        );

    \uart_drone.state_RNI62411_4_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__36617\,
            in1 => \N__36545\,
            in2 => \N__44552\,
            in3 => \N__36489\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => \uart_drone.un1_state_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI63LK2_3_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44548\,
            in2 => \N__36450\,
            in3 => \N__44451\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000110011"
        )
    port map (
            in0 => \N__36966\,
            in1 => \N__38000\,
            in2 => \_gnd_net_\,
            in3 => \N__37596\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37371\,
            in1 => \N__37359\,
            in2 => \N__37347\,
            in3 => \N__37332\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__42035\,
            in1 => \N__37713\,
            in2 => \N__36945\,
            in3 => \N__42348\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__41615\,
            in1 => \N__37275\,
            in2 => \N__37269\,
            in3 => \N__41380\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__43855\
        );

    \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__36939\,
            in1 => \N__42229\,
            in2 => \_gnd_net_\,
            in3 => \N__42034\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => \ppm_encoder_1.un1_init_pulses_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIN3352_0_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36963\,
            in2 => \N__37266\,
            in3 => \N__37592\,
            lcout => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_0_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__36964\,
            in1 => \N__37203\,
            in2 => \_gnd_net_\,
            in3 => \N__36996\,
            lcout => \ppm_encoder_1.throttleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__43855\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__41062\,
            in1 => \_gnd_net_\,
            in2 => \N__40930\,
            in3 => \N__36940\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_4_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__39846\,
            in1 => \N__41616\,
            in2 => \N__41411\,
            in3 => \N__37851\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47417\,
            ce => 'H',
            sr => \N__43861\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__42162\,
            in1 => \N__37469\,
            in2 => \_gnd_net_\,
            in3 => \N__41984\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_4_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37468\,
            in1 => \_gnd_net_\,
            in2 => \N__42037\,
            in3 => \N__42164\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__41063\,
            in1 => \N__37470\,
            in2 => \N__40983\,
            in3 => \N__37458\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_5_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__39831\,
            in1 => \N__41617\,
            in2 => \N__41412\,
            in3 => \N__37809\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47417\,
            ce => 'H',
            sr => \N__43861\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__42165\,
            in1 => \N__41991\,
            in2 => \_gnd_net_\,
            in3 => \N__37426\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37427\,
            in1 => \_gnd_net_\,
            in2 => \N__42036\,
            in3 => \N__42163\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__41064\,
            in1 => \N__37428\,
            in2 => \N__40984\,
            in3 => \N__37416\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_1_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__41423\,
            in1 => \N__39924\,
            in2 => \N__37953\,
            in3 => \N__41606\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47407\,
            ce => 'H',
            sr => \N__43872\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__37384\,
            in1 => \_gnd_net_\,
            in2 => \N__42230\,
            in3 => \N__41998\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__41997\,
            in1 => \N__42158\,
            in2 => \_gnd_net_\,
            in3 => \N__37385\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__40221\,
            in1 => \N__41419\,
            in2 => \N__41619\,
            in3 => \N__38175\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47407\,
            ce => 'H',
            sr => \N__43872\
        );

    \ppm_encoder_1.init_pulses_11_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__40194\,
            in1 => \N__41602\,
            in2 => \N__41446\,
            in3 => \N__38124\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47407\,
            ce => 'H',
            sr => \N__43872\
        );

    \ppm_encoder_1.init_pulses_12_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41601\,
            in1 => \N__40173\,
            in2 => \N__41447\,
            in3 => \N__38076\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47407\,
            ce => 'H',
            sr => \N__43872\
        );

    \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__37652\,
            in1 => \N__42324\,
            in2 => \N__37719\,
            in3 => \N__42003\,
            lcout => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__42325\,
            in1 => \N__37487\,
            in2 => \N__42039\,
            in3 => \N__37717\,
            lcout => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__37718\,
            in1 => \N__42326\,
            in2 => \N__42047\,
            in3 => \N__41337\,
            lcout => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_2_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41595\,
            in1 => \N__39894\,
            in2 => \N__41448\,
            in3 => \N__37917\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => 'H',
            sr => \N__43878\
        );

    \ppm_encoder_1.throttle_RNIR7352_2_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__37651\,
            in1 => \N__42323\,
            in2 => \N__37632\,
            in3 => \N__37574\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI5V123_2_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37497\,
            in3 => \N__37928\,
            lcout => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_6_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__39792\,
            in1 => \N__41445\,
            in2 => \N__41618\,
            in3 => \N__37773\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => 'H',
            sr => \N__43878\
        );

    \ppm_encoder_1.throttle_RNIVO123_0_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38016\,
            in2 => \N__38004\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37986\,
            in2 => \N__37974\,
            in3 => \N__37941\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37938\,
            in2 => \N__37932\,
            in3 => \N__37911\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37908\,
            in2 => \N__37902\,
            in3 => \N__37881\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37878\,
            in2 => \N__37869\,
            in3 => \N__37842\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37839\,
            in2 => \N__37832\,
            in3 => \N__37800\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37797\,
            in2 => \N__37788\,
            in3 => \N__37767\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38226\,
            in2 => \N__40247\,
            in3 => \N__38214\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38211\,
            in2 => \N__40622\,
            in3 => \N__38202\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38199\,
            in2 => \N__40575\,
            in3 => \N__38190\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38187\,
            in2 => \N__39029\,
            in3 => \N__38166\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38163\,
            in2 => \N__38151\,
            in3 => \N__38115\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38112\,
            in2 => \N__38100\,
            in3 => \N__38067\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38064\,
            in2 => \N__38052\,
            in3 => \N__38031\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41183\,
            in2 => \N__38028\,
            in3 => \N__38019\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42405\,
            in2 => \N__38451\,
            in3 => \N__38433\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38379\,
            in2 => \_gnd_net_\,
            in3 => \N__38430\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38427\,
            in2 => \_gnd_net_\,
            in3 => \N__38412\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38409\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__40644\,
            in1 => \N__41132\,
            in2 => \N__40992\,
            in3 => \N__38406\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40798\,
            in1 => \N__42273\,
            in2 => \_gnd_net_\,
            in3 => \N__41939\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38972\,
            in1 => \N__38372\,
            in2 => \_gnd_net_\,
            in3 => \N__38358\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_axb_0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38349\,
            in2 => \N__38334\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.un9_error_filt_add_1_axbZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_1_s_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38289\,
            in2 => \N__38274\,
            in3 => \N__38229\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_0\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_2_s_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38775\,
            in2 => \N__38760\,
            in3 => \N__38718\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_1\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_3_s_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38715\,
            in2 => \N__38700\,
            in3 => \N__38658\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_2\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_4_s_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39107\,
            in2 => \N__38655\,
            in3 => \N__38625\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_3\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_5_s_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38622\,
            in2 => \N__39124\,
            in3 => \N__38592\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_4\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_6_s_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39111\,
            in2 => \N__38589\,
            in3 => \N__38547\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_5\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_7_s_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38544\,
            in2 => \N__39125\,
            in3 => \N__38502\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_6\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_8_s_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39126\,
            in2 => \N__38499\,
            in3 => \N__38454\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_9_s_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39216\,
            in2 => \N__39132\,
            in3 => \N__39180\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_8\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_cry_10_s_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39130\,
            in2 => \N__39177\,
            in3 => \N__39135\,
            lcout => \pid_alt.un9_error_filt_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pid_alt.un9_error_filt_add_1_cry_9\,
            carryout => \pid_alt.un9_error_filt_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un9_error_filt_add_1_s_11_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39131\,
            in1 => \N__39081\,
            in2 => \_gnd_net_\,
            in3 => \N__39063\,
            lcout => \pid_alt.un9_error_filt_add_1_sZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40325\,
            lcout => \ppm_encoder_1.N_140_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41246\,
            in1 => \N__42289\,
            in2 => \_gnd_net_\,
            in3 => \N__41921\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__38947\,
            in1 => \N__40129\,
            in2 => \_gnd_net_\,
            in3 => \N__40425\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011111111"
        )
    port map (
            in0 => \N__39006\,
            in1 => \N__40990\,
            in2 => \N__41336\,
            in3 => \N__41147\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38948\,
            in1 => \N__38823\,
            in2 => \_gnd_net_\,
            in3 => \N__38808\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42610\,
            in2 => \N__38787\,
            in3 => \N__38784\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__42531\,
            sr => \N__43897\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42611\,
            in1 => \N__39447\,
            in2 => \_gnd_net_\,
            in3 => \N__40515\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__42531\,
            sr => \N__43897\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39432\,
            in1 => \N__42607\,
            in2 => \_gnd_net_\,
            in3 => \N__39417\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__42531\,
            sr => \N__43897\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42608\,
            in1 => \N__39411\,
            in2 => \_gnd_net_\,
            in3 => \N__39399\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__42531\,
            sr => \N__43897\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__39381\,
            in1 => \N__39363\,
            in2 => \N__39309\,
            in3 => \N__39354\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42609\,
            in1 => \N__39336\,
            in2 => \_gnd_net_\,
            in3 => \N__39321\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__42531\,
            sr => \N__43897\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__39300\,
            in1 => \N__39289\,
            in2 => \N__39273\,
            in3 => \N__39262\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__41289\,
            in1 => \N__39697\,
            in2 => \N__39228\,
            in3 => \N__39244\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_15_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__42369\,
            in1 => \N__39227\,
            in2 => \N__39746\,
            in3 => \N__41941\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47302\,
            ce => 'H',
            sr => \N__43900\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__39655\,
            in1 => \N__39755\,
            in2 => \N__39683\,
            in3 => \N__39780\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_17_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__41940\,
            in1 => \N__39742\,
            in2 => \N__39759\,
            in3 => \N__40754\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47302\,
            ce => 'H',
            sr => \N__43900\
        );

    \ppm_encoder_1.pulses2count_18_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__41651\,
            in1 => \N__39624\,
            in2 => \N__39747\,
            in3 => \N__41942\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47302\,
            ce => 'H',
            sr => \N__43900\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39698\,
            in1 => \N__39684\,
            in2 => \N__39660\,
            in3 => \N__39611\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39623\,
            in2 => \_gnd_net_\,
            in3 => \N__39610\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_0_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39594\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47279\,
            ce => \N__46798\,
            sr => \N__46585\
        );

    \pid_alt.error_i_reg_esr_3_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39561\,
            lcout => \pid_alt.error_i_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47279\,
            ce => \N__46798\,
            sr => \N__46585\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44485\,
            in2 => \_gnd_net_\,
            in3 => \N__44382\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_1_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__39494\,
            in1 => \N__39530\,
            in2 => \N__44495\,
            in3 => \N__44392\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47445\,
            ce => 'H',
            sr => \N__43856\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__40140\,
            in1 => \N__40491\,
            in2 => \_gnd_net_\,
            in3 => \N__39992\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39951\,
            in2 => \N__39942\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39930\,
            in2 => \_gnd_net_\,
            in3 => \N__39918\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39915\,
            in2 => \N__39906\,
            in3 => \N__39882\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39879\,
            in2 => \_gnd_net_\,
            in3 => \N__39855\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39852\,
            in2 => \_gnd_net_\,
            in3 => \N__39840\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39837\,
            in2 => \_gnd_net_\,
            in3 => \N__39825\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39822\,
            in2 => \N__39804\,
            in3 => \N__39783\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40722\,
            in3 => \N__40230\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40272\,
            in2 => \_gnd_net_\,
            in3 => \N__40227\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40584\,
            in2 => \_gnd_net_\,
            in3 => \N__40224\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41217\,
            in2 => \_gnd_net_\,
            in3 => \N__40215\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40212\,
            in2 => \_gnd_net_\,
            in3 => \N__40188\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40185\,
            in2 => \_gnd_net_\,
            in3 => \N__40167\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40164\,
            in2 => \N__40158\,
            in3 => \N__40146\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41172\,
            in2 => \_gnd_net_\,
            in3 => \N__40143\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42396\,
            in2 => \_gnd_net_\,
            in3 => \N__40503\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40782\,
            in3 => \N__40500\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41256\,
            in2 => \_gnd_net_\,
            in3 => \N__40497\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__42259\,
            in1 => \N__42023\,
            in2 => \N__41652\,
            in3 => \N__40494\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__40489\,
            in1 => \N__40421\,
            in2 => \N__40383\,
            in3 => \N__40326\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40275\,
            in3 => \N__44670\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__42022\,
            in1 => \N__40640\,
            in2 => \_gnd_net_\,
            in3 => \N__42258\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41599\,
            in1 => \N__40266\,
            in2 => \N__41473\,
            in3 => \N__40257\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47392\,
            ce => 'H',
            sr => \N__43888\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__40708\,
            in1 => \_gnd_net_\,
            in2 => \N__42040\,
            in3 => \N__42248\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__42247\,
            in1 => \N__42011\,
            in2 => \_gnd_net_\,
            in3 => \N__40709\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__40710\,
            in1 => \N__40978\,
            in2 => \N__41121\,
            in3 => \N__40695\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_8_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41600\,
            in1 => \N__40659\,
            in2 => \N__41474\,
            in3 => \N__40650\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47392\,
            ce => 'H',
            sr => \N__43888\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__40639\,
            in1 => \_gnd_net_\,
            in2 => \N__42041\,
            in3 => \N__42249\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__41610\,
            in1 => \N__40599\,
            in2 => \N__41496\,
            in3 => \N__40593\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47377\,
            ce => 'H',
            sr => \N__43893\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__42019\,
            in1 => \_gnd_net_\,
            in2 => \N__42284\,
            in3 => \N__40553\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40552\,
            in1 => \N__42254\,
            in2 => \_gnd_net_\,
            in3 => \N__42020\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__41094\,
            in1 => \N__40554\,
            in2 => \N__40542\,
            in3 => \N__40988\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__42021\,
            in1 => \_gnd_net_\,
            in2 => \N__42285\,
            in3 => \N__40741\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41242\,
            in1 => \N__42250\,
            in2 => \_gnd_net_\,
            in3 => \N__42018\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_14_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41612\,
            in1 => \N__41205\,
            in2 => \N__41497\,
            in3 => \N__41196\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47365\,
            ce => 'H',
            sr => \N__43895\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_14_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41158\,
            in1 => \N__42272\,
            in2 => \_gnd_net_\,
            in3 => \N__41938\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__41936\,
            in1 => \N__41159\,
            in2 => \_gnd_net_\,
            in3 => \N__42270\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__41160\,
            in1 => \N__41128\,
            in2 => \N__41025\,
            in3 => \N__40989\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_16_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41613\,
            in1 => \N__40824\,
            in2 => \N__41498\,
            in3 => \N__40815\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47365\,
            ce => 'H',
            sr => \N__43895\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__41937\,
            in1 => \N__40799\,
            in2 => \_gnd_net_\,
            in3 => \N__42271\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_17_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41614\,
            in1 => \N__40770\,
            in2 => \N__41499\,
            in3 => \N__40761\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47365\,
            ce => 'H',
            sr => \N__43895\
        );

    \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__42288\,
            in1 => \N__42361\,
            in2 => \N__42048\,
            in3 => \N__42346\,
            lcout => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__42362\,
            in1 => \N__42286\,
            in2 => \_gnd_net_\,
            in3 => \N__42042\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41608\,
            in1 => \N__42387\,
            in2 => \N__41501\,
            in3 => \N__42378\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__43896\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__42347\,
            in1 => \N__42287\,
            in2 => \N__41641\,
            in3 => \N__42043\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_18_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41609\,
            in1 => \N__41667\,
            in2 => \N__41502\,
            in3 => \N__41658\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__43896\
        );

    \ppm_encoder_1.init_pulses_13_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__41607\,
            in1 => \N__41514\,
            in2 => \N__41500\,
            in3 => \N__41346\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__43896\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42605\,
            in1 => \N__41307\,
            in2 => \_gnd_net_\,
            in3 => \N__41298\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__42539\,
            sr => \N__43898\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42604\,
            in1 => \N__41280\,
            in2 => \_gnd_net_\,
            in3 => \N__41268\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__42539\,
            sr => \N__43898\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42762\,
            in1 => \N__42606\,
            in2 => \_gnd_net_\,
            in3 => \N__42750\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__42539\,
            sr => \N__43898\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__42736\,
            in1 => \N__42660\,
            in2 => \N__42717\,
            in3 => \N__42707\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42616\,
            in1 => \N__42687\,
            in2 => \_gnd_net_\,
            in3 => \N__42672\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47322\,
            ce => \N__42538\,
            sr => \N__43901\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42612\,
            in1 => \N__42654\,
            in2 => \_gnd_net_\,
            in3 => \N__42642\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47322\,
            ce => \N__42538\,
            sr => \N__43901\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__42630\,
            in1 => \_gnd_net_\,
            in2 => \N__42618\,
            in3 => \N__42555\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47322\,
            ce => \N__42538\,
            sr => \N__43901\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__42489\,
            in1 => \N__42465\,
            in2 => \N__42459\,
            in3 => \N__42450\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42426\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43008\,
            in2 => \N__42417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43191\,
            in2 => \N__43068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42999\,
            in2 => \N__43179\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43167\,
            in2 => \N__43069\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43003\,
            in2 => \N__44565\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43161\,
            in2 => \N__43070\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43007\,
            in2 => \N__43155\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43146\,
            in2 => \N__43118\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43074\,
            in2 => \N__42771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44673\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44634\,
            in1 => \N__44625\,
            in2 => \N__44601\,
            in3 => \N__44589\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_0_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000101100"
        )
    port map (
            in0 => \N__44556\,
            in1 => \N__44378\,
            in2 => \N__44499\,
            in3 => \N__44469\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47465\,
            ce => 'H',
            sr => \N__43862\
        );

    \pid_alt.error_filt_prev_esr_21_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44343\,
            lcout => \pid_alt.error_filt_prevZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47453\,
            ce => \N__46819\,
            sr => \N__46600\
        );

    \Commands_frame_decoder.source_alt_ki_5_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44283\,
            in2 => \_gnd_net_\,
            in3 => \N__46675\,
            lcout => alt_ki_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47303\,
            ce => \N__44865\,
            sr => \_gnd_net_\
        );

    \GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_20_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44065\,
            lcout => \GB_BUFFER_reset_system_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_3_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43364\,
            in2 => \_gnd_net_\,
            in3 => \N__46680\,
            lcout => alt_ki_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47353\,
            ce => \N__44860\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_4_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43218\,
            lcout => \pid_alt.error_i_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47337\,
            ce => \N__46806\,
            sr => \N__46589\
        );

    \pid_alt.error_i_reg_esr_5_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45420\,
            lcout => \pid_alt.error_i_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47337\,
            ce => \N__46806\,
            sr => \N__46589\
        );

    \pid_alt.error_i_reg_esr_8_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45396\,
            lcout => \pid_alt.error_i_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47324\,
            ce => \N__46802\,
            sr => \N__46587\
        );

    \Commands_frame_decoder.source_alt_ki_4_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45366\,
            lcout => alt_ki_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47312\,
            ce => \N__44856\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_1_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45224\,
            in2 => \_gnd_net_\,
            in3 => \N__46676\,
            lcout => alt_ki_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47312\,
            ce => \N__44856\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_filt_prev_esr_19_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45066\,
            lcout => \pid_alt.error_filt_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47466\,
            ce => \N__46822\,
            sr => \N__46604\
        );

    \Commands_frame_decoder.source_alt_ki_7_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45013\,
            in2 => \_gnd_net_\,
            in3 => \N__46679\,
            lcout => alt_ki_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47338\,
            ce => \N__44864\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_10_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44772\,
            lcout => \pid_alt.error_i_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47325\,
            ce => \N__46803\,
            sr => \N__46588\
        );

    \pid_alt.error_i_reg_esr_11_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44739\,
            lcout => \pid_alt.error_i_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47339\,
            ce => \N__46807\,
            sr => \N__46590\
        );

    \pid_alt.error_i_reg_esr_12_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44706\,
            lcout => \pid_alt.error_i_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47339\,
            ce => \N__46807\,
            sr => \N__46590\
        );

    \pid_alt.error_i_reg_esr_13_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45831\,
            lcout => \pid_alt.error_i_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47339\,
            ce => \N__46807\,
            sr => \N__46590\
        );

    \pid_alt.error_filt_prev_esr_17_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45798\,
            lcout => \pid_alt.error_filt_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47473\,
            ce => \N__46824\,
            sr => \N__46611\
        );

    \pid_alt.error_filt_prev_esr_18_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45750\,
            lcout => \pid_alt.error_filt_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47473\,
            ce => \N__46824\,
            sr => \N__46611\
        );

    \pid_alt.error_filt_prev_esr_22_LC_24_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45702\,
            lcout => \pid_alt.error_filt_prevZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47473\,
            ce => \N__46824\,
            sr => \N__46611\
        );

    \pid_alt.error_filt_prev_esr_20_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45600\,
            lcout => \pid_alt.error_filt_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47471\,
            ce => \N__46823\,
            sr => \N__46607\
        );

    \pid_alt.error_filt_prev_esr_8_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45561\,
            lcout => \pid_alt.error_filt_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__46821\,
            sr => \N__46603\
        );

    \pid_alt.error_d_reg_esr_4_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45522\,
            lcout => \pid_alt.error_d_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__46820\,
            sr => \N__46601\
        );

    \pid_alt.error_filt_prev_esr_1_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45462\,
            lcout => \pid_alt.error_filt_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__46820\,
            sr => \N__46601\
        );

    \pid_alt.error_filt_prev_esr_2_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46176\,
            lcout => \pid_alt.error_filt_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__46820\,
            sr => \N__46601\
        );

    \pid_alt.error_filt_prev_esr_10_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46140\,
            lcout => \pid_alt.error_filt_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_11_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46104\,
            lcout => \pid_alt.error_filt_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_12_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46062\,
            lcout => \pid_alt.error_filt_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_13_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46023\,
            lcout => \pid_alt.error_filt_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_15_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45987\,
            lcout => \pid_alt.error_filt_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_16_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45942\,
            lcout => \pid_alt.error_filt_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__46818\,
            sr => \N__46599\
        );

    \pid_alt.error_filt_prev_esr_4_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45894\,
            lcout => \pid_alt.error_filt_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_5_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45864\,
            lcout => \pid_alt.error_filt_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_6_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46425\,
            lcout => \pid_alt.error_filt_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_7_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46392\,
            lcout => \pid_alt.error_filt_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_9_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46359\,
            lcout => \pid_alt.error_filt_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_3_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46314\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_filt_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__46817\,
            sr => \N__46597\
        );

    \pid_alt.error_filt_prev_esr_14_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46281\,
            lcout => \pid_alt.error_filt_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47429\,
            ce => \N__46816\,
            sr => \N__46596\
        );

    \pid_alt.error_i_reg_esr_7_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => \N__46813\,
            sr => \N__46595\
        );

    \pid_alt.error_i_reg_esr_6_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46224\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => \N__46813\,
            sr => \N__46595\
        );

    \pid_alt.error_i_reg_esr_15_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46203\,
            lcout => \pid_alt.error_i_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => \N__46811\,
            sr => \N__46594\
        );

    \pid_alt.error_i_reg_esr_9_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47625\,
            lcout => \pid_alt.error_i_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => \N__46811\,
            sr => \N__46594\
        );

    \pid_alt.error_i_reg_esr_14_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47604\,
            lcout => \pid_alt.error_i_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => \N__46811\,
            sr => \N__46594\
        );

    \pid_alt.error_i_reg_esr_20_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47586\,
            lcout => \pid_alt.error_i_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__46810\,
            sr => \N__46592\
        );

    \pid_alt.error_i_reg_esr_17_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47562\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__46810\,
            sr => \N__46592\
        );

    \pid_alt.error_i_reg_esr_18_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__46810\,
            sr => \N__46592\
        );

    \pid_alt.error_i_reg_esr_16_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47520\,
            lcout => \pid_alt.error_i_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__46810\,
            sr => \N__46592\
        );

    \pid_alt.error_i_reg_esr_19_LC_24_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47502\,
            lcout => \pid_alt.error_i_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => \N__46808\,
            sr => \N__46591\
        );
end \INTERFACE\;
