-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 16 2019 22:03:59

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_pc : in std_logic;
    debug_CH5_31B : out std_logic;
    debug_CH3_20A : out std_logic;
    debug_CH0_16A : out std_logic;
    uart_input_drone : in std_logic;
    ppm_output : out std_logic;
    debug_CH6_5B : out std_logic;
    debug_CH2_18A : out std_logic;
    debug_CH4_2A : out std_logic;
    debug_CH1_0A : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__52031\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51965\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51956\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51938\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51796\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51764\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51572\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51563\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51561\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51540\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51527\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51524\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51512\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51509\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51506\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51485\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51471\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51469\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51462\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51459\ : std_logic;
signal \N__51458\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51453\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51426\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51423\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51408\ : std_logic;
signal \N__51407\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51384\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51381\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51378\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51373\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51367\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51354\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51344\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51341\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51338\ : std_logic;
signal \N__51337\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51308\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50806\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50738\ : std_logic;
signal \N__50735\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50702\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50699\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50222\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50021\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49960\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49780\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49692\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49595\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49559\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49556\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49502\ : std_logic;
signal \N__49501\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41458\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40963\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40924\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pid_alt.O_1_12\ : std_logic;
signal \pid_alt.O_1_15\ : std_logic;
signal \pid_alt.O_1_16\ : std_logic;
signal \pid_alt.O_1_17\ : std_logic;
signal \pid_alt.O_1_19\ : std_logic;
signal \pid_alt.O_1_20\ : std_logic;
signal \pid_alt.O_1_7\ : std_logic;
signal \pid_alt.O_1_22\ : std_logic;
signal \pid_alt.O_1_23\ : std_logic;
signal \pid_alt.O_1_18\ : std_logic;
signal \pid_alt.O_1_24\ : std_logic;
signal \pid_alt.O_1_13\ : std_logic;
signal \pid_alt.O_1_14\ : std_logic;
signal \pid_alt.O_1_10\ : std_logic;
signal \pid_alt.O_1_21\ : std_logic;
signal \pid_alt.O_2_13\ : std_logic;
signal \pid_alt.O_2_21\ : std_logic;
signal \pid_alt.O_2_18\ : std_logic;
signal \pid_alt.O_2_20\ : std_logic;
signal \pid_alt.O_2_22\ : std_logic;
signal \pid_alt.O_2_11\ : std_logic;
signal \pid_alt.O_2_24\ : std_logic;
signal \pid_alt.O_2_7\ : std_logic;
signal \pid_alt.O_2_8\ : std_logic;
signal \pid_alt.O_2_23\ : std_logic;
signal \pid_alt.O_2_10\ : std_logic;
signal \pid_alt.O_2_9\ : std_logic;
signal \pid_alt.O_2_16\ : std_logic;
signal \pid_alt.O_2_17\ : std_logic;
signal \pid_alt.O_1_6\ : std_logic;
signal \pid_alt.O_2_12\ : std_logic;
signal \pid_alt.O_2_19\ : std_logic;
signal \pid_alt.O_2_14\ : std_logic;
signal \pid_alt.O_2_15\ : std_logic;
signal \pid_alt.O_1_5\ : std_logic;
signal \pid_side.O_0_9\ : std_logic;
signal \pid_side.O_0_19\ : std_logic;
signal \pid_side.O_0_14\ : std_logic;
signal \pid_side.O_0_8\ : std_logic;
signal \pid_side.O_0_10\ : std_logic;
signal \pid_side.O_0_23\ : std_logic;
signal \pid_side.O_0_15\ : std_logic;
signal \pid_side.O_0_18\ : std_logic;
signal \pid_side.O_0_11\ : std_logic;
signal \pid_side.O_0_6\ : std_logic;
signal \pid_side.O_0_17\ : std_logic;
signal \pid_side.O_0_16\ : std_logic;
signal \pid_side.O_0_12\ : std_logic;
signal \pid_side.O_0_20\ : std_logic;
signal \pid_side.O_0_21\ : std_logic;
signal \pid_side.O_0_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\ : std_logic;
signal \pid_alt.O_1_4\ : std_logic;
signal \pid_alt.O_3_4\ : std_logic;
signal \pid_alt.N_1505_i\ : std_logic;
signal \pid_alt.N_1505_i_cascade_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_axb_2_1\ : std_logic;
signal \pid_alt.N_1513_0_cascade_\ : std_logic;
signal \pid_alt.N_1505_i_0\ : std_logic;
signal \pid_alt.N_3_0\ : std_logic;
signal \pid_alt.N_1507_0\ : std_logic;
signal \pid_alt.N_5\ : std_logic;
signal \pid_alt.N_1511_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_0\ : std_logic;
signal \pid_alt.N_1505_i_1\ : std_logic;
signal \pid_alt.N_1507_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_1\ : std_logic;
signal \pid_alt.error_d_regZ0Z_1\ : std_logic;
signal \pid_alt.N_3_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\ : std_logic;
signal \pid_alt.error_d_regZ0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_2\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_3\ : std_logic;
signal \pid_alt.error_d_regZ0Z_3\ : std_logic;
signal \pid_alt.g0_4_0\ : std_logic;
signal \pid_alt.O_3_6\ : std_logic;
signal \pid_alt.error_p_regZ0Z_2\ : std_logic;
signal \pid_alt.O_3_7\ : std_logic;
signal \pid_alt.error_p_regZ0Z_3\ : std_logic;
signal \pid_alt.O_3_5\ : std_logic;
signal \pid_alt.error_p_regZ0Z_1\ : std_logic;
signal \pid_alt.O_3_12\ : std_logic;
signal \pid_alt.O_3_16\ : std_logic;
signal \pid_alt.O_3_17\ : std_logic;
signal \pid_alt.O_3_18\ : std_logic;
signal \pid_alt.O_3_24\ : std_logic;
signal \pid_alt.O_3_20\ : std_logic;
signal \pid_alt.O_3_21\ : std_logic;
signal \pid_alt.O_3_22\ : std_logic;
signal \pid_alt.O_3_23\ : std_logic;
signal \pid_alt.O_3_15\ : std_logic;
signal \pid_alt.O_3_19\ : std_logic;
signal \pid_alt.O_3_14\ : std_logic;
signal \pid_alt.O_3_8\ : std_logic;
signal \pid_alt.O_3_9\ : std_logic;
signal \pid_alt.O_3_10\ : std_logic;
signal \pid_alt.O_3_11\ : std_logic;
signal \pid_alt.O_3_13\ : std_logic;
signal \pid_alt.O_1_8\ : std_logic;
signal \pid_alt.O_1_11\ : std_logic;
signal alt_kd_6 : std_logic;
signal alt_kd_2 : std_logic;
signal alt_kd_7 : std_logic;
signal alt_kd_5 : std_logic;
signal alt_kd_1 : std_logic;
signal \pid_alt.O_1_9\ : std_logic;
signal alt_ki_0 : std_logic;
signal alt_ki_4 : std_logic;
signal alt_ki_1 : std_logic;
signal alt_ki_2 : std_logic;
signal alt_ki_3 : std_logic;
signal alt_ki_5 : std_logic;
signal \pid_alt.O_2_5\ : std_logic;
signal \pid_alt.O_2_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_4\ : std_logic;
signal \pid_alt.error_d_regZ0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_9\ : std_logic;
signal \pid_alt.error_p_regZ0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\ : std_logic;
signal \pid_alt.error_d_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_18\ : std_logic;
signal \pid_alt.error_p_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\ : std_logic;
signal \pid_alt.error_p_regZ0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_5\ : std_logic;
signal \pid_alt.error_d_regZ0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\ : std_logic;
signal \pid_alt.error_p_regZ0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_6\ : std_logic;
signal \pid_alt.error_d_regZ0Z_6\ : std_logic;
signal \pid_side.O_0_24\ : std_logic;
signal \pid_side.O_0_13\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_10\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_8\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_9\ : std_logic;
signal alt_kp_2 : std_logic;
signal alt_kp_3 : std_logic;
signal alt_kp_5 : std_logic;
signal alt_kp_6 : std_logic;
signal alt_kd_3 : std_logic;
signal alt_kd_0 : std_logic;
signal alt_kd_4 : std_logic;
signal \pid_alt.O_2_6\ : std_logic;
signal \pid_alt.N_850_0_g\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_6\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_10\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_8\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_1\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_0\ : std_logic;
signal \pid_alt.error_i_regZ0Z_2\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_1\ : std_logic;
signal \pid_alt.error_i_regZ0Z_3\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_2\ : std_logic;
signal \pid_alt.error_i_regZ0Z_4\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_3\ : std_logic;
signal \pid_alt.error_i_regZ0Z_5\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_4\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_6\ : std_logic;
signal \pid_alt.error_i_regZ0Z_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5\ : std_logic;
signal \pid_alt.error_i_regZ0Z_7\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_8\ : std_logic;
signal \pid_alt.error_i_regZ0Z_8\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_9\ : std_logic;
signal \pid_alt.error_i_regZ0Z_9\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_10\ : std_logic;
signal \pid_alt.error_i_regZ0Z_10\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9\ : std_logic;
signal \pid_alt.error_i_regZ0Z_11\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_10\ : std_logic;
signal \pid_alt.error_i_regZ0Z_12\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_11\ : std_logic;
signal \pid_alt.error_i_regZ0Z_13\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_12\ : std_logic;
signal \pid_alt.error_i_regZ0Z_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_13\ : std_logic;
signal \pid_alt.error_i_regZ0Z_15\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_15\ : std_logic;
signal \pid_alt.error_i_regZ0Z_16\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_16\ : std_logic;
signal \pid_alt.error_i_regZ0Z_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_17\ : std_logic;
signal \pid_alt.error_i_regZ0Z_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19\ : std_logic;
signal \pid_alt.error_i_regZ0Z_20\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\ : std_logic;
signal \pid_alt.error_p_regZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_17\ : std_logic;
signal \pid_alt.error_d_regZ0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\ : std_logic;
signal \pid_alt.error_d_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_16\ : std_logic;
signal \pid_alt.error_p_regZ0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_1_1_0\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \pid_alt.error_1\ : std_logic;
signal \pid_alt.error_cry_0\ : std_logic;
signal \pid_alt.error_2\ : std_logic;
signal \pid_alt.error_cry_1\ : std_logic;
signal \pid_alt.error_3\ : std_logic;
signal \pid_alt.error_cry_2\ : std_logic;
signal alt_command_0 : std_logic;
signal \pid_alt.error_4\ : std_logic;
signal \pid_alt.error_cry_3\ : std_logic;
signal drone_altitude_i_5 : std_logic;
signal alt_command_1 : std_logic;
signal \pid_alt.error_5\ : std_logic;
signal \pid_alt.error_cry_4\ : std_logic;
signal drone_altitude_i_6 : std_logic;
signal alt_command_2 : std_logic;
signal \pid_alt.error_6\ : std_logic;
signal \pid_alt.error_cry_5\ : std_logic;
signal drone_altitude_i_7 : std_logic;
signal alt_command_3 : std_logic;
signal \pid_alt.error_7\ : std_logic;
signal \pid_alt.error_cry_6\ : std_logic;
signal \pid_alt.error_cry_7\ : std_logic;
signal drone_altitude_i_8 : std_logic;
signal alt_command_4 : std_logic;
signal \pid_alt.error_8\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal drone_altitude_i_9 : std_logic;
signal alt_command_5 : std_logic;
signal \pid_alt.error_9\ : std_logic;
signal \pid_alt.error_cry_8\ : std_logic;
signal drone_altitude_i_10 : std_logic;
signal alt_command_6 : std_logic;
signal \pid_alt.error_10\ : std_logic;
signal \pid_alt.error_cry_9\ : std_logic;
signal alt_command_7 : std_logic;
signal \pid_alt.error_11\ : std_logic;
signal \pid_alt.error_cry_10\ : std_logic;
signal \pid_alt.error_12\ : std_logic;
signal \pid_alt.error_cry_11\ : std_logic;
signal \pid_alt.error_13\ : std_logic;
signal \pid_alt.error_cry_12\ : std_logic;
signal \pid_alt.error_14\ : std_logic;
signal \pid_alt.error_cry_13\ : std_logic;
signal drone_altitude_15 : std_logic;
signal \pid_alt.error_cry_14\ : std_logic;
signal \pid_alt.error_15\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_11\ : std_logic;
signal drone_altitude_i_11 : std_logic;
signal \pid_alt.error_i_acummZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_7\ : std_logic;
signal alt_kp_1 : std_logic;
signal alt_kp_7 : std_logic;
signal \Commands_frame_decoder.state_RNIRSI31Z0Z_11\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_3_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\ : std_logic;
signal \pid_alt.error_p_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_13\ : std_logic;
signal \pid_alt.error_d_regZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\ : std_logic;
signal \pid_alt.error_p_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_5\ : std_logic;
signal \pid_alt.N_295_cascade_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_1\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_3\ : std_logic;
signal \pid_alt.m39_i_a2_3\ : std_logic;
signal \pid_alt.m39_i_a2_4\ : std_logic;
signal \pid_alt.error_i_acumm7lto5\ : std_logic;
signal \pid_alt.N_294_cascade_\ : std_logic;
signal \pid_alt.N_294\ : std_logic;
signal \pid_alt.N_295\ : std_logic;
signal \pid_alt.error_i_acumm7lto4\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_4\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\ : std_logic;
signal \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_0\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_2\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_4\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_5\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_6\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_9\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_16\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_17\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_18\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_21\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_22\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_23\ : std_logic;
signal \pid_alt.error_axbZ0Z_13\ : std_logic;
signal drone_altitude_13 : std_logic;
signal \pid_alt.error_axbZ0Z_14\ : std_logic;
signal drone_altitude_14 : std_logic;
signal \pid_alt.error_axbZ0Z_2\ : std_logic;
signal \pid_alt.error_axbZ0Z_3\ : std_logic;
signal \pid_alt.error_d_reg_prev_i_0\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_8\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_9\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_10\ : std_logic;
signal \pid_alt.error_axbZ0Z_1\ : std_logic;
signal drone_altitude_12 : std_logic;
signal \pid_alt.error_axbZ0Z_12\ : std_logic;
signal \pid_side.error_axb_0\ : std_logic;
signal \bfn_4_21_0_\ : std_logic;
signal \pid_side.error_1\ : std_logic;
signal \pid_side.error_cry_0\ : std_logic;
signal \pid_side.error_2\ : std_logic;
signal \pid_side.error_cry_1\ : std_logic;
signal \pid_side.error_3\ : std_logic;
signal \pid_side.error_cry_2\ : std_logic;
signal \pid_side.error_4\ : std_logic;
signal \pid_side.error_cry_3\ : std_logic;
signal \pid_side.error_5\ : std_logic;
signal \pid_side.error_cry_0_0\ : std_logic;
signal \pid_side.error_6\ : std_logic;
signal \pid_side.error_cry_1_0\ : std_logic;
signal \pid_side.error_7\ : std_logic;
signal \pid_side.error_cry_2_0\ : std_logic;
signal \pid_side.error_cry_3_0\ : std_logic;
signal \drone_H_disp_side_i_8\ : std_logic;
signal \pid_side.error_8\ : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal \drone_H_disp_side_i_9\ : std_logic;
signal \pid_side.error_9\ : std_logic;
signal \pid_side.error_cry_4\ : std_logic;
signal \drone_H_disp_side_i_10\ : std_logic;
signal \pid_side.error_10\ : std_logic;
signal \pid_side.error_cry_5\ : std_logic;
signal \pid_side.error_11\ : std_logic;
signal \pid_side.error_cry_6\ : std_logic;
signal \pid_side.error_12\ : std_logic;
signal \pid_side.error_cry_7\ : std_logic;
signal \pid_side.error_13\ : std_logic;
signal \pid_side.error_cry_8\ : std_logic;
signal \pid_side.error_14\ : std_logic;
signal \pid_side.error_cry_9\ : std_logic;
signal \pid_side.error_cry_10\ : std_logic;
signal \pid_side.error_15\ : std_logic;
signal alt_kp_0 : std_logic;
signal \Commands_frame_decoder.N_418\ : std_logic;
signal \Commands_frame_decoder.N_382_2\ : std_logic;
signal \Commands_frame_decoder.N_383_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_0_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_11\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_0_2_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_3_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal \pid_alt.error_d_regZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_12\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\ : std_logic;
signal \pid_alt.error_p_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_10\ : std_logic;
signal \pid_alt.error_d_regZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\ : std_logic;
signal \pid_alt.error_d_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_11\ : std_logic;
signal \pid_alt.error_p_regZ0Z_11\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_11\ : std_logic;
signal \pid_alt.error_d_regZ0Z_0\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\ : std_logic;
signal \pid_alt.error_i_acumm7lto12\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_12\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_7\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_2\ : std_logic;
signal \pid_alt.un1_reset_1_i_a5_0_7_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_15\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_14\ : std_logic;
signal \pid_alt.un1_reset_1_i_a5_0_9\ : std_logic;
signal \pid_alt.un1_reset_1_i_a5_0_8\ : std_logic;
signal \pid_alt.N_557_cascade_\ : std_logic;
signal \pid_alt.un1_reset_1_i_a5_0_10\ : std_logic;
signal \pid_alt.N_304_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\ : std_logic;
signal \pid_alt.error_p_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_8\ : std_logic;
signal \pid_alt.error_d_regZ0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\ : std_logic;
signal \pid_alt.error_d_regZ0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_7\ : std_logic;
signal \pid_alt.error_p_regZ0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_20\ : std_logic;
signal \pid_alt.pid_preregZ0Z_19\ : std_logic;
signal \pid_alt.pid_preregZ0Z_22\ : std_logic;
signal \pid_alt.pid_preregZ0Z_17\ : std_logic;
signal \pid_alt.pid_preregZ0Z_21\ : std_logic;
signal \pid_alt.pid_preregZ0Z_15\ : std_logic;
signal \pid_alt.pid_preregZ0Z_23\ : std_logic;
signal \pid_alt.pid_preregZ0Z_18\ : std_logic;
signal \pid_alt.error_p_regZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\ : std_logic;
signal \pid_alt.error_d_regZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_19\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_20\ : std_logic;
signal \pid_alt.error_p_regZ0Z_20\ : std_logic;
signal \pid_alt.error_d_regZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_236_1_cascade_\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_236_1\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\ : std_logic;
signal drone_altitude_1 : std_logic;
signal drone_altitude_2 : std_logic;
signal drone_altitude_3 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_5\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_6\ : std_logic;
signal xy_kp_0 : std_logic;
signal xy_kp_2 : std_logic;
signal xy_kp_6 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_4\ : std_logic;
signal drone_altitude_i_4 : std_logic;
signal \pid_alt.error_i_regZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_0\ : std_logic;
signal \drone_H_disp_side_i_13\ : std_logic;
signal \drone_H_disp_side_i_6\ : std_logic;
signal side_command_0 : std_logic;
signal side_command_1 : std_logic;
signal side_command_2 : std_logic;
signal side_command_3 : std_logic;
signal side_command_4 : std_logic;
signal side_command_5 : std_logic;
signal side_command_6 : std_logic;
signal \drone_H_disp_side_15\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.WDT8lto13_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\ : std_logic;
signal \Commands_frame_decoder.preinitZ0\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0\ : std_logic;
signal \Commands_frame_decoder.N_377_0\ : std_logic;
signal \Commands_frame_decoder.N_377_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_384\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10lto13_1\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_3\ : std_logic;
signal \pid_alt.m7_e_4\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_19\ : std_logic;
signal \pid_alt.un1_reset_i_a5_1_10_7_cascade_\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_18\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_20\ : std_logic;
signal \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_16\ : std_logic;
signal \pid_alt.state_0_g_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_14\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_16\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_5\ : std_logic;
signal \dron_frame_decoder_1.N_755_0\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_7\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \drone_H_disp_side_i_4\ : std_logic;
signal \drone_H_disp_side_i_7\ : std_logic;
signal \drone_H_disp_side_i_5\ : std_logic;
signal \pid_side.error_axbZ0Z_2\ : std_logic;
signal \pid_side.error_axbZ0Z_3\ : std_logic;
signal alt_kp_4 : std_logic;
signal \Commands_frame_decoder.state_RNIF38SZ0Z_6\ : std_logic;
signal \pid_alt.state_RNIFCSD1Z0Z_0\ : std_logic;
signal \pid_alt.N_850_0\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_1__0__0_0\ : std_logic;
signal \Commands_frame_decoder.count_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \scaler_4.N_1684_i_l_ofxZ0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \Commands_frame_decoder.un1_state57_iZ0\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_8\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_11\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_12\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0\ : std_logic;
signal xy_kp_4 : std_logic;
signal \Commands_frame_decoder.stateZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_8\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_415\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_10\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_1\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_2\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_3\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_4\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_5\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_6\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_7\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_8\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_9\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_10\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_11\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_12\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_13\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_14\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_15\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_16\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_17\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_18\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_19\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_20\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \drone_H_disp_side_0\ : std_logic;
signal \drone_H_disp_side_2\ : std_logic;
signal \drone_H_disp_side_3\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_4\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_5\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_6\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_side_7\ : std_logic;
signal \dron_frame_decoder_1.N_747_0\ : std_logic;
signal alt_ki_7 : std_logic;
signal uart_input_pc_c : std_logic;
signal \uart_pc_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_1__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_3__0_Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_0\ : std_logic;
signal \debug_CH3_20A_c\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_422\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_AuxZ1Z_0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_412_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_14\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0\ : std_logic;
signal \dron_frame_decoder_1.N_177_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.N_412_4\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0\ : std_logic;
signal \dron_frame_decoder_1.N_175\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.N_431\ : std_logic;
signal \dron_frame_decoder_1.N_435\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_1\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_8_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.N_428\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_3\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_7_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_8\ : std_logic;
signal \pid_side.error_p_regZ0Z_11\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_10_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_3_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_4\ : std_logic;
signal \pid_side.error_p_regZ0Z_6\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_5_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_18_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_19\ : std_logic;
signal \pid_side.error_p_regZ0Z_15\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_14_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_14\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_13_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_16_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_17\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_19_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_20\ : std_logic;
signal \pid_side.error_p_regZ0Z_12\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_11_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_17_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_18\ : std_logic;
signal \pid_alt.error_d_reg_prevZ0Z_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_15\ : std_logic;
signal \pid_alt.error_d_regZ0Z_15\ : std_logic;
signal \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\ : std_logic;
signal \pid_side.error_axb_8_l_ofxZ0\ : std_logic;
signal side_command_7 : std_logic;
signal \pid_side.error_axbZ0Z_7\ : std_logic;
signal \drone_H_disp_front_2\ : std_logic;
signal \drone_H_disp_side_1\ : std_logic;
signal \pid_side.error_axbZ0Z_1\ : std_logic;
signal \pid_alt.state_1_0_0\ : std_logic;
signal \uart_pc.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_pc.N_143_cascade_\ : std_logic;
signal \uart_pc.data_rdyc_1\ : std_logic;
signal \uart_pc.data_rdyc_1_cascade_\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\ : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \scaler_4.debug_CH3_20A_c_0\ : std_logic;
signal \uart_pc.data_AuxZ1Z_2\ : std_logic;
signal \uart_pc.data_AuxZ1Z_1\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.data_rdyc_1_0\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_2\ : std_logic;
signal uart_drone_data_rdy : std_logic;
signal \pid_alt.pid_preregZ0Z_10\ : std_logic;
signal \pid_alt.un1_reset_i_a2_3_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_8\ : std_logic;
signal \pid_alt.un1_reset_i_a5_1_10_5_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_6\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_9_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_10\ : std_logic;
signal \pid_side.un1_reset_i_a2_3_cascade_\ : std_logic;
signal \pid_side.pid_preregZ0Z_18\ : std_logic;
signal \pid_side.pid_preregZ0Z_17\ : std_logic;
signal \pid_side.pid_preregZ0Z_19\ : std_logic;
signal \pid_side.pid_preregZ0Z_20\ : std_logic;
signal \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\ : std_logic;
signal \drone_H_disp_side_11\ : std_logic;
signal \drone_H_disp_side_13\ : std_logic;
signal \drone_H_disp_side_14\ : std_logic;
signal \dron_frame_decoder_1.N_739_0\ : std_logic;
signal \drone_H_disp_side_12\ : std_logic;
signal \drone_H_disp_side_i_12\ : std_logic;
signal \drone_H_disp_front_3\ : std_logic;
signal xy_kp_3 : std_logic;
signal \uart_drone_sync.aux_2__0__0_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.data_rdyc_1\ : std_logic;
signal \uart_drone_sync.aux_3__0__0_0\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa_cascade_\ : std_logic;
signal \uart_pc.N_145_cascade_\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \uart_pc.N_144_1_cascade_\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.N_152_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.CO0_cascade_\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \pid_alt.pid_preregZ0Z_9\ : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4\ : std_logic;
signal \pid_alt.un1_reset_i_a5_0_6_3\ : std_logic;
signal \pid_alt.N_306_5\ : std_logic;
signal \pid_alt.un1_reset_i_a5_0_6_2_cascade_\ : std_logic;
signal \pid_alt.un1_reset_i_a5_1_10_8\ : std_logic;
signal \pid_alt.un1_reset_i_a5_1_10_9\ : std_logic;
signal \pid_alt.un1_reset_i_a5_0_6_cascade_\ : std_logic;
signal \pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal \pid_alt.N_530\ : std_logic;
signal \pid_alt.N_535\ : std_logic;
signal \pid_alt.pid_preregZ0Z_5\ : std_logic;
signal \pid_alt.N_535_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_4\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_12\ : std_logic;
signal \pid_alt.pid_preregZ0Z_13\ : std_logic;
signal \pid_alt.pid_preregZ0Z_24\ : std_logic;
signal \pid_alt.N_551\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_6_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_7\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_2_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_16\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_15_THRU_CO\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_4_THRU_CO\ : std_logic;
signal \pid_side.error_p_regZ0Z_5\ : std_logic;
signal \pid_side.error_p_regZ0Z_13\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_12_THRU_CO\ : std_logic;
signal xy_kp_1 : std_logic;
signal xy_kp_7 : std_logic;
signal \pid_alt.stateZ0Z_0\ : std_logic;
signal \pid_alt.state_0_0\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \debug_CH0_16A_c\ : std_logic;
signal \uart_drone.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal scaler_4_data_6 : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal throttle_order_9 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal \pid_alt.N_72_i_1\ : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \pid_alt.pid_preregZ0Z_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_1\ : std_logic;
signal \pid_alt.pid_preregZ0Z_2\ : std_logic;
signal \pid_alt.pid_preregZ0Z_3\ : std_logic;
signal \pid_alt.N_472_1\ : std_logic;
signal \pid_alt.pid_preregZ0Z_11\ : std_logic;
signal \pid_alt.N_72_i\ : std_logic;
signal \pid_alt.N_299\ : std_logic;
signal \pid_alt.pid_preregZ0Z_7\ : std_logic;
signal \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\ : std_logic;
signal \ppm_encoder_1.N_292\ : std_logic;
signal \uart_drone.un1_state_7_0_cascade_\ : std_logic;
signal \uart_drone.N_152_cascade_\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal \pid_front.N_533_cascade_\ : std_logic;
signal \pid_front.N_10_1\ : std_logic;
signal \pid_front.un1_reset_i_a5_0_2_cascade_\ : std_logic;
signal \pid_front.un1_reset_i_a5_0_3\ : std_logic;
signal \pid_front.pid_preregZ0Z_1\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \uart_pc.state_srsts_i_0_2\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal scaler_4_data_11 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal throttle_order_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\ : std_logic;
signal throttle_order_2 : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal throttle_order_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal throttle_order_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\ : std_logic;
signal throttle_order_3 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\ : std_logic;
signal throttle_order_5 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\ : std_logic;
signal throttle_order_6 : std_logic;
signal \ppm_encoder_1.N_314_cascade_\ : std_logic;
signal \ppm_encoder_1.N_288_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_21\ : std_logic;
signal \pid_alt.N_557\ : std_logic;
signal \pid_alt.error_i_acumm7lto13\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_13\ : std_logic;
signal \pid_alt.N_72_i_0\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \ppm_encoder_1.N_291\ : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \uart_drone.N_145_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \debug_CH1_0A_c\ : std_logic;
signal \pid_side.state_ns_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_763_0\ : std_logic;
signal \pid_front.un1_reset_i_a5_0_5\ : std_logic;
signal \pid_front.un1_reset_i_1_cascade_\ : std_logic;
signal \pid_front.N_532\ : std_logic;
signal \pid_front.un1_reset_i_a2_3\ : std_logic;
signal \pid_front.stateZ0Z_1\ : std_logic;
signal \pid_front.N_287\ : std_logic;
signal \pid_front.N_533\ : std_logic;
signal \pid_front.state_0_1\ : std_logic;
signal \pid_front.pid_prereg_RNI2A6A6Z0Z_2\ : std_logic;
signal \pid_front.un1_reset_i_a5_1_6\ : std_logic;
signal \pid_front.N_315\ : std_logic;
signal \drone_H_disp_front_1\ : std_logic;
signal \pid_front.un1_reset_i_a5_1_5_cascade_\ : std_logic;
signal \pid_front.un1_reset_i_a5_1_8\ : std_logic;
signal \pid_front.pid_preregZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_8\ : std_logic;
signal \reset_module_System.reset6_15_cascade_\ : std_logic;
signal \reset_module_System.count_1_1\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_297_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.N_298_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal drone_altitude_0 : std_logic;
signal \pid_alt.drone_altitude_i_0\ : std_logic;
signal \pid_side.pid_preregZ0Z_10\ : std_logic;
signal side_order_11 : std_logic;
signal \pid_side.pid_preregZ0Z_6\ : std_logic;
signal \pid_side.pid_preregZ0Z_8\ : std_logic;
signal \pid_side.pid_preregZ0Z_9\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \pid_side.pid_preregZ0Z_11\ : std_logic;
signal \pid_side.pid_preregZ0Z_7\ : std_logic;
signal \pid_side.un1_reset_i_a5_1_5\ : std_logic;
signal \pid_side.pid_preregZ0Z_15\ : std_logic;
signal \pid_side.pid_preregZ0Z_14\ : std_logic;
signal \pid_side.m7_e_4\ : std_logic;
signal \pid_side.pid_preregZ0Z_16\ : std_logic;
signal \pid_side.un1_reset_i_a5_1_7\ : std_logic;
signal \pid_side.N_563_cascade_\ : std_logic;
signal \pid_side.un1_reset_i_a5_1_8\ : std_logic;
signal \pid_side.N_311_cascade_\ : std_logic;
signal \pid_side.un1_reset_i_a5_1_6\ : std_logic;
signal \pid_side.error_p_regZ0Z_2\ : std_logic;
signal \pid_side.un1_pid_prereg_cry_1_THRU_CO\ : std_logic;
signal \pid_side.un1_reset_i_a5_0_2\ : std_logic;
signal \pid_side.un1_reset_i_a5_0_3\ : std_logic;
signal \pid_front.N_569\ : std_logic;
signal \pid_front.pid_preregZ0Z_14\ : std_logic;
signal \pid_front.m7_e_4\ : std_logic;
signal \pid_front.pid_preregZ0Z_18\ : std_logic;
signal \pid_front.pid_preregZ0Z_19\ : std_logic;
signal \pid_front.pid_preregZ0Z_9\ : std_logic;
signal \pid_front.pid_preregZ0Z_11\ : std_logic;
signal \pid_front.pid_preregZ0Z_13\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.reset6_3_cascade_\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_313_cascade_\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.N_287\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\ : std_logic;
signal throttle_order_1 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.N_295\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10\ : std_logic;
signal \ppm_encoder_1.N_296\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal side_order_10 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal \pid_side.N_531\ : std_logic;
signal \pid_side.un1_reset_i_a5_0_5\ : std_logic;
signal \pid_side.un1_reset_i_1\ : std_logic;
signal side_order_1 : std_logic;
signal \pid_side.pid_preregZ0Z_2\ : std_logic;
signal side_order_2 : std_logic;
signal \pid_side.stateZ0Z_1\ : std_logic;
signal \pid_side.pid_preregZ0Z_3\ : std_logic;
signal \pid_side.N_291_cascade_\ : std_logic;
signal \pid_side.N_451_1\ : std_logic;
signal front_order_0 : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal front_order_1 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_1\ : std_logic;
signal front_order_3 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal front_order_9 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal front_order_11 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal front_order_12 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal \pid_front.pid_preregZ0Z_0\ : std_logic;
signal \pid_front.un1_reset_i_a5_1_7\ : std_logic;
signal uart_drone_data_7 : std_logic;
signal \pid_front.pid_preregZ0Z_17\ : std_logic;
signal \pid_front.pid_preregZ0Z_20\ : std_logic;
signal \pid_front.pid_preregZ0Z_7\ : std_logic;
signal \pid_front.pid_preregZ0Z_6\ : std_logic;
signal \pid_front.pid_preregZ0Z_12\ : std_logic;
signal \pid_front.pid_preregZ0Z_16\ : std_logic;
signal \pid_front.pid_preregZ0Z_2\ : std_logic;
signal \pid_front.pid_preregZ0Z_15\ : std_logic;
signal uart_drone_data_2 : std_logic;
signal uart_drone_data_3 : std_logic;
signal uart_drone_data_4 : std_logic;
signal uart_drone_data_5 : std_logic;
signal uart_drone_data_1 : std_logic;
signal scaler_4_data_4 : std_logic;
signal scaler_4_data_5 : std_logic;
signal \ppm_encoder_1.pid_altitude_dv_0\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8\ : std_logic;
signal \ppm_encoder_1.N_294_cascade_\ : std_logic;
signal side_order_8 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal front_order_8 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal throttle_order_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_1\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_m_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \pid_side.pid_preregZ0Z_12\ : std_logic;
signal side_order_12 : std_logic;
signal \pid_side.N_563\ : std_logic;
signal \pid_side.pid_preregZ0Z_21\ : std_logic;
signal \pid_side.pid_preregZ0Z_13\ : std_logic;
signal \pid_side.pid_preregZ0Z_4\ : std_logic;
signal \pid_side.N_534\ : std_logic;
signal \pid_side.N_291\ : std_logic;
signal \pid_side.pid_preregZ0Z_5\ : std_logic;
signal \pid_side.state_0_1\ : std_logic;
signal \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6\ : std_logic;
signal side_order_6 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\ : std_logic;
signal side_order_3 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\ : std_logic;
signal side_order_5 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal side_order_9 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal front_order_10 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal front_order_2 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\ : std_logic;
signal front_order_6 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal front_order_5 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal xy_kp_5 : std_logic;
signal \Commands_frame_decoder.state_RNIG48SZ0Z_7\ : std_logic;
signal \pid_front.pid_preregZ0Z_4\ : std_logic;
signal \pid_front.pid_preregZ0Z_5\ : std_logic;
signal \pid_front.pid_preregZ0Z_3\ : std_logic;
signal alt_ki_6 : std_logic;
signal \Commands_frame_decoder.state_RNIQRI31Z0Z_10\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_4\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_5\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_6\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_7\ : std_logic;
signal uart_pc_data_0 : std_logic;
signal uart_pc_data_1 : std_logic;
signal uart_pc_data_2 : std_logic;
signal uart_pc_data_3 : std_logic;
signal uart_pc_data_4 : std_logic;
signal uart_pc_data_5 : std_logic;
signal uart_pc_data_6 : std_logic;
signal uart_pc_data_7 : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_10\ : std_logic;
signal \dron_frame_decoder_1.drone_H_disp_front_9\ : std_logic;
signal front_command_7 : std_logic;
signal \drone_H_disp_front_11\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \debug_CH2_18A_c\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_6\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13\ : std_logic;
signal \ppm_encoder_1.N_299_cascade_\ : std_logic;
signal side_order_13 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal front_order_13 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal throttle_order_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.N_300_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\ : std_logic;
signal \pid_side.pid_preregZ0Z_0\ : std_logic;
signal \pid_side.state_0_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_53_d_cascade_\ : std_logic;
signal \ppm_encoder_1.N_134_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.N_221\ : std_logic;
signal \ppm_encoder_1.N_232_cascade_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.N_139\ : std_logic;
signal \ppm_encoder_1.N_232\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_3\ : std_logic;
signal \ppm_encoder_1.N_289\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_139_17\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal \pid_front.stateZ0Z_0\ : std_logic;
signal \pid_front.pid_preregZ0Z_8\ : std_logic;
signal uart_drone_data_0 : std_logic;
signal \dron_frame_decoder_1.N_731_0\ : std_logic;
signal \drone_H_disp_front_0\ : std_logic;
signal \pid_front.error_axb_0\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \pid_front.error_axbZ0Z_1\ : std_logic;
signal \pid_front.error_1\ : std_logic;
signal \pid_front.error_cry_0\ : std_logic;
signal \pid_front.error_axbZ0Z_2\ : std_logic;
signal \pid_front.error_2\ : std_logic;
signal \pid_front.error_cry_1\ : std_logic;
signal \pid_front.error_axbZ0Z_3\ : std_logic;
signal \pid_front.error_3\ : std_logic;
signal \pid_front.error_cry_2\ : std_logic;
signal front_command_0 : std_logic;
signal \drone_H_disp_front_i_4\ : std_logic;
signal \pid_front.error_4\ : std_logic;
signal \pid_front.error_cry_3\ : std_logic;
signal \drone_H_disp_front_i_5\ : std_logic;
signal front_command_1 : std_logic;
signal \pid_front.error_5\ : std_logic;
signal \pid_front.error_cry_0_0\ : std_logic;
signal \drone_H_disp_front_i_6\ : std_logic;
signal front_command_2 : std_logic;
signal \pid_front.error_6\ : std_logic;
signal \pid_front.error_cry_1_0\ : std_logic;
signal \drone_H_disp_front_i_7\ : std_logic;
signal front_command_3 : std_logic;
signal \pid_front.error_7\ : std_logic;
signal \pid_front.error_cry_2_0\ : std_logic;
signal \pid_front.error_cry_3_0\ : std_logic;
signal front_command_4 : std_logic;
signal \drone_H_disp_front_i_8\ : std_logic;
signal \pid_front.error_8\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \drone_H_disp_front_i_9\ : std_logic;
signal front_command_5 : std_logic;
signal \pid_front.error_9\ : std_logic;
signal \pid_front.error_cry_4\ : std_logic;
signal front_command_6 : std_logic;
signal \drone_H_disp_front_i_10\ : std_logic;
signal \pid_front.error_10\ : std_logic;
signal \pid_front.error_cry_5\ : std_logic;
signal \pid_front.error_axbZ0Z_7\ : std_logic;
signal \pid_front.error_11\ : std_logic;
signal \pid_front.error_cry_6\ : std_logic;
signal \pid_front.error_axb_8_l_ofx_0\ : std_logic;
signal \drone_H_disp_front_12\ : std_logic;
signal \pid_front.error_12\ : std_logic;
signal \pid_front.error_cry_7\ : std_logic;
signal \drone_H_disp_front_i_12\ : std_logic;
signal \drone_H_disp_front_13\ : std_logic;
signal \pid_front.error_13\ : std_logic;
signal \pid_front.error_cry_8\ : std_logic;
signal \drone_H_disp_front_i_13\ : std_logic;
signal \pid_front.error_14\ : std_logic;
signal \pid_front.error_cry_9\ : std_logic;
signal \drone_H_disp_front_15\ : std_logic;
signal \pid_front.error_cry_10\ : std_logic;
signal \pid_front.error_15\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal throttle_order_0 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_0\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.N_286_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_153_d\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_53_d\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal \ppm_encoder_1.N_1818_0\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7\ : std_logic;
signal \ppm_encoder_1.N_293_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal side_order_7 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal front_order_7 : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal throttle_order_7 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\ : std_logic;
signal side_order_4 : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\ : std_logic;
signal front_order_4 : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_290_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\ : std_logic;
signal throttle_order_4 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal pid_altitude_dv : std_logic;
signal side_order_0 : std_logic;
signal \ppm_encoder_1.aileronZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.N_1818_i\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.N_661_g\ : std_logic;
signal \bfn_18_22_0_\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_1_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_1\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_2_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_2\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_3_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_3\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_4_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_4\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_5_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_5\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_6_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_6\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_7_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_7\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_8\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_8_THRU_CO\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_9_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_9\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_10_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_10\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_11_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_11\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_12_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_12\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_13_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_13\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_14_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_14\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_15_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_15\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_16\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_16_THRU_CO\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_17_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_17\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_18_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_18\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_19_THRU_CO\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_19\ : std_logic;
signal \pid_front.un1_pid_prereg_cry_20\ : std_logic;
signal \pid_front.pid_preregZ0Z_21\ : std_logic;
signal \pid_front.state_0_0\ : std_logic;
signal uart_drone_data_6 : std_logic;
signal \drone_H_disp_front_14\ : std_logic;
signal \dron_frame_decoder_1.N_723_0\ : std_logic;
signal \GB_BUFFER_reset_system_g_THRU_CO\ : std_logic;
signal \pid_side.O_0_4\ : std_logic;
signal \pid_side.error_p_regZ0Z_0\ : std_logic;
signal \pid_side.O_0_5\ : std_logic;
signal \pid_side.state_RNINK4UZ0Z_1\ : std_logic;
signal \pid_side.O_0_7\ : std_logic;
signal \pid_side.error_p_regZ0Z_3\ : std_logic;
signal \pid_front.O_4\ : std_logic;
signal \pid_front.error_p_regZ0Z_0\ : std_logic;
signal \pid_side.stateZ0Z_0\ : std_logic;
signal \pid_side.error_p_regZ0Z_1\ : std_logic;
signal \pid_side.pid_preregZ0Z_1\ : std_logic;
signal reset_system_g : std_logic;
signal \pid_front.state_ns_0\ : std_logic;
signal reset_system : std_logic;
signal \pid_front.O_5\ : std_logic;
signal \pid_front.error_p_regZ0Z_1\ : std_logic;
signal \pid_front.O_13\ : std_logic;
signal \pid_front.error_p_regZ0Z_9\ : std_logic;
signal \pid_front.O_6\ : std_logic;
signal \pid_front.error_p_regZ0Z_2\ : std_logic;
signal \pid_front.O_9\ : std_logic;
signal \pid_front.error_p_regZ0Z_5\ : std_logic;
signal \pid_front.O_8\ : std_logic;
signal \pid_front.error_p_regZ0Z_4\ : std_logic;
signal \pid_front.O_18\ : std_logic;
signal \pid_front.error_p_regZ0Z_14\ : std_logic;
signal \pid_front.O_12\ : std_logic;
signal \pid_front.error_p_regZ0Z_8\ : std_logic;
signal \pid_front.O_14\ : std_logic;
signal \pid_front.error_p_regZ0Z_10\ : std_logic;
signal \pid_front.O_11\ : std_logic;
signal \pid_front.error_p_regZ0Z_7\ : std_logic;
signal \pid_front.O_7\ : std_logic;
signal \pid_front.error_p_regZ0Z_3\ : std_logic;
signal \pid_front.O_20\ : std_logic;
signal \pid_front.error_p_regZ0Z_16\ : std_logic;
signal \pid_front.O_10\ : std_logic;
signal \pid_front.error_p_regZ0Z_6\ : std_logic;
signal \pid_front.O_22\ : std_logic;
signal \pid_front.error_p_regZ0Z_18\ : std_logic;
signal \pid_front.O_23\ : std_logic;
signal \pid_front.error_p_regZ0Z_19\ : std_logic;
signal \pid_front.O_17\ : std_logic;
signal \pid_front.error_p_regZ0Z_13\ : std_logic;
signal \pid_front.O_19\ : std_logic;
signal \pid_front.error_p_regZ0Z_15\ : std_logic;
signal \pid_front.O_15\ : std_logic;
signal \pid_front.error_p_regZ0Z_11\ : std_logic;
signal \pid_front.O_16\ : std_logic;
signal \pid_front.error_p_regZ0Z_12\ : std_logic;
signal \pid_front.O_24\ : std_logic;
signal \pid_front.error_p_regZ0Z_20\ : std_logic;
signal \pid_front.state_RNIVIRQZ0Z_1\ : std_logic;
signal \pid_front.O_21\ : std_logic;
signal \pid_front.error_p_regZ0Z_17\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal \N_851_g\ : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_drone_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal \debug_CH2_18A_wire\ : std_logic;
signal \debug_CH0_16A_wire\ : std_logic;
signal \debug_CH1_0A_wire\ : std_logic;
signal \debug_CH5_31B_wire\ : std_logic;
signal \debug_CH4_2A_wire\ : std_logic;
signal ppm_output_wire : std_logic;
signal \debug_CH3_20A_wire\ : std_logic;
signal \debug_CH6_5B_wire\ : std_logic;
signal \pid_alt.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_front.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_side.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    clk_system_wire <= clk_system;
    uart_input_drone_wire <= uart_input_drone;
    uart_input_pc_wire <= uart_input_pc;
    debug_CH2_18A <= \debug_CH2_18A_wire\;
    debug_CH0_16A <= \debug_CH0_16A_wire\;
    debug_CH1_0A <= \debug_CH1_0A_wire\;
    debug_CH5_31B <= \debug_CH5_31B_wire\;
    debug_CH4_2A <= \debug_CH4_2A_wire\;
    ppm_output <= ppm_output_wire;
    debug_CH3_20A <= \debug_CH3_20A_wire\;
    debug_CH6_5B <= \debug_CH6_5B_wire\;
    \pid_alt.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_A_wire\ <= \N__22032\&\N__22089\&\N__21468\&\N__21520\&\N__21573\&\N__21630\&\N__21696\&\N__21759\&\N__21810\&\N__21873\&\N__21169\&\N__21225\&\N__21303\&\N__21342\&\N__21396\&\N__34334\;
    \pid_alt.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21944\&\N__20234\&\N__20246\&\N__25973\&\N__20261\&\N__20273\&\N__21956\&\N__23333\;
    \pid_alt.O_3_24\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_3_23\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_3_22\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_3_21\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_3_20\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_3_19\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_3_18\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_3_17\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_3_16\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_3_15\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_3_14\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_3_13\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_3_12\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_3_11\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_3_10\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_3_9\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_3_8\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_3_7\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_3_6\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_3_5\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_3_4\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__22033\&\N__22090\&\N__21475\&\N__21519\&\N__21574\&\N__21631\&\N__21697\&\N__21763\&\N__21811\&\N__21883\&\N__21165\&\N__21232\&\N__21304\&\N__21343\&\N__21397\&\N__34327\;
    \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27089\&\N__38870\&\N__19781\&\N__19697\&\N__19661\&\N__19673\&\N__19685\&\N__19709\;
    \pid_alt.O_2_24\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_2_23\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_2_22\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_2_21\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_2_20\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_2_19\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_2_18\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_2_17\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_2_16\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_2_15\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_2_14\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_2_13\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_2_12\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_2_11\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_2_10\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_2_9\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_2_8\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_2_7\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_2_6\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_2_5\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_2_4\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\ <= \N__22037\&\N__22097\&\N__21479\&\N__21527\&\N__21575\&\N__21635\&\N__21701\&\N__21767\&\N__21815\&\N__21884\&\N__21170\&\N__21239\&\N__21308\&\N__21350\&\N__21398\&\N__34326\;
    \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19583\&\N__19601\&\N__19745\&\N__20198\&\N__20222\&\N__19592\&\N__19733\&\N__20210\;
    \pid_alt.O_1_24\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_1_23\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_1_22\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_1_21\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_1_20\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_1_19\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_1_18\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_1_17\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_1_16\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_1_15\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_1_14\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_1_13\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_1_12\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_1_11\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_1_10\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_1_9\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_1_8\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_1_7\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_1_6\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_1_5\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_1_4\ <= \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\(4);
    \pid_front.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_mulonly_0_24_0_A_wire\ <= \N__43391\&\N__43424\&\N__43451\&\N__43499\&\N__43553\&\N__43577\&\N__43610\&\N__42875\&\N__42914\&\N__42947\&\N__42980\&\N__43013\&\N__43046\&\N__43076\&\N__42443\&\N__42482\;
    \pid_front.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_front.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30757\&\N__25076\&\N__39067\&\N__26756\&\N__29504\&\N__25112\&\N__30796\&\N__25142\;
    \pid_front.O_24\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_front.O_23\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_front.O_22\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_front.O_21\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_front.O_20\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_front.O_19\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_front.O_18\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_front.O_17\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_front.O_16\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_front.O_15\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_front.O_14\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_front.O_13\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_front.O_12\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_front.O_11\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_front.O_10\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_front.O_9\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_front.O_8\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_front.O_7\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_front.O_6\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_front.O_5\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_front.O_4\ <= \pid_front.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_side.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_mulonly_0_24_0_A_wire\ <= \N__23345\&\N__23366\&\N__23384\&\N__23402\&\N__23420\&\N__23438\&\N__23468\&\N__23495\&\N__23216\&\N__23234\&\N__23249\&\N__23264\&\N__23282\&\N__23297\&\N__23315\&\N__27158\;
    \pid_side.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_side.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__30758\&\N__25069\&\N__39071\&\N__26755\&\N__29503\&\N__25105\&\N__30797\&\N__25141\;
    \pid_side.O_0_24\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_side.O_0_23\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_side.O_0_22\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_side.O_0_21\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_side.O_0_20\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_side.O_0_19\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_side.O_0_18\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_side.O_0_17\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_side.O_0_16\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_side.O_0_15\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_side.O_0_14\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_side.O_0_13\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_side.O_0_12\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_side.O_0_11\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_side.O_0_10\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_side.O_0_9\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_side.O_0_8\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_side.O_0_7\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_side.O_0_6\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_side.O_0_5\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_side.O_0_4\ <= \pid_side.un2_error_mulonly_0_24_0_O_wire\(4);

    \pid_alt.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48236\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48235\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48206\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48199\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_2_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48230\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48229\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_2_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_2_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_2_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_2_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_2_mulonly_0_24_0_O_wire\
        );

    \pid_front.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48234\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48233\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_front.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_front.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_front.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_front.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_front.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_side.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__48193\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__48192\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_side.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_side.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_side.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_side.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_side.un2_error_mulonly_0_24_0_O_wire\
        );

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__52029\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52031\,
            DIN => \N__52030\,
            DOUT => \N__52029\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52031\,
            PADOUT => \N__52030\,
            PADIN => \N__52029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52020\,
            DIN => \N__52019\,
            DOUT => \N__52018\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52020\,
            PADOUT => \N__52019\,
            PADIN => \N__52018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52011\,
            DIN => \N__52010\,
            DOUT => \N__52009\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52011\,
            PADOUT => \N__52010\,
            PADIN => \N__52009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH2_18A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52002\,
            DIN => \N__52001\,
            DOUT => \N__52000\,
            PACKAGEPIN => \debug_CH2_18A_wire\
        );

    \debug_CH2_18A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52002\,
            PADOUT => \N__52001\,
            PADIN => \N__52000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__40706\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH0_16A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51993\,
            DIN => \N__51992\,
            DOUT => \N__51991\,
            PACKAGEPIN => \debug_CH0_16A_wire\
        );

    \debug_CH0_16A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51993\,
            PADOUT => \N__51992\,
            PADIN => \N__51991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH1_0A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51984\,
            DIN => \N__51983\,
            DOUT => \N__51982\,
            PACKAGEPIN => \debug_CH1_0A_wire\
        );

    \debug_CH1_0A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51984\,
            PADOUT => \N__51983\,
            PADIN => \N__51982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH5_31B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51975\,
            DIN => \N__51974\,
            DOUT => \N__51973\,
            PACKAGEPIN => \debug_CH5_31B_wire\
        );

    \debug_CH5_31B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51975\,
            PADOUT => \N__51974\,
            PADIN => \N__51973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH4_2A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51966\,
            DIN => \N__51965\,
            DOUT => \N__51964\,
            PACKAGEPIN => \debug_CH4_2A_wire\
        );

    \debug_CH4_2A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51966\,
            PADOUT => \N__51965\,
            PADIN => \N__51964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51957\,
            DIN => \N__51956\,
            DOUT => \N__51955\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51957\,
            PADOUT => \N__51956\,
            PADIN => \N__51955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32519\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH3_20A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51948\,
            DIN => \N__51947\,
            DOUT => \N__51946\,
            PACKAGEPIN => \debug_CH3_20A_wire\
        );

    \debug_CH3_20A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51948\,
            PADOUT => \N__51947\,
            PADIN => \N__51946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27203\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH6_5B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51939\,
            DIN => \N__51938\,
            DOUT => \N__51937\,
            PACKAGEPIN => \debug_CH6_5B_wire\
        );

    \debug_CH6_5B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__51939\,
            PADOUT => \N__51938\,
            PADIN => \N__51937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12609\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51917\
        );

    \I__12608\ : LocalMux
    port map (
            O => \N__51917\,
            I => \N__51914\
        );

    \I__12607\ : Odrv4
    port map (
            O => \N__51914\,
            I => \pid_front.O_23\
        );

    \I__12606\ : CascadeMux
    port map (
            O => \N__51911\,
            I => \N__51908\
        );

    \I__12605\ : InMux
    port map (
            O => \N__51908\,
            I => \N__51904\
        );

    \I__12604\ : InMux
    port map (
            O => \N__51907\,
            I => \N__51901\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__51904\,
            I => \N__51898\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__51901\,
            I => \N__51895\
        );

    \I__12601\ : Sp12to4
    port map (
            O => \N__51898\,
            I => \N__51892\
        );

    \I__12600\ : Span4Mux_h
    port map (
            O => \N__51895\,
            I => \N__51888\
        );

    \I__12599\ : Span12Mux_h
    port map (
            O => \N__51892\,
            I => \N__51885\
        );

    \I__12598\ : InMux
    port map (
            O => \N__51891\,
            I => \N__51882\
        );

    \I__12597\ : Span4Mux_h
    port map (
            O => \N__51888\,
            I => \N__51879\
        );

    \I__12596\ : Odrv12
    port map (
            O => \N__51885\,
            I => \pid_front.error_p_regZ0Z_19\
        );

    \I__12595\ : LocalMux
    port map (
            O => \N__51882\,
            I => \pid_front.error_p_regZ0Z_19\
        );

    \I__12594\ : Odrv4
    port map (
            O => \N__51879\,
            I => \pid_front.error_p_regZ0Z_19\
        );

    \I__12593\ : InMux
    port map (
            O => \N__51872\,
            I => \N__51869\
        );

    \I__12592\ : LocalMux
    port map (
            O => \N__51869\,
            I => \N__51866\
        );

    \I__12591\ : Odrv4
    port map (
            O => \N__51866\,
            I => \pid_front.O_17\
        );

    \I__12590\ : InMux
    port map (
            O => \N__51863\,
            I => \N__51860\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__51860\,
            I => \N__51857\
        );

    \I__12588\ : Span4Mux_h
    port map (
            O => \N__51857\,
            I => \N__51852\
        );

    \I__12587\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51849\
        );

    \I__12586\ : InMux
    port map (
            O => \N__51855\,
            I => \N__51846\
        );

    \I__12585\ : Sp12to4
    port map (
            O => \N__51852\,
            I => \N__51841\
        );

    \I__12584\ : LocalMux
    port map (
            O => \N__51849\,
            I => \N__51841\
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__51846\,
            I => \pid_front.error_p_regZ0Z_13\
        );

    \I__12582\ : Odrv12
    port map (
            O => \N__51841\,
            I => \pid_front.error_p_regZ0Z_13\
        );

    \I__12581\ : InMux
    port map (
            O => \N__51836\,
            I => \N__51833\
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__51833\,
            I => \N__51830\
        );

    \I__12579\ : Odrv4
    port map (
            O => \N__51830\,
            I => \pid_front.O_19\
        );

    \I__12578\ : InMux
    port map (
            O => \N__51827\,
            I => \N__51824\
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__51824\,
            I => \N__51819\
        );

    \I__12576\ : InMux
    port map (
            O => \N__51823\,
            I => \N__51816\
        );

    \I__12575\ : InMux
    port map (
            O => \N__51822\,
            I => \N__51813\
        );

    \I__12574\ : Sp12to4
    port map (
            O => \N__51819\,
            I => \N__51808\
        );

    \I__12573\ : LocalMux
    port map (
            O => \N__51816\,
            I => \N__51808\
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__51813\,
            I => \pid_front.error_p_regZ0Z_15\
        );

    \I__12571\ : Odrv12
    port map (
            O => \N__51808\,
            I => \pid_front.error_p_regZ0Z_15\
        );

    \I__12570\ : InMux
    port map (
            O => \N__51803\,
            I => \N__51800\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__51800\,
            I => \pid_front.O_15\
        );

    \I__12568\ : InMux
    port map (
            O => \N__51797\,
            I => \N__51792\
        );

    \I__12567\ : InMux
    port map (
            O => \N__51796\,
            I => \N__51789\
        );

    \I__12566\ : InMux
    port map (
            O => \N__51795\,
            I => \N__51786\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__51792\,
            I => \N__51781\
        );

    \I__12564\ : LocalMux
    port map (
            O => \N__51789\,
            I => \N__51781\
        );

    \I__12563\ : LocalMux
    port map (
            O => \N__51786\,
            I => \pid_front.error_p_regZ0Z_11\
        );

    \I__12562\ : Odrv12
    port map (
            O => \N__51781\,
            I => \pid_front.error_p_regZ0Z_11\
        );

    \I__12561\ : InMux
    port map (
            O => \N__51776\,
            I => \N__51773\
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__51773\,
            I => \N__51770\
        );

    \I__12559\ : Odrv4
    port map (
            O => \N__51770\,
            I => \pid_front.O_16\
        );

    \I__12558\ : InMux
    port map (
            O => \N__51767\,
            I => \N__51764\
        );

    \I__12557\ : LocalMux
    port map (
            O => \N__51764\,
            I => \N__51761\
        );

    \I__12556\ : Span4Mux_h
    port map (
            O => \N__51761\,
            I => \N__51757\
        );

    \I__12555\ : InMux
    port map (
            O => \N__51760\,
            I => \N__51754\
        );

    \I__12554\ : Span4Mux_h
    port map (
            O => \N__51757\,
            I => \N__51751\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__51754\,
            I => \N__51747\
        );

    \I__12552\ : Span4Mux_h
    port map (
            O => \N__51751\,
            I => \N__51744\
        );

    \I__12551\ : InMux
    port map (
            O => \N__51750\,
            I => \N__51741\
        );

    \I__12550\ : Span4Mux_h
    port map (
            O => \N__51747\,
            I => \N__51738\
        );

    \I__12549\ : Odrv4
    port map (
            O => \N__51744\,
            I => \pid_front.error_p_regZ0Z_12\
        );

    \I__12548\ : LocalMux
    port map (
            O => \N__51741\,
            I => \pid_front.error_p_regZ0Z_12\
        );

    \I__12547\ : Odrv4
    port map (
            O => \N__51738\,
            I => \pid_front.error_p_regZ0Z_12\
        );

    \I__12546\ : InMux
    port map (
            O => \N__51731\,
            I => \N__51728\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__51728\,
            I => \N__51725\
        );

    \I__12544\ : Odrv4
    port map (
            O => \N__51725\,
            I => \pid_front.O_24\
        );

    \I__12543\ : CascadeMux
    port map (
            O => \N__51722\,
            I => \N__51719\
        );

    \I__12542\ : InMux
    port map (
            O => \N__51719\,
            I => \N__51716\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__51716\,
            I => \N__51713\
        );

    \I__12540\ : Span4Mux_h
    port map (
            O => \N__51713\,
            I => \N__51708\
        );

    \I__12539\ : InMux
    port map (
            O => \N__51712\,
            I => \N__51703\
        );

    \I__12538\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51703\
        );

    \I__12537\ : Span4Mux_h
    port map (
            O => \N__51708\,
            I => \N__51700\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__51703\,
            I => \N__51696\
        );

    \I__12535\ : Span4Mux_h
    port map (
            O => \N__51700\,
            I => \N__51693\
        );

    \I__12534\ : InMux
    port map (
            O => \N__51699\,
            I => \N__51690\
        );

    \I__12533\ : Span4Mux_h
    port map (
            O => \N__51696\,
            I => \N__51687\
        );

    \I__12532\ : Odrv4
    port map (
            O => \N__51693\,
            I => \pid_front.error_p_regZ0Z_20\
        );

    \I__12531\ : LocalMux
    port map (
            O => \N__51690\,
            I => \pid_front.error_p_regZ0Z_20\
        );

    \I__12530\ : Odrv4
    port map (
            O => \N__51687\,
            I => \pid_front.error_p_regZ0Z_20\
        );

    \I__12529\ : CascadeMux
    port map (
            O => \N__51680\,
            I => \N__51672\
        );

    \I__12528\ : InMux
    port map (
            O => \N__51679\,
            I => \N__51652\
        );

    \I__12527\ : InMux
    port map (
            O => \N__51678\,
            I => \N__51652\
        );

    \I__12526\ : InMux
    port map (
            O => \N__51677\,
            I => \N__51645\
        );

    \I__12525\ : InMux
    port map (
            O => \N__51676\,
            I => \N__51645\
        );

    \I__12524\ : InMux
    port map (
            O => \N__51675\,
            I => \N__51645\
        );

    \I__12523\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51640\
        );

    \I__12522\ : InMux
    port map (
            O => \N__51671\,
            I => \N__51640\
        );

    \I__12521\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51629\
        );

    \I__12520\ : InMux
    port map (
            O => \N__51669\,
            I => \N__51629\
        );

    \I__12519\ : InMux
    port map (
            O => \N__51668\,
            I => \N__51629\
        );

    \I__12518\ : InMux
    port map (
            O => \N__51667\,
            I => \N__51629\
        );

    \I__12517\ : InMux
    port map (
            O => \N__51666\,
            I => \N__51629\
        );

    \I__12516\ : InMux
    port map (
            O => \N__51665\,
            I => \N__51618\
        );

    \I__12515\ : InMux
    port map (
            O => \N__51664\,
            I => \N__51618\
        );

    \I__12514\ : InMux
    port map (
            O => \N__51663\,
            I => \N__51618\
        );

    \I__12513\ : InMux
    port map (
            O => \N__51662\,
            I => \N__51618\
        );

    \I__12512\ : InMux
    port map (
            O => \N__51661\,
            I => \N__51618\
        );

    \I__12511\ : InMux
    port map (
            O => \N__51660\,
            I => \N__51613\
        );

    \I__12510\ : InMux
    port map (
            O => \N__51659\,
            I => \N__51613\
        );

    \I__12509\ : InMux
    port map (
            O => \N__51658\,
            I => \N__51610\
        );

    \I__12508\ : InMux
    port map (
            O => \N__51657\,
            I => \N__51607\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__51652\,
            I => \N__51602\
        );

    \I__12506\ : LocalMux
    port map (
            O => \N__51645\,
            I => \N__51602\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__51640\,
            I => \N__51595\
        );

    \I__12504\ : LocalMux
    port map (
            O => \N__51629\,
            I => \N__51595\
        );

    \I__12503\ : LocalMux
    port map (
            O => \N__51618\,
            I => \N__51595\
        );

    \I__12502\ : LocalMux
    port map (
            O => \N__51613\,
            I => \N__51592\
        );

    \I__12501\ : LocalMux
    port map (
            O => \N__51610\,
            I => \N__51587\
        );

    \I__12500\ : LocalMux
    port map (
            O => \N__51607\,
            I => \N__51587\
        );

    \I__12499\ : Span4Mux_v
    port map (
            O => \N__51602\,
            I => \N__51582\
        );

    \I__12498\ : Span4Mux_v
    port map (
            O => \N__51595\,
            I => \N__51582\
        );

    \I__12497\ : Odrv4
    port map (
            O => \N__51592\,
            I => \pid_front.state_RNIVIRQZ0Z_1\
        );

    \I__12496\ : Odrv4
    port map (
            O => \N__51587\,
            I => \pid_front.state_RNIVIRQZ0Z_1\
        );

    \I__12495\ : Odrv4
    port map (
            O => \N__51582\,
            I => \pid_front.state_RNIVIRQZ0Z_1\
        );

    \I__12494\ : InMux
    port map (
            O => \N__51575\,
            I => \N__51572\
        );

    \I__12493\ : LocalMux
    port map (
            O => \N__51572\,
            I => \pid_front.O_21\
        );

    \I__12492\ : InMux
    port map (
            O => \N__51569\,
            I => \N__51566\
        );

    \I__12491\ : LocalMux
    port map (
            O => \N__51566\,
            I => \N__51563\
        );

    \I__12490\ : Span4Mux_v
    port map (
            O => \N__51563\,
            I => \N__51558\
        );

    \I__12489\ : InMux
    port map (
            O => \N__51562\,
            I => \N__51555\
        );

    \I__12488\ : InMux
    port map (
            O => \N__51561\,
            I => \N__51552\
        );

    \I__12487\ : Sp12to4
    port map (
            O => \N__51558\,
            I => \N__51547\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__51555\,
            I => \N__51547\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__51552\,
            I => \pid_front.error_p_regZ0Z_17\
        );

    \I__12484\ : Odrv12
    port map (
            O => \N__51547\,
            I => \pid_front.error_p_regZ0Z_17\
        );

    \I__12483\ : ClkMux
    port map (
            O => \N__51542\,
            I => \N__50831\
        );

    \I__12482\ : ClkMux
    port map (
            O => \N__51541\,
            I => \N__50831\
        );

    \I__12481\ : ClkMux
    port map (
            O => \N__51540\,
            I => \N__50831\
        );

    \I__12480\ : ClkMux
    port map (
            O => \N__51539\,
            I => \N__50831\
        );

    \I__12479\ : ClkMux
    port map (
            O => \N__51538\,
            I => \N__50831\
        );

    \I__12478\ : ClkMux
    port map (
            O => \N__51537\,
            I => \N__50831\
        );

    \I__12477\ : ClkMux
    port map (
            O => \N__51536\,
            I => \N__50831\
        );

    \I__12476\ : ClkMux
    port map (
            O => \N__51535\,
            I => \N__50831\
        );

    \I__12475\ : ClkMux
    port map (
            O => \N__51534\,
            I => \N__50831\
        );

    \I__12474\ : ClkMux
    port map (
            O => \N__51533\,
            I => \N__50831\
        );

    \I__12473\ : ClkMux
    port map (
            O => \N__51532\,
            I => \N__50831\
        );

    \I__12472\ : ClkMux
    port map (
            O => \N__51531\,
            I => \N__50831\
        );

    \I__12471\ : ClkMux
    port map (
            O => \N__51530\,
            I => \N__50831\
        );

    \I__12470\ : ClkMux
    port map (
            O => \N__51529\,
            I => \N__50831\
        );

    \I__12469\ : ClkMux
    port map (
            O => \N__51528\,
            I => \N__50831\
        );

    \I__12468\ : ClkMux
    port map (
            O => \N__51527\,
            I => \N__50831\
        );

    \I__12467\ : ClkMux
    port map (
            O => \N__51526\,
            I => \N__50831\
        );

    \I__12466\ : ClkMux
    port map (
            O => \N__51525\,
            I => \N__50831\
        );

    \I__12465\ : ClkMux
    port map (
            O => \N__51524\,
            I => \N__50831\
        );

    \I__12464\ : ClkMux
    port map (
            O => \N__51523\,
            I => \N__50831\
        );

    \I__12463\ : ClkMux
    port map (
            O => \N__51522\,
            I => \N__50831\
        );

    \I__12462\ : ClkMux
    port map (
            O => \N__51521\,
            I => \N__50831\
        );

    \I__12461\ : ClkMux
    port map (
            O => \N__51520\,
            I => \N__50831\
        );

    \I__12460\ : ClkMux
    port map (
            O => \N__51519\,
            I => \N__50831\
        );

    \I__12459\ : ClkMux
    port map (
            O => \N__51518\,
            I => \N__50831\
        );

    \I__12458\ : ClkMux
    port map (
            O => \N__51517\,
            I => \N__50831\
        );

    \I__12457\ : ClkMux
    port map (
            O => \N__51516\,
            I => \N__50831\
        );

    \I__12456\ : ClkMux
    port map (
            O => \N__51515\,
            I => \N__50831\
        );

    \I__12455\ : ClkMux
    port map (
            O => \N__51514\,
            I => \N__50831\
        );

    \I__12454\ : ClkMux
    port map (
            O => \N__51513\,
            I => \N__50831\
        );

    \I__12453\ : ClkMux
    port map (
            O => \N__51512\,
            I => \N__50831\
        );

    \I__12452\ : ClkMux
    port map (
            O => \N__51511\,
            I => \N__50831\
        );

    \I__12451\ : ClkMux
    port map (
            O => \N__51510\,
            I => \N__50831\
        );

    \I__12450\ : ClkMux
    port map (
            O => \N__51509\,
            I => \N__50831\
        );

    \I__12449\ : ClkMux
    port map (
            O => \N__51508\,
            I => \N__50831\
        );

    \I__12448\ : ClkMux
    port map (
            O => \N__51507\,
            I => \N__50831\
        );

    \I__12447\ : ClkMux
    port map (
            O => \N__51506\,
            I => \N__50831\
        );

    \I__12446\ : ClkMux
    port map (
            O => \N__51505\,
            I => \N__50831\
        );

    \I__12445\ : ClkMux
    port map (
            O => \N__51504\,
            I => \N__50831\
        );

    \I__12444\ : ClkMux
    port map (
            O => \N__51503\,
            I => \N__50831\
        );

    \I__12443\ : ClkMux
    port map (
            O => \N__51502\,
            I => \N__50831\
        );

    \I__12442\ : ClkMux
    port map (
            O => \N__51501\,
            I => \N__50831\
        );

    \I__12441\ : ClkMux
    port map (
            O => \N__51500\,
            I => \N__50831\
        );

    \I__12440\ : ClkMux
    port map (
            O => \N__51499\,
            I => \N__50831\
        );

    \I__12439\ : ClkMux
    port map (
            O => \N__51498\,
            I => \N__50831\
        );

    \I__12438\ : ClkMux
    port map (
            O => \N__51497\,
            I => \N__50831\
        );

    \I__12437\ : ClkMux
    port map (
            O => \N__51496\,
            I => \N__50831\
        );

    \I__12436\ : ClkMux
    port map (
            O => \N__51495\,
            I => \N__50831\
        );

    \I__12435\ : ClkMux
    port map (
            O => \N__51494\,
            I => \N__50831\
        );

    \I__12434\ : ClkMux
    port map (
            O => \N__51493\,
            I => \N__50831\
        );

    \I__12433\ : ClkMux
    port map (
            O => \N__51492\,
            I => \N__50831\
        );

    \I__12432\ : ClkMux
    port map (
            O => \N__51491\,
            I => \N__50831\
        );

    \I__12431\ : ClkMux
    port map (
            O => \N__51490\,
            I => \N__50831\
        );

    \I__12430\ : ClkMux
    port map (
            O => \N__51489\,
            I => \N__50831\
        );

    \I__12429\ : ClkMux
    port map (
            O => \N__51488\,
            I => \N__50831\
        );

    \I__12428\ : ClkMux
    port map (
            O => \N__51487\,
            I => \N__50831\
        );

    \I__12427\ : ClkMux
    port map (
            O => \N__51486\,
            I => \N__50831\
        );

    \I__12426\ : ClkMux
    port map (
            O => \N__51485\,
            I => \N__50831\
        );

    \I__12425\ : ClkMux
    port map (
            O => \N__51484\,
            I => \N__50831\
        );

    \I__12424\ : ClkMux
    port map (
            O => \N__51483\,
            I => \N__50831\
        );

    \I__12423\ : ClkMux
    port map (
            O => \N__51482\,
            I => \N__50831\
        );

    \I__12422\ : ClkMux
    port map (
            O => \N__51481\,
            I => \N__50831\
        );

    \I__12421\ : ClkMux
    port map (
            O => \N__51480\,
            I => \N__50831\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__51479\,
            I => \N__50831\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__51478\,
            I => \N__50831\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__51477\,
            I => \N__50831\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__51476\,
            I => \N__50831\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__51475\,
            I => \N__50831\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__51474\,
            I => \N__50831\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__51473\,
            I => \N__50831\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__51472\,
            I => \N__50831\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__51471\,
            I => \N__50831\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__51470\,
            I => \N__50831\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__51469\,
            I => \N__50831\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__51468\,
            I => \N__50831\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__51467\,
            I => \N__50831\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__51466\,
            I => \N__50831\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__51465\,
            I => \N__50831\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__51464\,
            I => \N__50831\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__51463\,
            I => \N__50831\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__51462\,
            I => \N__50831\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__51461\,
            I => \N__50831\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__51460\,
            I => \N__50831\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__51459\,
            I => \N__50831\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__51458\,
            I => \N__50831\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__51457\,
            I => \N__50831\
        );

    \I__12397\ : ClkMux
    port map (
            O => \N__51456\,
            I => \N__50831\
        );

    \I__12396\ : ClkMux
    port map (
            O => \N__51455\,
            I => \N__50831\
        );

    \I__12395\ : ClkMux
    port map (
            O => \N__51454\,
            I => \N__50831\
        );

    \I__12394\ : ClkMux
    port map (
            O => \N__51453\,
            I => \N__50831\
        );

    \I__12393\ : ClkMux
    port map (
            O => \N__51452\,
            I => \N__50831\
        );

    \I__12392\ : ClkMux
    port map (
            O => \N__51451\,
            I => \N__50831\
        );

    \I__12391\ : ClkMux
    port map (
            O => \N__51450\,
            I => \N__50831\
        );

    \I__12390\ : ClkMux
    port map (
            O => \N__51449\,
            I => \N__50831\
        );

    \I__12389\ : ClkMux
    port map (
            O => \N__51448\,
            I => \N__50831\
        );

    \I__12388\ : ClkMux
    port map (
            O => \N__51447\,
            I => \N__50831\
        );

    \I__12387\ : ClkMux
    port map (
            O => \N__51446\,
            I => \N__50831\
        );

    \I__12386\ : ClkMux
    port map (
            O => \N__51445\,
            I => \N__50831\
        );

    \I__12385\ : ClkMux
    port map (
            O => \N__51444\,
            I => \N__50831\
        );

    \I__12384\ : ClkMux
    port map (
            O => \N__51443\,
            I => \N__50831\
        );

    \I__12383\ : ClkMux
    port map (
            O => \N__51442\,
            I => \N__50831\
        );

    \I__12382\ : ClkMux
    port map (
            O => \N__51441\,
            I => \N__50831\
        );

    \I__12381\ : ClkMux
    port map (
            O => \N__51440\,
            I => \N__50831\
        );

    \I__12380\ : ClkMux
    port map (
            O => \N__51439\,
            I => \N__50831\
        );

    \I__12379\ : ClkMux
    port map (
            O => \N__51438\,
            I => \N__50831\
        );

    \I__12378\ : ClkMux
    port map (
            O => \N__51437\,
            I => \N__50831\
        );

    \I__12377\ : ClkMux
    port map (
            O => \N__51436\,
            I => \N__50831\
        );

    \I__12376\ : ClkMux
    port map (
            O => \N__51435\,
            I => \N__50831\
        );

    \I__12375\ : ClkMux
    port map (
            O => \N__51434\,
            I => \N__50831\
        );

    \I__12374\ : ClkMux
    port map (
            O => \N__51433\,
            I => \N__50831\
        );

    \I__12373\ : ClkMux
    port map (
            O => \N__51432\,
            I => \N__50831\
        );

    \I__12372\ : ClkMux
    port map (
            O => \N__51431\,
            I => \N__50831\
        );

    \I__12371\ : ClkMux
    port map (
            O => \N__51430\,
            I => \N__50831\
        );

    \I__12370\ : ClkMux
    port map (
            O => \N__51429\,
            I => \N__50831\
        );

    \I__12369\ : ClkMux
    port map (
            O => \N__51428\,
            I => \N__50831\
        );

    \I__12368\ : ClkMux
    port map (
            O => \N__51427\,
            I => \N__50831\
        );

    \I__12367\ : ClkMux
    port map (
            O => \N__51426\,
            I => \N__50831\
        );

    \I__12366\ : ClkMux
    port map (
            O => \N__51425\,
            I => \N__50831\
        );

    \I__12365\ : ClkMux
    port map (
            O => \N__51424\,
            I => \N__50831\
        );

    \I__12364\ : ClkMux
    port map (
            O => \N__51423\,
            I => \N__50831\
        );

    \I__12363\ : ClkMux
    port map (
            O => \N__51422\,
            I => \N__50831\
        );

    \I__12362\ : ClkMux
    port map (
            O => \N__51421\,
            I => \N__50831\
        );

    \I__12361\ : ClkMux
    port map (
            O => \N__51420\,
            I => \N__50831\
        );

    \I__12360\ : ClkMux
    port map (
            O => \N__51419\,
            I => \N__50831\
        );

    \I__12359\ : ClkMux
    port map (
            O => \N__51418\,
            I => \N__50831\
        );

    \I__12358\ : ClkMux
    port map (
            O => \N__51417\,
            I => \N__50831\
        );

    \I__12357\ : ClkMux
    port map (
            O => \N__51416\,
            I => \N__50831\
        );

    \I__12356\ : ClkMux
    port map (
            O => \N__51415\,
            I => \N__50831\
        );

    \I__12355\ : ClkMux
    port map (
            O => \N__51414\,
            I => \N__50831\
        );

    \I__12354\ : ClkMux
    port map (
            O => \N__51413\,
            I => \N__50831\
        );

    \I__12353\ : ClkMux
    port map (
            O => \N__51412\,
            I => \N__50831\
        );

    \I__12352\ : ClkMux
    port map (
            O => \N__51411\,
            I => \N__50831\
        );

    \I__12351\ : ClkMux
    port map (
            O => \N__51410\,
            I => \N__50831\
        );

    \I__12350\ : ClkMux
    port map (
            O => \N__51409\,
            I => \N__50831\
        );

    \I__12349\ : ClkMux
    port map (
            O => \N__51408\,
            I => \N__50831\
        );

    \I__12348\ : ClkMux
    port map (
            O => \N__51407\,
            I => \N__50831\
        );

    \I__12347\ : ClkMux
    port map (
            O => \N__51406\,
            I => \N__50831\
        );

    \I__12346\ : ClkMux
    port map (
            O => \N__51405\,
            I => \N__50831\
        );

    \I__12345\ : ClkMux
    port map (
            O => \N__51404\,
            I => \N__50831\
        );

    \I__12344\ : ClkMux
    port map (
            O => \N__51403\,
            I => \N__50831\
        );

    \I__12343\ : ClkMux
    port map (
            O => \N__51402\,
            I => \N__50831\
        );

    \I__12342\ : ClkMux
    port map (
            O => \N__51401\,
            I => \N__50831\
        );

    \I__12341\ : ClkMux
    port map (
            O => \N__51400\,
            I => \N__50831\
        );

    \I__12340\ : ClkMux
    port map (
            O => \N__51399\,
            I => \N__50831\
        );

    \I__12339\ : ClkMux
    port map (
            O => \N__51398\,
            I => \N__50831\
        );

    \I__12338\ : ClkMux
    port map (
            O => \N__51397\,
            I => \N__50831\
        );

    \I__12337\ : ClkMux
    port map (
            O => \N__51396\,
            I => \N__50831\
        );

    \I__12336\ : ClkMux
    port map (
            O => \N__51395\,
            I => \N__50831\
        );

    \I__12335\ : ClkMux
    port map (
            O => \N__51394\,
            I => \N__50831\
        );

    \I__12334\ : ClkMux
    port map (
            O => \N__51393\,
            I => \N__50831\
        );

    \I__12333\ : ClkMux
    port map (
            O => \N__51392\,
            I => \N__50831\
        );

    \I__12332\ : ClkMux
    port map (
            O => \N__51391\,
            I => \N__50831\
        );

    \I__12331\ : ClkMux
    port map (
            O => \N__51390\,
            I => \N__50831\
        );

    \I__12330\ : ClkMux
    port map (
            O => \N__51389\,
            I => \N__50831\
        );

    \I__12329\ : ClkMux
    port map (
            O => \N__51388\,
            I => \N__50831\
        );

    \I__12328\ : ClkMux
    port map (
            O => \N__51387\,
            I => \N__50831\
        );

    \I__12327\ : ClkMux
    port map (
            O => \N__51386\,
            I => \N__50831\
        );

    \I__12326\ : ClkMux
    port map (
            O => \N__51385\,
            I => \N__50831\
        );

    \I__12325\ : ClkMux
    port map (
            O => \N__51384\,
            I => \N__50831\
        );

    \I__12324\ : ClkMux
    port map (
            O => \N__51383\,
            I => \N__50831\
        );

    \I__12323\ : ClkMux
    port map (
            O => \N__51382\,
            I => \N__50831\
        );

    \I__12322\ : ClkMux
    port map (
            O => \N__51381\,
            I => \N__50831\
        );

    \I__12321\ : ClkMux
    port map (
            O => \N__51380\,
            I => \N__50831\
        );

    \I__12320\ : ClkMux
    port map (
            O => \N__51379\,
            I => \N__50831\
        );

    \I__12319\ : ClkMux
    port map (
            O => \N__51378\,
            I => \N__50831\
        );

    \I__12318\ : ClkMux
    port map (
            O => \N__51377\,
            I => \N__50831\
        );

    \I__12317\ : ClkMux
    port map (
            O => \N__51376\,
            I => \N__50831\
        );

    \I__12316\ : ClkMux
    port map (
            O => \N__51375\,
            I => \N__50831\
        );

    \I__12315\ : ClkMux
    port map (
            O => \N__51374\,
            I => \N__50831\
        );

    \I__12314\ : ClkMux
    port map (
            O => \N__51373\,
            I => \N__50831\
        );

    \I__12313\ : ClkMux
    port map (
            O => \N__51372\,
            I => \N__50831\
        );

    \I__12312\ : ClkMux
    port map (
            O => \N__51371\,
            I => \N__50831\
        );

    \I__12311\ : ClkMux
    port map (
            O => \N__51370\,
            I => \N__50831\
        );

    \I__12310\ : ClkMux
    port map (
            O => \N__51369\,
            I => \N__50831\
        );

    \I__12309\ : ClkMux
    port map (
            O => \N__51368\,
            I => \N__50831\
        );

    \I__12308\ : ClkMux
    port map (
            O => \N__51367\,
            I => \N__50831\
        );

    \I__12307\ : ClkMux
    port map (
            O => \N__51366\,
            I => \N__50831\
        );

    \I__12306\ : ClkMux
    port map (
            O => \N__51365\,
            I => \N__50831\
        );

    \I__12305\ : ClkMux
    port map (
            O => \N__51364\,
            I => \N__50831\
        );

    \I__12304\ : ClkMux
    port map (
            O => \N__51363\,
            I => \N__50831\
        );

    \I__12303\ : ClkMux
    port map (
            O => \N__51362\,
            I => \N__50831\
        );

    \I__12302\ : ClkMux
    port map (
            O => \N__51361\,
            I => \N__50831\
        );

    \I__12301\ : ClkMux
    port map (
            O => \N__51360\,
            I => \N__50831\
        );

    \I__12300\ : ClkMux
    port map (
            O => \N__51359\,
            I => \N__50831\
        );

    \I__12299\ : ClkMux
    port map (
            O => \N__51358\,
            I => \N__50831\
        );

    \I__12298\ : ClkMux
    port map (
            O => \N__51357\,
            I => \N__50831\
        );

    \I__12297\ : ClkMux
    port map (
            O => \N__51356\,
            I => \N__50831\
        );

    \I__12296\ : ClkMux
    port map (
            O => \N__51355\,
            I => \N__50831\
        );

    \I__12295\ : ClkMux
    port map (
            O => \N__51354\,
            I => \N__50831\
        );

    \I__12294\ : ClkMux
    port map (
            O => \N__51353\,
            I => \N__50831\
        );

    \I__12293\ : ClkMux
    port map (
            O => \N__51352\,
            I => \N__50831\
        );

    \I__12292\ : ClkMux
    port map (
            O => \N__51351\,
            I => \N__50831\
        );

    \I__12291\ : ClkMux
    port map (
            O => \N__51350\,
            I => \N__50831\
        );

    \I__12290\ : ClkMux
    port map (
            O => \N__51349\,
            I => \N__50831\
        );

    \I__12289\ : ClkMux
    port map (
            O => \N__51348\,
            I => \N__50831\
        );

    \I__12288\ : ClkMux
    port map (
            O => \N__51347\,
            I => \N__50831\
        );

    \I__12287\ : ClkMux
    port map (
            O => \N__51346\,
            I => \N__50831\
        );

    \I__12286\ : ClkMux
    port map (
            O => \N__51345\,
            I => \N__50831\
        );

    \I__12285\ : ClkMux
    port map (
            O => \N__51344\,
            I => \N__50831\
        );

    \I__12284\ : ClkMux
    port map (
            O => \N__51343\,
            I => \N__50831\
        );

    \I__12283\ : ClkMux
    port map (
            O => \N__51342\,
            I => \N__50831\
        );

    \I__12282\ : ClkMux
    port map (
            O => \N__51341\,
            I => \N__50831\
        );

    \I__12281\ : ClkMux
    port map (
            O => \N__51340\,
            I => \N__50831\
        );

    \I__12280\ : ClkMux
    port map (
            O => \N__51339\,
            I => \N__50831\
        );

    \I__12279\ : ClkMux
    port map (
            O => \N__51338\,
            I => \N__50831\
        );

    \I__12278\ : ClkMux
    port map (
            O => \N__51337\,
            I => \N__50831\
        );

    \I__12277\ : ClkMux
    port map (
            O => \N__51336\,
            I => \N__50831\
        );

    \I__12276\ : ClkMux
    port map (
            O => \N__51335\,
            I => \N__50831\
        );

    \I__12275\ : ClkMux
    port map (
            O => \N__51334\,
            I => \N__50831\
        );

    \I__12274\ : ClkMux
    port map (
            O => \N__51333\,
            I => \N__50831\
        );

    \I__12273\ : ClkMux
    port map (
            O => \N__51332\,
            I => \N__50831\
        );

    \I__12272\ : ClkMux
    port map (
            O => \N__51331\,
            I => \N__50831\
        );

    \I__12271\ : ClkMux
    port map (
            O => \N__51330\,
            I => \N__50831\
        );

    \I__12270\ : ClkMux
    port map (
            O => \N__51329\,
            I => \N__50831\
        );

    \I__12269\ : ClkMux
    port map (
            O => \N__51328\,
            I => \N__50831\
        );

    \I__12268\ : ClkMux
    port map (
            O => \N__51327\,
            I => \N__50831\
        );

    \I__12267\ : ClkMux
    port map (
            O => \N__51326\,
            I => \N__50831\
        );

    \I__12266\ : ClkMux
    port map (
            O => \N__51325\,
            I => \N__50831\
        );

    \I__12265\ : ClkMux
    port map (
            O => \N__51324\,
            I => \N__50831\
        );

    \I__12264\ : ClkMux
    port map (
            O => \N__51323\,
            I => \N__50831\
        );

    \I__12263\ : ClkMux
    port map (
            O => \N__51322\,
            I => \N__50831\
        );

    \I__12262\ : ClkMux
    port map (
            O => \N__51321\,
            I => \N__50831\
        );

    \I__12261\ : ClkMux
    port map (
            O => \N__51320\,
            I => \N__50831\
        );

    \I__12260\ : ClkMux
    port map (
            O => \N__51319\,
            I => \N__50831\
        );

    \I__12259\ : ClkMux
    port map (
            O => \N__51318\,
            I => \N__50831\
        );

    \I__12258\ : ClkMux
    port map (
            O => \N__51317\,
            I => \N__50831\
        );

    \I__12257\ : ClkMux
    port map (
            O => \N__51316\,
            I => \N__50831\
        );

    \I__12256\ : ClkMux
    port map (
            O => \N__51315\,
            I => \N__50831\
        );

    \I__12255\ : ClkMux
    port map (
            O => \N__51314\,
            I => \N__50831\
        );

    \I__12254\ : ClkMux
    port map (
            O => \N__51313\,
            I => \N__50831\
        );

    \I__12253\ : ClkMux
    port map (
            O => \N__51312\,
            I => \N__50831\
        );

    \I__12252\ : ClkMux
    port map (
            O => \N__51311\,
            I => \N__50831\
        );

    \I__12251\ : ClkMux
    port map (
            O => \N__51310\,
            I => \N__50831\
        );

    \I__12250\ : ClkMux
    port map (
            O => \N__51309\,
            I => \N__50831\
        );

    \I__12249\ : ClkMux
    port map (
            O => \N__51308\,
            I => \N__50831\
        );

    \I__12248\ : ClkMux
    port map (
            O => \N__51307\,
            I => \N__50831\
        );

    \I__12247\ : ClkMux
    port map (
            O => \N__51306\,
            I => \N__50831\
        );

    \I__12246\ : GlobalMux
    port map (
            O => \N__50831\,
            I => \N__50828\
        );

    \I__12245\ : gio2CtrlBuf
    port map (
            O => \N__50828\,
            I => clk_system_c_g
        );

    \I__12244\ : InMux
    port map (
            O => \N__50825\,
            I => \N__50788\
        );

    \I__12243\ : InMux
    port map (
            O => \N__50824\,
            I => \N__50788\
        );

    \I__12242\ : InMux
    port map (
            O => \N__50823\,
            I => \N__50788\
        );

    \I__12241\ : InMux
    port map (
            O => \N__50822\,
            I => \N__50781\
        );

    \I__12240\ : InMux
    port map (
            O => \N__50821\,
            I => \N__50781\
        );

    \I__12239\ : InMux
    port map (
            O => \N__50820\,
            I => \N__50781\
        );

    \I__12238\ : InMux
    port map (
            O => \N__50819\,
            I => \N__50776\
        );

    \I__12237\ : InMux
    port map (
            O => \N__50818\,
            I => \N__50776\
        );

    \I__12236\ : InMux
    port map (
            O => \N__50817\,
            I => \N__50773\
        );

    \I__12235\ : InMux
    port map (
            O => \N__50816\,
            I => \N__50762\
        );

    \I__12234\ : InMux
    port map (
            O => \N__50815\,
            I => \N__50762\
        );

    \I__12233\ : InMux
    port map (
            O => \N__50814\,
            I => \N__50762\
        );

    \I__12232\ : InMux
    port map (
            O => \N__50813\,
            I => \N__50762\
        );

    \I__12231\ : InMux
    port map (
            O => \N__50812\,
            I => \N__50762\
        );

    \I__12230\ : InMux
    port map (
            O => \N__50811\,
            I => \N__50755\
        );

    \I__12229\ : InMux
    port map (
            O => \N__50810\,
            I => \N__50755\
        );

    \I__12228\ : InMux
    port map (
            O => \N__50809\,
            I => \N__50755\
        );

    \I__12227\ : InMux
    port map (
            O => \N__50808\,
            I => \N__50746\
        );

    \I__12226\ : InMux
    port map (
            O => \N__50807\,
            I => \N__50746\
        );

    \I__12225\ : InMux
    port map (
            O => \N__50806\,
            I => \N__50746\
        );

    \I__12224\ : InMux
    port map (
            O => \N__50805\,
            I => \N__50746\
        );

    \I__12223\ : InMux
    port map (
            O => \N__50804\,
            I => \N__50741\
        );

    \I__12222\ : InMux
    port map (
            O => \N__50803\,
            I => \N__50741\
        );

    \I__12221\ : InMux
    port map (
            O => \N__50802\,
            I => \N__50738\
        );

    \I__12220\ : InMux
    port map (
            O => \N__50801\,
            I => \N__50735\
        );

    \I__12219\ : InMux
    port map (
            O => \N__50800\,
            I => \N__50730\
        );

    \I__12218\ : InMux
    port map (
            O => \N__50799\,
            I => \N__50730\
        );

    \I__12217\ : InMux
    port map (
            O => \N__50798\,
            I => \N__50727\
        );

    \I__12216\ : InMux
    port map (
            O => \N__50797\,
            I => \N__50724\
        );

    \I__12215\ : InMux
    port map (
            O => \N__50796\,
            I => \N__50721\
        );

    \I__12214\ : InMux
    port map (
            O => \N__50795\,
            I => \N__50718\
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__50788\,
            I => \N__50687\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__50781\,
            I => \N__50684\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__50776\,
            I => \N__50681\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__50773\,
            I => \N__50678\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__50762\,
            I => \N__50675\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__50755\,
            I => \N__50672\
        );

    \I__12207\ : LocalMux
    port map (
            O => \N__50746\,
            I => \N__50669\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__50741\,
            I => \N__50666\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__50738\,
            I => \N__50663\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__50735\,
            I => \N__50660\
        );

    \I__12203\ : LocalMux
    port map (
            O => \N__50730\,
            I => \N__50657\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__50727\,
            I => \N__50654\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__50724\,
            I => \N__50651\
        );

    \I__12200\ : LocalMux
    port map (
            O => \N__50721\,
            I => \N__50648\
        );

    \I__12199\ : LocalMux
    port map (
            O => \N__50718\,
            I => \N__50645\
        );

    \I__12198\ : SRMux
    port map (
            O => \N__50717\,
            I => \N__50558\
        );

    \I__12197\ : SRMux
    port map (
            O => \N__50716\,
            I => \N__50558\
        );

    \I__12196\ : SRMux
    port map (
            O => \N__50715\,
            I => \N__50558\
        );

    \I__12195\ : SRMux
    port map (
            O => \N__50714\,
            I => \N__50558\
        );

    \I__12194\ : SRMux
    port map (
            O => \N__50713\,
            I => \N__50558\
        );

    \I__12193\ : SRMux
    port map (
            O => \N__50712\,
            I => \N__50558\
        );

    \I__12192\ : SRMux
    port map (
            O => \N__50711\,
            I => \N__50558\
        );

    \I__12191\ : SRMux
    port map (
            O => \N__50710\,
            I => \N__50558\
        );

    \I__12190\ : SRMux
    port map (
            O => \N__50709\,
            I => \N__50558\
        );

    \I__12189\ : SRMux
    port map (
            O => \N__50708\,
            I => \N__50558\
        );

    \I__12188\ : SRMux
    port map (
            O => \N__50707\,
            I => \N__50558\
        );

    \I__12187\ : SRMux
    port map (
            O => \N__50706\,
            I => \N__50558\
        );

    \I__12186\ : SRMux
    port map (
            O => \N__50705\,
            I => \N__50558\
        );

    \I__12185\ : SRMux
    port map (
            O => \N__50704\,
            I => \N__50558\
        );

    \I__12184\ : SRMux
    port map (
            O => \N__50703\,
            I => \N__50558\
        );

    \I__12183\ : SRMux
    port map (
            O => \N__50702\,
            I => \N__50558\
        );

    \I__12182\ : SRMux
    port map (
            O => \N__50701\,
            I => \N__50558\
        );

    \I__12181\ : SRMux
    port map (
            O => \N__50700\,
            I => \N__50558\
        );

    \I__12180\ : SRMux
    port map (
            O => \N__50699\,
            I => \N__50558\
        );

    \I__12179\ : SRMux
    port map (
            O => \N__50698\,
            I => \N__50558\
        );

    \I__12178\ : SRMux
    port map (
            O => \N__50697\,
            I => \N__50558\
        );

    \I__12177\ : SRMux
    port map (
            O => \N__50696\,
            I => \N__50558\
        );

    \I__12176\ : SRMux
    port map (
            O => \N__50695\,
            I => \N__50558\
        );

    \I__12175\ : SRMux
    port map (
            O => \N__50694\,
            I => \N__50558\
        );

    \I__12174\ : SRMux
    port map (
            O => \N__50693\,
            I => \N__50558\
        );

    \I__12173\ : SRMux
    port map (
            O => \N__50692\,
            I => \N__50558\
        );

    \I__12172\ : SRMux
    port map (
            O => \N__50691\,
            I => \N__50558\
        );

    \I__12171\ : SRMux
    port map (
            O => \N__50690\,
            I => \N__50558\
        );

    \I__12170\ : Glb2LocalMux
    port map (
            O => \N__50687\,
            I => \N__50558\
        );

    \I__12169\ : Glb2LocalMux
    port map (
            O => \N__50684\,
            I => \N__50558\
        );

    \I__12168\ : Glb2LocalMux
    port map (
            O => \N__50681\,
            I => \N__50558\
        );

    \I__12167\ : Glb2LocalMux
    port map (
            O => \N__50678\,
            I => \N__50558\
        );

    \I__12166\ : Glb2LocalMux
    port map (
            O => \N__50675\,
            I => \N__50558\
        );

    \I__12165\ : Glb2LocalMux
    port map (
            O => \N__50672\,
            I => \N__50558\
        );

    \I__12164\ : Glb2LocalMux
    port map (
            O => \N__50669\,
            I => \N__50558\
        );

    \I__12163\ : Glb2LocalMux
    port map (
            O => \N__50666\,
            I => \N__50558\
        );

    \I__12162\ : Glb2LocalMux
    port map (
            O => \N__50663\,
            I => \N__50558\
        );

    \I__12161\ : Glb2LocalMux
    port map (
            O => \N__50660\,
            I => \N__50558\
        );

    \I__12160\ : Glb2LocalMux
    port map (
            O => \N__50657\,
            I => \N__50558\
        );

    \I__12159\ : Glb2LocalMux
    port map (
            O => \N__50654\,
            I => \N__50558\
        );

    \I__12158\ : Glb2LocalMux
    port map (
            O => \N__50651\,
            I => \N__50558\
        );

    \I__12157\ : Glb2LocalMux
    port map (
            O => \N__50648\,
            I => \N__50558\
        );

    \I__12156\ : Glb2LocalMux
    port map (
            O => \N__50645\,
            I => \N__50558\
        );

    \I__12155\ : GlobalMux
    port map (
            O => \N__50558\,
            I => \N__50555\
        );

    \I__12154\ : gio2CtrlBuf
    port map (
            O => \N__50555\,
            I => \N_851_g\
        );

    \I__12153\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50549\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__50549\,
            I => \N__50546\
        );

    \I__12151\ : Odrv4
    port map (
            O => \N__50546\,
            I => \pid_front.O_18\
        );

    \I__12150\ : InMux
    port map (
            O => \N__50543\,
            I => \N__50540\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__50540\,
            I => \N__50536\
        );

    \I__12148\ : InMux
    port map (
            O => \N__50539\,
            I => \N__50533\
        );

    \I__12147\ : Span4Mux_h
    port map (
            O => \N__50536\,
            I => \N__50530\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__50533\,
            I => \N__50527\
        );

    \I__12145\ : Span4Mux_h
    port map (
            O => \N__50530\,
            I => \N__50524\
        );

    \I__12144\ : Span4Mux_h
    port map (
            O => \N__50527\,
            I => \N__50520\
        );

    \I__12143\ : Span4Mux_h
    port map (
            O => \N__50524\,
            I => \N__50517\
        );

    \I__12142\ : InMux
    port map (
            O => \N__50523\,
            I => \N__50514\
        );

    \I__12141\ : Span4Mux_h
    port map (
            O => \N__50520\,
            I => \N__50511\
        );

    \I__12140\ : Odrv4
    port map (
            O => \N__50517\,
            I => \pid_front.error_p_regZ0Z_14\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__50514\,
            I => \pid_front.error_p_regZ0Z_14\
        );

    \I__12138\ : Odrv4
    port map (
            O => \N__50511\,
            I => \pid_front.error_p_regZ0Z_14\
        );

    \I__12137\ : InMux
    port map (
            O => \N__50504\,
            I => \N__50501\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__50501\,
            I => \N__50498\
        );

    \I__12135\ : Odrv4
    port map (
            O => \N__50498\,
            I => \pid_front.O_12\
        );

    \I__12134\ : InMux
    port map (
            O => \N__50495\,
            I => \N__50492\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__50492\,
            I => \N__50488\
        );

    \I__12132\ : InMux
    port map (
            O => \N__50491\,
            I => \N__50485\
        );

    \I__12131\ : Span4Mux_v
    port map (
            O => \N__50488\,
            I => \N__50479\
        );

    \I__12130\ : LocalMux
    port map (
            O => \N__50485\,
            I => \N__50479\
        );

    \I__12129\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50476\
        );

    \I__12128\ : Span4Mux_h
    port map (
            O => \N__50479\,
            I => \N__50473\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__50476\,
            I => \pid_front.error_p_regZ0Z_8\
        );

    \I__12126\ : Odrv4
    port map (
            O => \N__50473\,
            I => \pid_front.error_p_regZ0Z_8\
        );

    \I__12125\ : InMux
    port map (
            O => \N__50468\,
            I => \N__50465\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__50465\,
            I => \N__50462\
        );

    \I__12123\ : Odrv4
    port map (
            O => \N__50462\,
            I => \pid_front.O_14\
        );

    \I__12122\ : InMux
    port map (
            O => \N__50459\,
            I => \N__50456\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__50456\,
            I => \N__50453\
        );

    \I__12120\ : Span4Mux_v
    port map (
            O => \N__50453\,
            I => \N__50449\
        );

    \I__12119\ : InMux
    port map (
            O => \N__50452\,
            I => \N__50446\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__50449\,
            I => \N__50442\
        );

    \I__12117\ : LocalMux
    port map (
            O => \N__50446\,
            I => \N__50439\
        );

    \I__12116\ : InMux
    port map (
            O => \N__50445\,
            I => \N__50436\
        );

    \I__12115\ : Sp12to4
    port map (
            O => \N__50442\,
            I => \N__50431\
        );

    \I__12114\ : Span12Mux_s8_v
    port map (
            O => \N__50439\,
            I => \N__50431\
        );

    \I__12113\ : LocalMux
    port map (
            O => \N__50436\,
            I => \pid_front.error_p_regZ0Z_10\
        );

    \I__12112\ : Odrv12
    port map (
            O => \N__50431\,
            I => \pid_front.error_p_regZ0Z_10\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50426\,
            I => \N__50423\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__50423\,
            I => \N__50420\
        );

    \I__12109\ : Odrv4
    port map (
            O => \N__50420\,
            I => \pid_front.O_11\
        );

    \I__12108\ : InMux
    port map (
            O => \N__50417\,
            I => \N__50413\
        );

    \I__12107\ : CascadeMux
    port map (
            O => \N__50416\,
            I => \N__50410\
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__50413\,
            I => \N__50406\
        );

    \I__12105\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50403\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50400\
        );

    \I__12103\ : Span12Mux_h
    port map (
            O => \N__50406\,
            I => \N__50395\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__50403\,
            I => \N__50395\
        );

    \I__12101\ : LocalMux
    port map (
            O => \N__50400\,
            I => \pid_front.error_p_regZ0Z_7\
        );

    \I__12100\ : Odrv12
    port map (
            O => \N__50395\,
            I => \pid_front.error_p_regZ0Z_7\
        );

    \I__12099\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50387\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__50387\,
            I => \pid_front.O_7\
        );

    \I__12097\ : InMux
    port map (
            O => \N__50384\,
            I => \N__50381\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__50381\,
            I => \N__50378\
        );

    \I__12095\ : Span4Mux_h
    port map (
            O => \N__50378\,
            I => \N__50374\
        );

    \I__12094\ : InMux
    port map (
            O => \N__50377\,
            I => \N__50370\
        );

    \I__12093\ : Span4Mux_h
    port map (
            O => \N__50374\,
            I => \N__50367\
        );

    \I__12092\ : InMux
    port map (
            O => \N__50373\,
            I => \N__50364\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__50370\,
            I => \N__50361\
        );

    \I__12090\ : Odrv4
    port map (
            O => \N__50367\,
            I => \pid_front.error_p_regZ0Z_3\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__50364\,
            I => \pid_front.error_p_regZ0Z_3\
        );

    \I__12088\ : Odrv12
    port map (
            O => \N__50361\,
            I => \pid_front.error_p_regZ0Z_3\
        );

    \I__12087\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50351\
        );

    \I__12086\ : LocalMux
    port map (
            O => \N__50351\,
            I => \N__50348\
        );

    \I__12085\ : Odrv4
    port map (
            O => \N__50348\,
            I => \pid_front.O_20\
        );

    \I__12084\ : InMux
    port map (
            O => \N__50345\,
            I => \N__50342\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__50342\,
            I => \N__50338\
        );

    \I__12082\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50335\
        );

    \I__12081\ : Span4Mux_h
    port map (
            O => \N__50338\,
            I => \N__50329\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__50335\,
            I => \N__50329\
        );

    \I__12079\ : InMux
    port map (
            O => \N__50334\,
            I => \N__50326\
        );

    \I__12078\ : Span4Mux_h
    port map (
            O => \N__50329\,
            I => \N__50323\
        );

    \I__12077\ : LocalMux
    port map (
            O => \N__50326\,
            I => \pid_front.error_p_regZ0Z_16\
        );

    \I__12076\ : Odrv4
    port map (
            O => \N__50323\,
            I => \pid_front.error_p_regZ0Z_16\
        );

    \I__12075\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50315\
        );

    \I__12074\ : LocalMux
    port map (
            O => \N__50315\,
            I => \pid_front.O_10\
        );

    \I__12073\ : InMux
    port map (
            O => \N__50312\,
            I => \N__50308\
        );

    \I__12072\ : CascadeMux
    port map (
            O => \N__50311\,
            I => \N__50305\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__50308\,
            I => \N__50302\
        );

    \I__12070\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50299\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__50302\,
            I => \N__50296\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__50299\,
            I => \N__50293\
        );

    \I__12067\ : Span4Mux_h
    port map (
            O => \N__50296\,
            I => \N__50289\
        );

    \I__12066\ : Span4Mux_v
    port map (
            O => \N__50293\,
            I => \N__50286\
        );

    \I__12065\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50283\
        );

    \I__12064\ : Span4Mux_h
    port map (
            O => \N__50289\,
            I => \N__50278\
        );

    \I__12063\ : Span4Mux_h
    port map (
            O => \N__50286\,
            I => \N__50278\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__50283\,
            I => \pid_front.error_p_regZ0Z_6\
        );

    \I__12061\ : Odrv4
    port map (
            O => \N__50278\,
            I => \pid_front.error_p_regZ0Z_6\
        );

    \I__12060\ : InMux
    port map (
            O => \N__50273\,
            I => \N__50270\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__50270\,
            I => \N__50267\
        );

    \I__12058\ : Odrv4
    port map (
            O => \N__50267\,
            I => \pid_front.O_22\
        );

    \I__12057\ : CascadeMux
    port map (
            O => \N__50264\,
            I => \N__50261\
        );

    \I__12056\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50258\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__50258\,
            I => \N__50255\
        );

    \I__12054\ : Span4Mux_v
    port map (
            O => \N__50255\,
            I => \N__50252\
        );

    \I__12053\ : Span4Mux_h
    port map (
            O => \N__50252\,
            I => \N__50248\
        );

    \I__12052\ : InMux
    port map (
            O => \N__50251\,
            I => \N__50245\
        );

    \I__12051\ : Sp12to4
    port map (
            O => \N__50248\,
            I => \N__50239\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__50245\,
            I => \N__50239\
        );

    \I__12049\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50236\
        );

    \I__12048\ : Span12Mux_s7_v
    port map (
            O => \N__50239\,
            I => \N__50233\
        );

    \I__12047\ : LocalMux
    port map (
            O => \N__50236\,
            I => \pid_front.error_p_regZ0Z_18\
        );

    \I__12046\ : Odrv12
    port map (
            O => \N__50233\,
            I => \pid_front.error_p_regZ0Z_18\
        );

    \I__12045\ : CascadeMux
    port map (
            O => \N__50228\,
            I => \N__50223\
        );

    \I__12044\ : CascadeMux
    port map (
            O => \N__50227\,
            I => \N__50219\
        );

    \I__12043\ : CascadeMux
    port map (
            O => \N__50226\,
            I => \N__50209\
        );

    \I__12042\ : InMux
    port map (
            O => \N__50223\,
            I => \N__50197\
        );

    \I__12041\ : InMux
    port map (
            O => \N__50222\,
            I => \N__50197\
        );

    \I__12040\ : InMux
    port map (
            O => \N__50219\,
            I => \N__50180\
        );

    \I__12039\ : InMux
    port map (
            O => \N__50218\,
            I => \N__50180\
        );

    \I__12038\ : InMux
    port map (
            O => \N__50217\,
            I => \N__50180\
        );

    \I__12037\ : InMux
    port map (
            O => \N__50216\,
            I => \N__50180\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50215\,
            I => \N__50180\
        );

    \I__12035\ : InMux
    port map (
            O => \N__50214\,
            I => \N__50180\
        );

    \I__12034\ : InMux
    port map (
            O => \N__50213\,
            I => \N__50180\
        );

    \I__12033\ : InMux
    port map (
            O => \N__50212\,
            I => \N__50180\
        );

    \I__12032\ : InMux
    port map (
            O => \N__50209\,
            I => \N__50160\
        );

    \I__12031\ : InMux
    port map (
            O => \N__50208\,
            I => \N__50160\
        );

    \I__12030\ : InMux
    port map (
            O => \N__50207\,
            I => \N__50160\
        );

    \I__12029\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50160\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50160\
        );

    \I__12027\ : InMux
    port map (
            O => \N__50204\,
            I => \N__50160\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50203\,
            I => \N__50160\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50202\,
            I => \N__50160\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__50197\,
            I => \N__50155\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50180\,
            I => \N__50155\
        );

    \I__12022\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50152\
        );

    \I__12021\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50147\
        );

    \I__12020\ : InMux
    port map (
            O => \N__50177\,
            I => \N__50147\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__50160\,
            I => \N__50144\
        );

    \I__12018\ : Span4Mux_v
    port map (
            O => \N__50155\,
            I => \N__50141\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50136\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__50147\,
            I => \N__50136\
        );

    \I__12015\ : Span12Mux_s3_h
    port map (
            O => \N__50144\,
            I => \N__50131\
        );

    \I__12014\ : Sp12to4
    port map (
            O => \N__50141\,
            I => \N__50131\
        );

    \I__12013\ : Odrv12
    port map (
            O => \N__50136\,
            I => \pid_side.state_RNINK4UZ0Z_1\
        );

    \I__12012\ : Odrv12
    port map (
            O => \N__50131\,
            I => \pid_side.state_RNINK4UZ0Z_1\
        );

    \I__12011\ : InMux
    port map (
            O => \N__50126\,
            I => \N__50123\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__50123\,
            I => \N__50120\
        );

    \I__12009\ : Span12Mux_h
    port map (
            O => \N__50120\,
            I => \N__50117\
        );

    \I__12008\ : Odrv12
    port map (
            O => \N__50117\,
            I => \pid_side.O_0_7\
        );

    \I__12007\ : InMux
    port map (
            O => \N__50114\,
            I => \N__50111\
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__50111\,
            I => \N__50108\
        );

    \I__12005\ : Span4Mux_h
    port map (
            O => \N__50108\,
            I => \N__50104\
        );

    \I__12004\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50101\
        );

    \I__12003\ : Sp12to4
    port map (
            O => \N__50104\,
            I => \N__50096\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50101\,
            I => \N__50096\
        );

    \I__12001\ : Span12Mux_v
    port map (
            O => \N__50096\,
            I => \N__50092\
        );

    \I__12000\ : InMux
    port map (
            O => \N__50095\,
            I => \N__50089\
        );

    \I__11999\ : Span12Mux_h
    port map (
            O => \N__50092\,
            I => \N__50086\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50089\,
            I => \pid_side.error_p_regZ0Z_3\
        );

    \I__11997\ : Odrv12
    port map (
            O => \N__50086\,
            I => \pid_side.error_p_regZ0Z_3\
        );

    \I__11996\ : InMux
    port map (
            O => \N__50081\,
            I => \N__50078\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50078\,
            I => \N__50075\
        );

    \I__11994\ : Odrv12
    port map (
            O => \N__50075\,
            I => \pid_front.O_4\
        );

    \I__11993\ : InMux
    port map (
            O => \N__50072\,
            I => \N__50069\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__50069\,
            I => \N__50066\
        );

    \I__11991\ : Span4Mux_v
    port map (
            O => \N__50066\,
            I => \N__50063\
        );

    \I__11990\ : Span4Mux_v
    port map (
            O => \N__50063\,
            I => \N__50060\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__50060\,
            I => \N__50056\
        );

    \I__11988\ : InMux
    port map (
            O => \N__50059\,
            I => \N__50053\
        );

    \I__11987\ : Odrv4
    port map (
            O => \N__50056\,
            I => \pid_front.error_p_regZ0Z_0\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__50053\,
            I => \pid_front.error_p_regZ0Z_0\
        );

    \I__11985\ : InMux
    port map (
            O => \N__50048\,
            I => \N__50041\
        );

    \I__11984\ : CascadeMux
    port map (
            O => \N__50047\,
            I => \N__50036\
        );

    \I__11983\ : CascadeMux
    port map (
            O => \N__50046\,
            I => \N__50031\
        );

    \I__11982\ : CascadeMux
    port map (
            O => \N__50045\,
            I => \N__50028\
        );

    \I__11981\ : CascadeMux
    port map (
            O => \N__50044\,
            I => \N__50024\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50041\,
            I => \N__50016\
        );

    \I__11979\ : CascadeMux
    port map (
            O => \N__50040\,
            I => \N__50013\
        );

    \I__11978\ : CascadeMux
    port map (
            O => \N__50039\,
            I => \N__50009\
        );

    \I__11977\ : InMux
    port map (
            O => \N__50036\,
            I => \N__50006\
        );

    \I__11976\ : InMux
    port map (
            O => \N__50035\,
            I => \N__50003\
        );

    \I__11975\ : InMux
    port map (
            O => \N__50034\,
            I => \N__49996\
        );

    \I__11974\ : InMux
    port map (
            O => \N__50031\,
            I => \N__49996\
        );

    \I__11973\ : InMux
    port map (
            O => \N__50028\,
            I => \N__49996\
        );

    \I__11972\ : InMux
    port map (
            O => \N__50027\,
            I => \N__49989\
        );

    \I__11971\ : InMux
    port map (
            O => \N__50024\,
            I => \N__49989\
        );

    \I__11970\ : InMux
    port map (
            O => \N__50023\,
            I => \N__49989\
        );

    \I__11969\ : CascadeMux
    port map (
            O => \N__50022\,
            I => \N__49986\
        );

    \I__11968\ : CascadeMux
    port map (
            O => \N__50021\,
            I => \N__49982\
        );

    \I__11967\ : CascadeMux
    port map (
            O => \N__50020\,
            I => \N__49979\
        );

    \I__11966\ : InMux
    port map (
            O => \N__50019\,
            I => \N__49971\
        );

    \I__11965\ : Span4Mux_h
    port map (
            O => \N__50016\,
            I => \N__49968\
        );

    \I__11964\ : InMux
    port map (
            O => \N__50013\,
            I => \N__49963\
        );

    \I__11963\ : InMux
    port map (
            O => \N__50012\,
            I => \N__49963\
        );

    \I__11962\ : InMux
    port map (
            O => \N__50009\,
            I => \N__49960\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__50006\,
            I => \N__49957\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__50003\,
            I => \N__49950\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__49996\,
            I => \N__49950\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__49989\,
            I => \N__49950\
        );

    \I__11957\ : InMux
    port map (
            O => \N__49986\,
            I => \N__49945\
        );

    \I__11956\ : InMux
    port map (
            O => \N__49985\,
            I => \N__49945\
        );

    \I__11955\ : InMux
    port map (
            O => \N__49982\,
            I => \N__49940\
        );

    \I__11954\ : InMux
    port map (
            O => \N__49979\,
            I => \N__49940\
        );

    \I__11953\ : CascadeMux
    port map (
            O => \N__49978\,
            I => \N__49937\
        );

    \I__11952\ : CascadeMux
    port map (
            O => \N__49977\,
            I => \N__49934\
        );

    \I__11951\ : CascadeMux
    port map (
            O => \N__49976\,
            I => \N__49931\
        );

    \I__11950\ : CascadeMux
    port map (
            O => \N__49975\,
            I => \N__49927\
        );

    \I__11949\ : InMux
    port map (
            O => \N__49974\,
            I => \N__49923\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__49971\,
            I => \N__49918\
        );

    \I__11947\ : Span4Mux_h
    port map (
            O => \N__49968\,
            I => \N__49918\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__49963\,
            I => \N__49915\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__49960\,
            I => \N__49912\
        );

    \I__11944\ : Span4Mux_v
    port map (
            O => \N__49957\,
            I => \N__49903\
        );

    \I__11943\ : Span4Mux_v
    port map (
            O => \N__49950\,
            I => \N__49903\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__49945\,
            I => \N__49903\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__49940\,
            I => \N__49903\
        );

    \I__11940\ : InMux
    port map (
            O => \N__49937\,
            I => \N__49900\
        );

    \I__11939\ : InMux
    port map (
            O => \N__49934\,
            I => \N__49891\
        );

    \I__11938\ : InMux
    port map (
            O => \N__49931\,
            I => \N__49891\
        );

    \I__11937\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49891\
        );

    \I__11936\ : InMux
    port map (
            O => \N__49927\,
            I => \N__49891\
        );

    \I__11935\ : InMux
    port map (
            O => \N__49926\,
            I => \N__49888\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__49923\,
            I => \N__49881\
        );

    \I__11933\ : Span4Mux_h
    port map (
            O => \N__49918\,
            I => \N__49881\
        );

    \I__11932\ : Span4Mux_h
    port map (
            O => \N__49915\,
            I => \N__49881\
        );

    \I__11931\ : Odrv12
    port map (
            O => \N__49912\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11930\ : Odrv4
    port map (
            O => \N__49903\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__49900\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__49891\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__49888\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11926\ : Odrv4
    port map (
            O => \N__49881\,
            I => \pid_side.stateZ0Z_0\
        );

    \I__11925\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49864\
        );

    \I__11924\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49861\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__49864\,
            I => \N__49858\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__49861\,
            I => \N__49855\
        );

    \I__11921\ : Span4Mux_v
    port map (
            O => \N__49858\,
            I => \N__49851\
        );

    \I__11920\ : Span4Mux_v
    port map (
            O => \N__49855\,
            I => \N__49848\
        );

    \I__11919\ : InMux
    port map (
            O => \N__49854\,
            I => \N__49845\
        );

    \I__11918\ : Sp12to4
    port map (
            O => \N__49851\,
            I => \N__49842\
        );

    \I__11917\ : Odrv4
    port map (
            O => \N__49848\,
            I => \pid_side.error_p_regZ0Z_1\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__49845\,
            I => \pid_side.error_p_regZ0Z_1\
        );

    \I__11915\ : Odrv12
    port map (
            O => \N__49842\,
            I => \pid_side.error_p_regZ0Z_1\
        );

    \I__11914\ : CascadeMux
    port map (
            O => \N__49835\,
            I => \N__49832\
        );

    \I__11913\ : InMux
    port map (
            O => \N__49832\,
            I => \N__49827\
        );

    \I__11912\ : InMux
    port map (
            O => \N__49831\,
            I => \N__49822\
        );

    \I__11911\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49822\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__49827\,
            I => \N__49818\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__49822\,
            I => \N__49815\
        );

    \I__11908\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49812\
        );

    \I__11907\ : Span4Mux_v
    port map (
            O => \N__49818\,
            I => \N__49807\
        );

    \I__11906\ : Span4Mux_h
    port map (
            O => \N__49815\,
            I => \N__49807\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__49812\,
            I => \N__49802\
        );

    \I__11904\ : Span4Mux_h
    port map (
            O => \N__49807\,
            I => \N__49802\
        );

    \I__11903\ : Odrv4
    port map (
            O => \N__49802\,
            I => \pid_side.pid_preregZ0Z_1\
        );

    \I__11902\ : CascadeMux
    port map (
            O => \N__49799\,
            I => \N__49792\
        );

    \I__11901\ : CascadeMux
    port map (
            O => \N__49798\,
            I => \N__49789\
        );

    \I__11900\ : CascadeMux
    port map (
            O => \N__49797\,
            I => \N__49786\
        );

    \I__11899\ : CascadeMux
    port map (
            O => \N__49796\,
            I => \N__49761\
        );

    \I__11898\ : InMux
    port map (
            O => \N__49795\,
            I => \N__49743\
        );

    \I__11897\ : InMux
    port map (
            O => \N__49792\,
            I => \N__49738\
        );

    \I__11896\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49738\
        );

    \I__11895\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49729\
        );

    \I__11894\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49729\
        );

    \I__11893\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49729\
        );

    \I__11892\ : InMux
    port map (
            O => \N__49783\,
            I => \N__49729\
        );

    \I__11891\ : InMux
    port map (
            O => \N__49782\,
            I => \N__49726\
        );

    \I__11890\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49723\
        );

    \I__11889\ : InMux
    port map (
            O => \N__49780\,
            I => \N__49718\
        );

    \I__11888\ : InMux
    port map (
            O => \N__49779\,
            I => \N__49718\
        );

    \I__11887\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49715\
        );

    \I__11886\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49712\
        );

    \I__11885\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49709\
        );

    \I__11884\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49704\
        );

    \I__11883\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49704\
        );

    \I__11882\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49701\
        );

    \I__11881\ : InMux
    port map (
            O => \N__49772\,
            I => \N__49698\
        );

    \I__11880\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49695\
        );

    \I__11879\ : InMux
    port map (
            O => \N__49770\,
            I => \N__49692\
        );

    \I__11878\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49689\
        );

    \I__11877\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49686\
        );

    \I__11876\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49683\
        );

    \I__11875\ : InMux
    port map (
            O => \N__49766\,
            I => \N__49678\
        );

    \I__11874\ : InMux
    port map (
            O => \N__49765\,
            I => \N__49678\
        );

    \I__11873\ : InMux
    port map (
            O => \N__49764\,
            I => \N__49675\
        );

    \I__11872\ : InMux
    port map (
            O => \N__49761\,
            I => \N__49672\
        );

    \I__11871\ : InMux
    port map (
            O => \N__49760\,
            I => \N__49669\
        );

    \I__11870\ : InMux
    port map (
            O => \N__49759\,
            I => \N__49666\
        );

    \I__11869\ : InMux
    port map (
            O => \N__49758\,
            I => \N__49663\
        );

    \I__11868\ : InMux
    port map (
            O => \N__49757\,
            I => \N__49658\
        );

    \I__11867\ : InMux
    port map (
            O => \N__49756\,
            I => \N__49658\
        );

    \I__11866\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49655\
        );

    \I__11865\ : InMux
    port map (
            O => \N__49754\,
            I => \N__49652\
        );

    \I__11864\ : InMux
    port map (
            O => \N__49753\,
            I => \N__49649\
        );

    \I__11863\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49646\
        );

    \I__11862\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49643\
        );

    \I__11861\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49638\
        );

    \I__11860\ : InMux
    port map (
            O => \N__49749\,
            I => \N__49638\
        );

    \I__11859\ : InMux
    port map (
            O => \N__49748\,
            I => \N__49635\
        );

    \I__11858\ : InMux
    port map (
            O => \N__49747\,
            I => \N__49632\
        );

    \I__11857\ : InMux
    port map (
            O => \N__49746\,
            I => \N__49629\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__49743\,
            I => \N__49495\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__49738\,
            I => \N__49492\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__49729\,
            I => \N__49489\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49726\,
            I => \N__49486\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__49723\,
            I => \N__49483\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__49718\,
            I => \N__49480\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__49715\,
            I => \N__49477\
        );

    \I__11849\ : LocalMux
    port map (
            O => \N__49712\,
            I => \N__49474\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__49709\,
            I => \N__49471\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__49704\,
            I => \N__49468\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__49701\,
            I => \N__49465\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__49698\,
            I => \N__49462\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__49695\,
            I => \N__49459\
        );

    \I__11843\ : LocalMux
    port map (
            O => \N__49692\,
            I => \N__49456\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__49689\,
            I => \N__49453\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__49686\,
            I => \N__49450\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__49683\,
            I => \N__49447\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__49678\,
            I => \N__49444\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__49675\,
            I => \N__49441\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__49672\,
            I => \N__49438\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__49669\,
            I => \N__49435\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__49666\,
            I => \N__49432\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__49663\,
            I => \N__49429\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__49658\,
            I => \N__49426\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__49655\,
            I => \N__49423\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__49652\,
            I => \N__49420\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__49649\,
            I => \N__49417\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__49646\,
            I => \N__49414\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__49643\,
            I => \N__49411\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49638\,
            I => \N__49408\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__49635\,
            I => \N__49405\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__49632\,
            I => \N__49402\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__49629\,
            I => \N__49399\
        );

    \I__11823\ : SRMux
    port map (
            O => \N__49628\,
            I => \N__49070\
        );

    \I__11822\ : SRMux
    port map (
            O => \N__49627\,
            I => \N__49070\
        );

    \I__11821\ : SRMux
    port map (
            O => \N__49626\,
            I => \N__49070\
        );

    \I__11820\ : SRMux
    port map (
            O => \N__49625\,
            I => \N__49070\
        );

    \I__11819\ : SRMux
    port map (
            O => \N__49624\,
            I => \N__49070\
        );

    \I__11818\ : SRMux
    port map (
            O => \N__49623\,
            I => \N__49070\
        );

    \I__11817\ : SRMux
    port map (
            O => \N__49622\,
            I => \N__49070\
        );

    \I__11816\ : SRMux
    port map (
            O => \N__49621\,
            I => \N__49070\
        );

    \I__11815\ : SRMux
    port map (
            O => \N__49620\,
            I => \N__49070\
        );

    \I__11814\ : SRMux
    port map (
            O => \N__49619\,
            I => \N__49070\
        );

    \I__11813\ : SRMux
    port map (
            O => \N__49618\,
            I => \N__49070\
        );

    \I__11812\ : SRMux
    port map (
            O => \N__49617\,
            I => \N__49070\
        );

    \I__11811\ : SRMux
    port map (
            O => \N__49616\,
            I => \N__49070\
        );

    \I__11810\ : SRMux
    port map (
            O => \N__49615\,
            I => \N__49070\
        );

    \I__11809\ : SRMux
    port map (
            O => \N__49614\,
            I => \N__49070\
        );

    \I__11808\ : SRMux
    port map (
            O => \N__49613\,
            I => \N__49070\
        );

    \I__11807\ : SRMux
    port map (
            O => \N__49612\,
            I => \N__49070\
        );

    \I__11806\ : SRMux
    port map (
            O => \N__49611\,
            I => \N__49070\
        );

    \I__11805\ : SRMux
    port map (
            O => \N__49610\,
            I => \N__49070\
        );

    \I__11804\ : SRMux
    port map (
            O => \N__49609\,
            I => \N__49070\
        );

    \I__11803\ : SRMux
    port map (
            O => \N__49608\,
            I => \N__49070\
        );

    \I__11802\ : SRMux
    port map (
            O => \N__49607\,
            I => \N__49070\
        );

    \I__11801\ : SRMux
    port map (
            O => \N__49606\,
            I => \N__49070\
        );

    \I__11800\ : SRMux
    port map (
            O => \N__49605\,
            I => \N__49070\
        );

    \I__11799\ : SRMux
    port map (
            O => \N__49604\,
            I => \N__49070\
        );

    \I__11798\ : SRMux
    port map (
            O => \N__49603\,
            I => \N__49070\
        );

    \I__11797\ : SRMux
    port map (
            O => \N__49602\,
            I => \N__49070\
        );

    \I__11796\ : SRMux
    port map (
            O => \N__49601\,
            I => \N__49070\
        );

    \I__11795\ : SRMux
    port map (
            O => \N__49600\,
            I => \N__49070\
        );

    \I__11794\ : SRMux
    port map (
            O => \N__49599\,
            I => \N__49070\
        );

    \I__11793\ : SRMux
    port map (
            O => \N__49598\,
            I => \N__49070\
        );

    \I__11792\ : SRMux
    port map (
            O => \N__49597\,
            I => \N__49070\
        );

    \I__11791\ : SRMux
    port map (
            O => \N__49596\,
            I => \N__49070\
        );

    \I__11790\ : SRMux
    port map (
            O => \N__49595\,
            I => \N__49070\
        );

    \I__11789\ : SRMux
    port map (
            O => \N__49594\,
            I => \N__49070\
        );

    \I__11788\ : SRMux
    port map (
            O => \N__49593\,
            I => \N__49070\
        );

    \I__11787\ : SRMux
    port map (
            O => \N__49592\,
            I => \N__49070\
        );

    \I__11786\ : SRMux
    port map (
            O => \N__49591\,
            I => \N__49070\
        );

    \I__11785\ : SRMux
    port map (
            O => \N__49590\,
            I => \N__49070\
        );

    \I__11784\ : SRMux
    port map (
            O => \N__49589\,
            I => \N__49070\
        );

    \I__11783\ : SRMux
    port map (
            O => \N__49588\,
            I => \N__49070\
        );

    \I__11782\ : SRMux
    port map (
            O => \N__49587\,
            I => \N__49070\
        );

    \I__11781\ : SRMux
    port map (
            O => \N__49586\,
            I => \N__49070\
        );

    \I__11780\ : SRMux
    port map (
            O => \N__49585\,
            I => \N__49070\
        );

    \I__11779\ : SRMux
    port map (
            O => \N__49584\,
            I => \N__49070\
        );

    \I__11778\ : SRMux
    port map (
            O => \N__49583\,
            I => \N__49070\
        );

    \I__11777\ : SRMux
    port map (
            O => \N__49582\,
            I => \N__49070\
        );

    \I__11776\ : SRMux
    port map (
            O => \N__49581\,
            I => \N__49070\
        );

    \I__11775\ : SRMux
    port map (
            O => \N__49580\,
            I => \N__49070\
        );

    \I__11774\ : SRMux
    port map (
            O => \N__49579\,
            I => \N__49070\
        );

    \I__11773\ : SRMux
    port map (
            O => \N__49578\,
            I => \N__49070\
        );

    \I__11772\ : SRMux
    port map (
            O => \N__49577\,
            I => \N__49070\
        );

    \I__11771\ : SRMux
    port map (
            O => \N__49576\,
            I => \N__49070\
        );

    \I__11770\ : SRMux
    port map (
            O => \N__49575\,
            I => \N__49070\
        );

    \I__11769\ : SRMux
    port map (
            O => \N__49574\,
            I => \N__49070\
        );

    \I__11768\ : SRMux
    port map (
            O => \N__49573\,
            I => \N__49070\
        );

    \I__11767\ : SRMux
    port map (
            O => \N__49572\,
            I => \N__49070\
        );

    \I__11766\ : SRMux
    port map (
            O => \N__49571\,
            I => \N__49070\
        );

    \I__11765\ : SRMux
    port map (
            O => \N__49570\,
            I => \N__49070\
        );

    \I__11764\ : SRMux
    port map (
            O => \N__49569\,
            I => \N__49070\
        );

    \I__11763\ : SRMux
    port map (
            O => \N__49568\,
            I => \N__49070\
        );

    \I__11762\ : SRMux
    port map (
            O => \N__49567\,
            I => \N__49070\
        );

    \I__11761\ : SRMux
    port map (
            O => \N__49566\,
            I => \N__49070\
        );

    \I__11760\ : SRMux
    port map (
            O => \N__49565\,
            I => \N__49070\
        );

    \I__11759\ : SRMux
    port map (
            O => \N__49564\,
            I => \N__49070\
        );

    \I__11758\ : SRMux
    port map (
            O => \N__49563\,
            I => \N__49070\
        );

    \I__11757\ : SRMux
    port map (
            O => \N__49562\,
            I => \N__49070\
        );

    \I__11756\ : SRMux
    port map (
            O => \N__49561\,
            I => \N__49070\
        );

    \I__11755\ : SRMux
    port map (
            O => \N__49560\,
            I => \N__49070\
        );

    \I__11754\ : SRMux
    port map (
            O => \N__49559\,
            I => \N__49070\
        );

    \I__11753\ : SRMux
    port map (
            O => \N__49558\,
            I => \N__49070\
        );

    \I__11752\ : SRMux
    port map (
            O => \N__49557\,
            I => \N__49070\
        );

    \I__11751\ : SRMux
    port map (
            O => \N__49556\,
            I => \N__49070\
        );

    \I__11750\ : SRMux
    port map (
            O => \N__49555\,
            I => \N__49070\
        );

    \I__11749\ : SRMux
    port map (
            O => \N__49554\,
            I => \N__49070\
        );

    \I__11748\ : SRMux
    port map (
            O => \N__49553\,
            I => \N__49070\
        );

    \I__11747\ : SRMux
    port map (
            O => \N__49552\,
            I => \N__49070\
        );

    \I__11746\ : SRMux
    port map (
            O => \N__49551\,
            I => \N__49070\
        );

    \I__11745\ : SRMux
    port map (
            O => \N__49550\,
            I => \N__49070\
        );

    \I__11744\ : SRMux
    port map (
            O => \N__49549\,
            I => \N__49070\
        );

    \I__11743\ : SRMux
    port map (
            O => \N__49548\,
            I => \N__49070\
        );

    \I__11742\ : SRMux
    port map (
            O => \N__49547\,
            I => \N__49070\
        );

    \I__11741\ : SRMux
    port map (
            O => \N__49546\,
            I => \N__49070\
        );

    \I__11740\ : SRMux
    port map (
            O => \N__49545\,
            I => \N__49070\
        );

    \I__11739\ : SRMux
    port map (
            O => \N__49544\,
            I => \N__49070\
        );

    \I__11738\ : SRMux
    port map (
            O => \N__49543\,
            I => \N__49070\
        );

    \I__11737\ : SRMux
    port map (
            O => \N__49542\,
            I => \N__49070\
        );

    \I__11736\ : SRMux
    port map (
            O => \N__49541\,
            I => \N__49070\
        );

    \I__11735\ : SRMux
    port map (
            O => \N__49540\,
            I => \N__49070\
        );

    \I__11734\ : SRMux
    port map (
            O => \N__49539\,
            I => \N__49070\
        );

    \I__11733\ : SRMux
    port map (
            O => \N__49538\,
            I => \N__49070\
        );

    \I__11732\ : SRMux
    port map (
            O => \N__49537\,
            I => \N__49070\
        );

    \I__11731\ : SRMux
    port map (
            O => \N__49536\,
            I => \N__49070\
        );

    \I__11730\ : SRMux
    port map (
            O => \N__49535\,
            I => \N__49070\
        );

    \I__11729\ : SRMux
    port map (
            O => \N__49534\,
            I => \N__49070\
        );

    \I__11728\ : SRMux
    port map (
            O => \N__49533\,
            I => \N__49070\
        );

    \I__11727\ : SRMux
    port map (
            O => \N__49532\,
            I => \N__49070\
        );

    \I__11726\ : SRMux
    port map (
            O => \N__49531\,
            I => \N__49070\
        );

    \I__11725\ : SRMux
    port map (
            O => \N__49530\,
            I => \N__49070\
        );

    \I__11724\ : SRMux
    port map (
            O => \N__49529\,
            I => \N__49070\
        );

    \I__11723\ : SRMux
    port map (
            O => \N__49528\,
            I => \N__49070\
        );

    \I__11722\ : SRMux
    port map (
            O => \N__49527\,
            I => \N__49070\
        );

    \I__11721\ : SRMux
    port map (
            O => \N__49526\,
            I => \N__49070\
        );

    \I__11720\ : SRMux
    port map (
            O => \N__49525\,
            I => \N__49070\
        );

    \I__11719\ : SRMux
    port map (
            O => \N__49524\,
            I => \N__49070\
        );

    \I__11718\ : SRMux
    port map (
            O => \N__49523\,
            I => \N__49070\
        );

    \I__11717\ : SRMux
    port map (
            O => \N__49522\,
            I => \N__49070\
        );

    \I__11716\ : SRMux
    port map (
            O => \N__49521\,
            I => \N__49070\
        );

    \I__11715\ : SRMux
    port map (
            O => \N__49520\,
            I => \N__49070\
        );

    \I__11714\ : SRMux
    port map (
            O => \N__49519\,
            I => \N__49070\
        );

    \I__11713\ : SRMux
    port map (
            O => \N__49518\,
            I => \N__49070\
        );

    \I__11712\ : SRMux
    port map (
            O => \N__49517\,
            I => \N__49070\
        );

    \I__11711\ : SRMux
    port map (
            O => \N__49516\,
            I => \N__49070\
        );

    \I__11710\ : SRMux
    port map (
            O => \N__49515\,
            I => \N__49070\
        );

    \I__11709\ : SRMux
    port map (
            O => \N__49514\,
            I => \N__49070\
        );

    \I__11708\ : SRMux
    port map (
            O => \N__49513\,
            I => \N__49070\
        );

    \I__11707\ : SRMux
    port map (
            O => \N__49512\,
            I => \N__49070\
        );

    \I__11706\ : SRMux
    port map (
            O => \N__49511\,
            I => \N__49070\
        );

    \I__11705\ : SRMux
    port map (
            O => \N__49510\,
            I => \N__49070\
        );

    \I__11704\ : SRMux
    port map (
            O => \N__49509\,
            I => \N__49070\
        );

    \I__11703\ : SRMux
    port map (
            O => \N__49508\,
            I => \N__49070\
        );

    \I__11702\ : SRMux
    port map (
            O => \N__49507\,
            I => \N__49070\
        );

    \I__11701\ : SRMux
    port map (
            O => \N__49506\,
            I => \N__49070\
        );

    \I__11700\ : SRMux
    port map (
            O => \N__49505\,
            I => \N__49070\
        );

    \I__11699\ : SRMux
    port map (
            O => \N__49504\,
            I => \N__49070\
        );

    \I__11698\ : SRMux
    port map (
            O => \N__49503\,
            I => \N__49070\
        );

    \I__11697\ : SRMux
    port map (
            O => \N__49502\,
            I => \N__49070\
        );

    \I__11696\ : SRMux
    port map (
            O => \N__49501\,
            I => \N__49070\
        );

    \I__11695\ : SRMux
    port map (
            O => \N__49500\,
            I => \N__49070\
        );

    \I__11694\ : SRMux
    port map (
            O => \N__49499\,
            I => \N__49070\
        );

    \I__11693\ : SRMux
    port map (
            O => \N__49498\,
            I => \N__49070\
        );

    \I__11692\ : Glb2LocalMux
    port map (
            O => \N__49495\,
            I => \N__49070\
        );

    \I__11691\ : Glb2LocalMux
    port map (
            O => \N__49492\,
            I => \N__49070\
        );

    \I__11690\ : Glb2LocalMux
    port map (
            O => \N__49489\,
            I => \N__49070\
        );

    \I__11689\ : Glb2LocalMux
    port map (
            O => \N__49486\,
            I => \N__49070\
        );

    \I__11688\ : Glb2LocalMux
    port map (
            O => \N__49483\,
            I => \N__49070\
        );

    \I__11687\ : Glb2LocalMux
    port map (
            O => \N__49480\,
            I => \N__49070\
        );

    \I__11686\ : Glb2LocalMux
    port map (
            O => \N__49477\,
            I => \N__49070\
        );

    \I__11685\ : Glb2LocalMux
    port map (
            O => \N__49474\,
            I => \N__49070\
        );

    \I__11684\ : Glb2LocalMux
    port map (
            O => \N__49471\,
            I => \N__49070\
        );

    \I__11683\ : Glb2LocalMux
    port map (
            O => \N__49468\,
            I => \N__49070\
        );

    \I__11682\ : Glb2LocalMux
    port map (
            O => \N__49465\,
            I => \N__49070\
        );

    \I__11681\ : Glb2LocalMux
    port map (
            O => \N__49462\,
            I => \N__49070\
        );

    \I__11680\ : Glb2LocalMux
    port map (
            O => \N__49459\,
            I => \N__49070\
        );

    \I__11679\ : Glb2LocalMux
    port map (
            O => \N__49456\,
            I => \N__49070\
        );

    \I__11678\ : Glb2LocalMux
    port map (
            O => \N__49453\,
            I => \N__49070\
        );

    \I__11677\ : Glb2LocalMux
    port map (
            O => \N__49450\,
            I => \N__49070\
        );

    \I__11676\ : Glb2LocalMux
    port map (
            O => \N__49447\,
            I => \N__49070\
        );

    \I__11675\ : Glb2LocalMux
    port map (
            O => \N__49444\,
            I => \N__49070\
        );

    \I__11674\ : Glb2LocalMux
    port map (
            O => \N__49441\,
            I => \N__49070\
        );

    \I__11673\ : Glb2LocalMux
    port map (
            O => \N__49438\,
            I => \N__49070\
        );

    \I__11672\ : Glb2LocalMux
    port map (
            O => \N__49435\,
            I => \N__49070\
        );

    \I__11671\ : Glb2LocalMux
    port map (
            O => \N__49432\,
            I => \N__49070\
        );

    \I__11670\ : Glb2LocalMux
    port map (
            O => \N__49429\,
            I => \N__49070\
        );

    \I__11669\ : Glb2LocalMux
    port map (
            O => \N__49426\,
            I => \N__49070\
        );

    \I__11668\ : Glb2LocalMux
    port map (
            O => \N__49423\,
            I => \N__49070\
        );

    \I__11667\ : Glb2LocalMux
    port map (
            O => \N__49420\,
            I => \N__49070\
        );

    \I__11666\ : Glb2LocalMux
    port map (
            O => \N__49417\,
            I => \N__49070\
        );

    \I__11665\ : Glb2LocalMux
    port map (
            O => \N__49414\,
            I => \N__49070\
        );

    \I__11664\ : Glb2LocalMux
    port map (
            O => \N__49411\,
            I => \N__49070\
        );

    \I__11663\ : Glb2LocalMux
    port map (
            O => \N__49408\,
            I => \N__49070\
        );

    \I__11662\ : Glb2LocalMux
    port map (
            O => \N__49405\,
            I => \N__49070\
        );

    \I__11661\ : Glb2LocalMux
    port map (
            O => \N__49402\,
            I => \N__49070\
        );

    \I__11660\ : Glb2LocalMux
    port map (
            O => \N__49399\,
            I => \N__49070\
        );

    \I__11659\ : GlobalMux
    port map (
            O => \N__49070\,
            I => \N__49067\
        );

    \I__11658\ : gio2CtrlBuf
    port map (
            O => \N__49067\,
            I => reset_system_g
        );

    \I__11657\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49061\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__49061\,
            I => \N__49058\
        );

    \I__11655\ : Span4Mux_v
    port map (
            O => \N__49058\,
            I => \N__49055\
        );

    \I__11654\ : Span4Mux_h
    port map (
            O => \N__49055\,
            I => \N__49052\
        );

    \I__11653\ : Span4Mux_h
    port map (
            O => \N__49052\,
            I => \N__49049\
        );

    \I__11652\ : Odrv4
    port map (
            O => \N__49049\,
            I => \pid_front.state_ns_0\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49046\,
            I => \N__49043\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__49043\,
            I => \N__49039\
        );

    \I__11649\ : InMux
    port map (
            O => \N__49042\,
            I => \N__49035\
        );

    \I__11648\ : Span4Mux_v
    port map (
            O => \N__49039\,
            I => \N__49030\
        );

    \I__11647\ : InMux
    port map (
            O => \N__49038\,
            I => \N__49027\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__49035\,
            I => \N__49019\
        );

    \I__11645\ : IoInMux
    port map (
            O => \N__49034\,
            I => \N__49016\
        );

    \I__11644\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49011\
        );

    \I__11643\ : Span4Mux_h
    port map (
            O => \N__49030\,
            I => \N__49005\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__49027\,
            I => \N__49005\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49026\,
            I => \N__49000\
        );

    \I__11640\ : InMux
    port map (
            O => \N__49025\,
            I => \N__49000\
        );

    \I__11639\ : InMux
    port map (
            O => \N__49024\,
            I => \N__48997\
        );

    \I__11638\ : InMux
    port map (
            O => \N__49023\,
            I => \N__48994\
        );

    \I__11637\ : InMux
    port map (
            O => \N__49022\,
            I => \N__48990\
        );

    \I__11636\ : Span4Mux_v
    port map (
            O => \N__49019\,
            I => \N__48984\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__49016\,
            I => \N__48981\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49015\,
            I => \N__48974\
        );

    \I__11633\ : InMux
    port map (
            O => \N__49014\,
            I => \N__48971\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__49011\,
            I => \N__48962\
        );

    \I__11631\ : InMux
    port map (
            O => \N__49010\,
            I => \N__48958\
        );

    \I__11630\ : Span4Mux_v
    port map (
            O => \N__49005\,
            I => \N__48953\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48946\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__48997\,
            I => \N__48946\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__48994\,
            I => \N__48946\
        );

    \I__11626\ : InMux
    port map (
            O => \N__48993\,
            I => \N__48943\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__48990\,
            I => \N__48940\
        );

    \I__11624\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48933\
        );

    \I__11623\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48933\
        );

    \I__11622\ : InMux
    port map (
            O => \N__48987\,
            I => \N__48933\
        );

    \I__11621\ : Span4Mux_v
    port map (
            O => \N__48984\,
            I => \N__48930\
        );

    \I__11620\ : Span4Mux_s1_v
    port map (
            O => \N__48981\,
            I => \N__48927\
        );

    \I__11619\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48922\
        );

    \I__11618\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48922\
        );

    \I__11617\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48919\
        );

    \I__11616\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48916\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__48974\,
            I => \N__48911\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__48971\,
            I => \N__48911\
        );

    \I__11613\ : InMux
    port map (
            O => \N__48970\,
            I => \N__48905\
        );

    \I__11612\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48905\
        );

    \I__11611\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48900\
        );

    \I__11610\ : InMux
    port map (
            O => \N__48967\,
            I => \N__48900\
        );

    \I__11609\ : InMux
    port map (
            O => \N__48966\,
            I => \N__48895\
        );

    \I__11608\ : InMux
    port map (
            O => \N__48965\,
            I => \N__48895\
        );

    \I__11607\ : Span4Mux_h
    port map (
            O => \N__48962\,
            I => \N__48892\
        );

    \I__11606\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48889\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__48958\,
            I => \N__48886\
        );

    \I__11604\ : InMux
    port map (
            O => \N__48957\,
            I => \N__48881\
        );

    \I__11603\ : InMux
    port map (
            O => \N__48956\,
            I => \N__48881\
        );

    \I__11602\ : Span4Mux_h
    port map (
            O => \N__48953\,
            I => \N__48876\
        );

    \I__11601\ : Span4Mux_v
    port map (
            O => \N__48946\,
            I => \N__48876\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__48943\,
            I => \N__48869\
        );

    \I__11599\ : Span4Mux_v
    port map (
            O => \N__48940\,
            I => \N__48869\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__48933\,
            I => \N__48869\
        );

    \I__11597\ : Span4Mux_v
    port map (
            O => \N__48930\,
            I => \N__48864\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__48927\,
            I => \N__48864\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__48922\,
            I => \N__48859\
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__48919\,
            I => \N__48859\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__48916\,
            I => \N__48856\
        );

    \I__11592\ : Span4Mux_v
    port map (
            O => \N__48911\,
            I => \N__48853\
        );

    \I__11591\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48850\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__48905\,
            I => \N__48839\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__48900\,
            I => \N__48839\
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__48895\,
            I => \N__48839\
        );

    \I__11587\ : Sp12to4
    port map (
            O => \N__48892\,
            I => \N__48839\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__48889\,
            I => \N__48839\
        );

    \I__11585\ : Span4Mux_v
    port map (
            O => \N__48886\,
            I => \N__48836\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__48881\,
            I => \N__48831\
        );

    \I__11583\ : Span4Mux_v
    port map (
            O => \N__48876\,
            I => \N__48831\
        );

    \I__11582\ : Span4Mux_v
    port map (
            O => \N__48869\,
            I => \N__48826\
        );

    \I__11581\ : Span4Mux_h
    port map (
            O => \N__48864\,
            I => \N__48826\
        );

    \I__11580\ : Span4Mux_v
    port map (
            O => \N__48859\,
            I => \N__48823\
        );

    \I__11579\ : Span4Mux_h
    port map (
            O => \N__48856\,
            I => \N__48820\
        );

    \I__11578\ : Span4Mux_v
    port map (
            O => \N__48853\,
            I => \N__48817\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__48850\,
            I => \N__48812\
        );

    \I__11576\ : Span12Mux_v
    port map (
            O => \N__48839\,
            I => \N__48812\
        );

    \I__11575\ : Span4Mux_v
    port map (
            O => \N__48836\,
            I => \N__48805\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__48831\,
            I => \N__48805\
        );

    \I__11573\ : Span4Mux_h
    port map (
            O => \N__48826\,
            I => \N__48805\
        );

    \I__11572\ : Odrv4
    port map (
            O => \N__48823\,
            I => reset_system
        );

    \I__11571\ : Odrv4
    port map (
            O => \N__48820\,
            I => reset_system
        );

    \I__11570\ : Odrv4
    port map (
            O => \N__48817\,
            I => reset_system
        );

    \I__11569\ : Odrv12
    port map (
            O => \N__48812\,
            I => reset_system
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__48805\,
            I => reset_system
        );

    \I__11567\ : InMux
    port map (
            O => \N__48794\,
            I => \N__48791\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__48791\,
            I => \N__48788\
        );

    \I__11565\ : Odrv12
    port map (
            O => \N__48788\,
            I => \pid_front.O_5\
        );

    \I__11564\ : InMux
    port map (
            O => \N__48785\,
            I => \N__48781\
        );

    \I__11563\ : InMux
    port map (
            O => \N__48784\,
            I => \N__48778\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48775\
        );

    \I__11561\ : LocalMux
    port map (
            O => \N__48778\,
            I => \N__48771\
        );

    \I__11560\ : Span12Mux_v
    port map (
            O => \N__48775\,
            I => \N__48768\
        );

    \I__11559\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48765\
        );

    \I__11558\ : Span4Mux_h
    port map (
            O => \N__48771\,
            I => \N__48762\
        );

    \I__11557\ : Odrv12
    port map (
            O => \N__48768\,
            I => \pid_front.error_p_regZ0Z_1\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__48765\,
            I => \pid_front.error_p_regZ0Z_1\
        );

    \I__11555\ : Odrv4
    port map (
            O => \N__48762\,
            I => \pid_front.error_p_regZ0Z_1\
        );

    \I__11554\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48752\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__48752\,
            I => \N__48749\
        );

    \I__11552\ : Span4Mux_h
    port map (
            O => \N__48749\,
            I => \N__48746\
        );

    \I__11551\ : Odrv4
    port map (
            O => \N__48746\,
            I => \pid_front.O_13\
        );

    \I__11550\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48740\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__48740\,
            I => \N__48735\
        );

    \I__11548\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48732\
        );

    \I__11547\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48729\
        );

    \I__11546\ : Span12Mux_h
    port map (
            O => \N__48735\,
            I => \N__48724\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__48732\,
            I => \N__48724\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__48729\,
            I => \pid_front.error_p_regZ0Z_9\
        );

    \I__11543\ : Odrv12
    port map (
            O => \N__48724\,
            I => \pid_front.error_p_regZ0Z_9\
        );

    \I__11542\ : InMux
    port map (
            O => \N__48719\,
            I => \N__48716\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__48716\,
            I => \N__48713\
        );

    \I__11540\ : Odrv4
    port map (
            O => \N__48713\,
            I => \pid_front.O_6\
        );

    \I__11539\ : InMux
    port map (
            O => \N__48710\,
            I => \N__48706\
        );

    \I__11538\ : InMux
    port map (
            O => \N__48709\,
            I => \N__48703\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__48706\,
            I => \N__48699\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__48703\,
            I => \N__48696\
        );

    \I__11535\ : InMux
    port map (
            O => \N__48702\,
            I => \N__48693\
        );

    \I__11534\ : Span4Mux_h
    port map (
            O => \N__48699\,
            I => \N__48690\
        );

    \I__11533\ : Odrv12
    port map (
            O => \N__48696\,
            I => \pid_front.error_p_regZ0Z_2\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__48693\,
            I => \pid_front.error_p_regZ0Z_2\
        );

    \I__11531\ : Odrv4
    port map (
            O => \N__48690\,
            I => \pid_front.error_p_regZ0Z_2\
        );

    \I__11530\ : InMux
    port map (
            O => \N__48683\,
            I => \N__48680\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__48680\,
            I => \N__48677\
        );

    \I__11528\ : Span4Mux_v
    port map (
            O => \N__48677\,
            I => \N__48674\
        );

    \I__11527\ : Odrv4
    port map (
            O => \N__48674\,
            I => \pid_front.O_9\
        );

    \I__11526\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48668\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__48668\,
            I => \N__48664\
        );

    \I__11524\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48661\
        );

    \I__11523\ : Span4Mux_v
    port map (
            O => \N__48664\,
            I => \N__48657\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__48661\,
            I => \N__48654\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48660\,
            I => \N__48651\
        );

    \I__11520\ : Span4Mux_h
    port map (
            O => \N__48657\,
            I => \N__48648\
        );

    \I__11519\ : Span12Mux_h
    port map (
            O => \N__48654\,
            I => \N__48645\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__48651\,
            I => \pid_front.error_p_regZ0Z_5\
        );

    \I__11517\ : Odrv4
    port map (
            O => \N__48648\,
            I => \pid_front.error_p_regZ0Z_5\
        );

    \I__11516\ : Odrv12
    port map (
            O => \N__48645\,
            I => \pid_front.error_p_regZ0Z_5\
        );

    \I__11515\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48635\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__48635\,
            I => \N__48632\
        );

    \I__11513\ : Span4Mux_v
    port map (
            O => \N__48632\,
            I => \N__48629\
        );

    \I__11512\ : Odrv4
    port map (
            O => \N__48629\,
            I => \pid_front.O_8\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48626\,
            I => \N__48622\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48619\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__48622\,
            I => \N__48616\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__48619\,
            I => \N__48613\
        );

    \I__11507\ : Span4Mux_v
    port map (
            O => \N__48616\,
            I => \N__48609\
        );

    \I__11506\ : Span4Mux_h
    port map (
            O => \N__48613\,
            I => \N__48606\
        );

    \I__11505\ : InMux
    port map (
            O => \N__48612\,
            I => \N__48603\
        );

    \I__11504\ : Span4Mux_h
    port map (
            O => \N__48609\,
            I => \N__48600\
        );

    \I__11503\ : Span4Mux_h
    port map (
            O => \N__48606\,
            I => \N__48597\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__48603\,
            I => \pid_front.error_p_regZ0Z_4\
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__48600\,
            I => \pid_front.error_p_regZ0Z_4\
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__48597\,
            I => \pid_front.error_p_regZ0Z_4\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48590\,
            I => \N__48587\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__48587\,
            I => \N__48584\
        );

    \I__11497\ : Span4Mux_h
    port map (
            O => \N__48584\,
            I => \N__48581\
        );

    \I__11496\ : Odrv4
    port map (
            O => \N__48581\,
            I => \pid_front.un1_pid_prereg_cry_17_THRU_CO\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48578\,
            I => \pid_front.un1_pid_prereg_cry_17\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48572\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__48572\,
            I => \N__48569\
        );

    \I__11492\ : Span4Mux_v
    port map (
            O => \N__48569\,
            I => \N__48566\
        );

    \I__11491\ : Odrv4
    port map (
            O => \N__48566\,
            I => \pid_front.un1_pid_prereg_cry_18_THRU_CO\
        );

    \I__11490\ : InMux
    port map (
            O => \N__48563\,
            I => \pid_front.un1_pid_prereg_cry_18\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48560\,
            I => \N__48557\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__48557\,
            I => \N__48554\
        );

    \I__11487\ : Span4Mux_v
    port map (
            O => \N__48554\,
            I => \N__48551\
        );

    \I__11486\ : Odrv4
    port map (
            O => \N__48551\,
            I => \pid_front.un1_pid_prereg_cry_19_THRU_CO\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48548\,
            I => \pid_front.un1_pid_prereg_cry_19\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48545\,
            I => \pid_front.un1_pid_prereg_cry_20\
        );

    \I__11483\ : CascadeMux
    port map (
            O => \N__48542\,
            I => \N__48539\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48539\,
            I => \N__48530\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48538\,
            I => \N__48530\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48527\
        );

    \I__11479\ : CascadeMux
    port map (
            O => \N__48536\,
            I => \N__48524\
        );

    \I__11478\ : CascadeMux
    port map (
            O => \N__48535\,
            I => \N__48521\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48530\,
            I => \N__48516\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__48527\,
            I => \N__48516\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48513\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48521\,
            I => \N__48510\
        );

    \I__11473\ : Span4Mux_h
    port map (
            O => \N__48516\,
            I => \N__48507\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__48513\,
            I => \N__48504\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48501\
        );

    \I__11470\ : Span4Mux_v
    port map (
            O => \N__48507\,
            I => \N__48498\
        );

    \I__11469\ : Span4Mux_h
    port map (
            O => \N__48504\,
            I => \N__48493\
        );

    \I__11468\ : Span4Mux_v
    port map (
            O => \N__48501\,
            I => \N__48493\
        );

    \I__11467\ : Span4Mux_h
    port map (
            O => \N__48498\,
            I => \N__48490\
        );

    \I__11466\ : Span4Mux_h
    port map (
            O => \N__48493\,
            I => \N__48487\
        );

    \I__11465\ : Odrv4
    port map (
            O => \N__48490\,
            I => \pid_front.pid_preregZ0Z_21\
        );

    \I__11464\ : Odrv4
    port map (
            O => \N__48487\,
            I => \pid_front.pid_preregZ0Z_21\
        );

    \I__11463\ : CEMux
    port map (
            O => \N__48482\,
            I => \N__48478\
        );

    \I__11462\ : CEMux
    port map (
            O => \N__48481\,
            I => \N__48475\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__48478\,
            I => \N__48472\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__48475\,
            I => \N__48469\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__48472\,
            I => \N__48466\
        );

    \I__11458\ : Span4Mux_v
    port map (
            O => \N__48469\,
            I => \N__48463\
        );

    \I__11457\ : Span4Mux_h
    port map (
            O => \N__48466\,
            I => \N__48458\
        );

    \I__11456\ : Span4Mux_h
    port map (
            O => \N__48463\,
            I => \N__48458\
        );

    \I__11455\ : Odrv4
    port map (
            O => \N__48458\,
            I => \pid_front.state_0_0\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48455\,
            I => \N__48452\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__48452\,
            I => \N__48449\
        );

    \I__11452\ : Span4Mux_h
    port map (
            O => \N__48449\,
            I => \N__48445\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48448\,
            I => \N__48442\
        );

    \I__11450\ : Span4Mux_v
    port map (
            O => \N__48445\,
            I => \N__48437\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__48442\,
            I => \N__48437\
        );

    \I__11448\ : Span4Mux_h
    port map (
            O => \N__48437\,
            I => \N__48430\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48427\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48423\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48434\,
            I => \N__48420\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48433\,
            I => \N__48417\
        );

    \I__11443\ : Span4Mux_h
    port map (
            O => \N__48430\,
            I => \N__48412\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48412\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48409\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48423\,
            I => \N__48403\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__48420\,
            I => \N__48403\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__48417\,
            I => \N__48400\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__48412\,
            I => \N__48397\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48409\,
            I => \N__48394\
        );

    \I__11435\ : CascadeMux
    port map (
            O => \N__48408\,
            I => \N__48391\
        );

    \I__11434\ : Span12Mux_s10_h
    port map (
            O => \N__48403\,
            I => \N__48386\
        );

    \I__11433\ : Span12Mux_s11_v
    port map (
            O => \N__48400\,
            I => \N__48386\
        );

    \I__11432\ : Span4Mux_v
    port map (
            O => \N__48397\,
            I => \N__48381\
        );

    \I__11431\ : Span4Mux_v
    port map (
            O => \N__48394\,
            I => \N__48381\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48378\
        );

    \I__11429\ : Odrv12
    port map (
            O => \N__48386\,
            I => uart_drone_data_6
        );

    \I__11428\ : Odrv4
    port map (
            O => \N__48381\,
            I => uart_drone_data_6
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__48378\,
            I => uart_drone_data_6
        );

    \I__11426\ : CascadeMux
    port map (
            O => \N__48371\,
            I => \N__48367\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48370\,
            I => \N__48362\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48367\,
            I => \N__48362\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__48362\,
            I => \drone_H_disp_front_14\
        );

    \I__11422\ : CEMux
    port map (
            O => \N__48359\,
            I => \N__48356\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__48356\,
            I => \N__48351\
        );

    \I__11420\ : CEMux
    port map (
            O => \N__48355\,
            I => \N__48348\
        );

    \I__11419\ : CEMux
    port map (
            O => \N__48354\,
            I => \N__48345\
        );

    \I__11418\ : Span4Mux_v
    port map (
            O => \N__48351\,
            I => \N__48341\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48348\,
            I => \N__48336\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__48345\,
            I => \N__48336\
        );

    \I__11415\ : CEMux
    port map (
            O => \N__48344\,
            I => \N__48333\
        );

    \I__11414\ : Span4Mux_h
    port map (
            O => \N__48341\,
            I => \N__48326\
        );

    \I__11413\ : Span4Mux_v
    port map (
            O => \N__48336\,
            I => \N__48326\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48333\,
            I => \N__48326\
        );

    \I__11411\ : Span4Mux_h
    port map (
            O => \N__48326\,
            I => \N__48323\
        );

    \I__11410\ : Span4Mux_v
    port map (
            O => \N__48323\,
            I => \N__48320\
        );

    \I__11409\ : Span4Mux_v
    port map (
            O => \N__48320\,
            I => \N__48317\
        );

    \I__11408\ : Odrv4
    port map (
            O => \N__48317\,
            I => \dron_frame_decoder_1.N_723_0\
        );

    \I__11407\ : IoInMux
    port map (
            O => \N__48314\,
            I => \N__48311\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48311\,
            I => \GB_BUFFER_reset_system_g_THRU_CO\
        );

    \I__11405\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48305\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48305\,
            I => \N__48302\
        );

    \I__11403\ : Span12Mux_h
    port map (
            O => \N__48302\,
            I => \N__48299\
        );

    \I__11402\ : Odrv12
    port map (
            O => \N__48299\,
            I => \pid_side.O_0_4\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48296\,
            I => \N__48293\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48290\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__48290\,
            I => \N__48286\
        );

    \I__11398\ : InMux
    port map (
            O => \N__48289\,
            I => \N__48283\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__48286\,
            I => \pid_side.error_p_regZ0Z_0\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__48283\,
            I => \pid_side.error_p_regZ0Z_0\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48275\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48272\
        );

    \I__11393\ : Span12Mux_h
    port map (
            O => \N__48272\,
            I => \N__48269\
        );

    \I__11392\ : Odrv12
    port map (
            O => \N__48269\,
            I => \pid_side.O_0_5\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48263\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48263\,
            I => \N__48260\
        );

    \I__11389\ : Span4Mux_h
    port map (
            O => \N__48260\,
            I => \N__48257\
        );

    \I__11388\ : Odrv4
    port map (
            O => \N__48257\,
            I => \pid_front.un1_pid_prereg_cry_9_THRU_CO\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48254\,
            I => \pid_front.un1_pid_prereg_cry_9\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48251\,
            I => \N__48248\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__48248\,
            I => \N__48245\
        );

    \I__11384\ : Span4Mux_h
    port map (
            O => \N__48245\,
            I => \N__48242\
        );

    \I__11383\ : Odrv4
    port map (
            O => \N__48242\,
            I => \pid_front.un1_pid_prereg_cry_10_THRU_CO\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48239\,
            I => \pid_front.un1_pid_prereg_cry_10\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48226\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48223\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48234\,
            I => \N__48220\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48217\
        );

    \I__11377\ : CascadeMux
    port map (
            O => \N__48232\,
            I => \N__48214\
        );

    \I__11376\ : CascadeMux
    port map (
            O => \N__48231\,
            I => \N__48211\
        );

    \I__11375\ : InMux
    port map (
            O => \N__48230\,
            I => \N__48203\
        );

    \I__11374\ : InMux
    port map (
            O => \N__48229\,
            I => \N__48200\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48226\,
            I => \N__48194\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48194\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__48220\,
            I => \N__48185\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__48217\,
            I => \N__48185\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48180\
        );

    \I__11368\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48180\
        );

    \I__11367\ : CascadeMux
    port map (
            O => \N__48210\,
            I => \N__48177\
        );

    \I__11366\ : CascadeMux
    port map (
            O => \N__48209\,
            I => \N__48170\
        );

    \I__11365\ : CascadeMux
    port map (
            O => \N__48208\,
            I => \N__48166\
        );

    \I__11364\ : CascadeMux
    port map (
            O => \N__48207\,
            I => \N__48162\
        );

    \I__11363\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48158\
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__48203\,
            I => \N__48155\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__48200\,
            I => \N__48152\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48149\
        );

    \I__11359\ : Span4Mux_v
    port map (
            O => \N__48194\,
            I => \N__48146\
        );

    \I__11358\ : InMux
    port map (
            O => \N__48193\,
            I => \N__48143\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48140\
        );

    \I__11356\ : CascadeMux
    port map (
            O => \N__48191\,
            I => \N__48137\
        );

    \I__11355\ : CascadeMux
    port map (
            O => \N__48190\,
            I => \N__48133\
        );

    \I__11354\ : Span4Mux_v
    port map (
            O => \N__48185\,
            I => \N__48125\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48180\,
            I => \N__48122\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48119\
        );

    \I__11351\ : CascadeMux
    port map (
            O => \N__48176\,
            I => \N__48116\
        );

    \I__11350\ : CascadeMux
    port map (
            O => \N__48175\,
            I => \N__48113\
        );

    \I__11349\ : CascadeMux
    port map (
            O => \N__48174\,
            I => \N__48110\
        );

    \I__11348\ : CascadeMux
    port map (
            O => \N__48173\,
            I => \N__48107\
        );

    \I__11347\ : InMux
    port map (
            O => \N__48170\,
            I => \N__48099\
        );

    \I__11346\ : InMux
    port map (
            O => \N__48169\,
            I => \N__48099\
        );

    \I__11345\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48096\
        );

    \I__11344\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48091\
        );

    \I__11343\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48091\
        );

    \I__11342\ : CascadeMux
    port map (
            O => \N__48161\,
            I => \N__48088\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__48158\,
            I => \N__48081\
        );

    \I__11340\ : Span4Mux_v
    port map (
            O => \N__48155\,
            I => \N__48074\
        );

    \I__11339\ : Span4Mux_v
    port map (
            O => \N__48152\,
            I => \N__48074\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__48149\,
            I => \N__48074\
        );

    \I__11337\ : Span4Mux_v
    port map (
            O => \N__48146\,
            I => \N__48069\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__48143\,
            I => \N__48069\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__48140\,
            I => \N__48066\
        );

    \I__11334\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48059\
        );

    \I__11333\ : InMux
    port map (
            O => \N__48136\,
            I => \N__48059\
        );

    \I__11332\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48059\
        );

    \I__11331\ : CascadeMux
    port map (
            O => \N__48132\,
            I => \N__48056\
        );

    \I__11330\ : CascadeMux
    port map (
            O => \N__48131\,
            I => \N__48053\
        );

    \I__11329\ : CascadeMux
    port map (
            O => \N__48130\,
            I => \N__48050\
        );

    \I__11328\ : CascadeMux
    port map (
            O => \N__48129\,
            I => \N__48047\
        );

    \I__11327\ : CascadeMux
    port map (
            O => \N__48128\,
            I => \N__48044\
        );

    \I__11326\ : Span4Mux_h
    port map (
            O => \N__48125\,
            I => \N__48037\
        );

    \I__11325\ : Span4Mux_v
    port map (
            O => \N__48122\,
            I => \N__48032\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__48119\,
            I => \N__48032\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48116\,
            I => \N__48023\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48113\,
            I => \N__48023\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48110\,
            I => \N__48023\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48023\
        );

    \I__11319\ : CascadeMux
    port map (
            O => \N__48106\,
            I => \N__48020\
        );

    \I__11318\ : CascadeMux
    port map (
            O => \N__48105\,
            I => \N__48017\
        );

    \I__11317\ : CascadeMux
    port map (
            O => \N__48104\,
            I => \N__48014\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__48011\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__48096\,
            I => \N__48006\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48091\,
            I => \N__48006\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48003\
        );

    \I__11312\ : CascadeMux
    port map (
            O => \N__48087\,
            I => \N__48000\
        );

    \I__11311\ : CascadeMux
    port map (
            O => \N__48086\,
            I => \N__47997\
        );

    \I__11310\ : CascadeMux
    port map (
            O => \N__48085\,
            I => \N__47994\
        );

    \I__11309\ : CascadeMux
    port map (
            O => \N__48084\,
            I => \N__47991\
        );

    \I__11308\ : Span4Mux_v
    port map (
            O => \N__48081\,
            I => \N__47982\
        );

    \I__11307\ : Span4Mux_v
    port map (
            O => \N__48074\,
            I => \N__47982\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__48069\,
            I => \N__47982\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__48066\,
            I => \N__47979\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__48059\,
            I => \N__47976\
        );

    \I__11303\ : InMux
    port map (
            O => \N__48056\,
            I => \N__47971\
        );

    \I__11302\ : InMux
    port map (
            O => \N__48053\,
            I => \N__47971\
        );

    \I__11301\ : InMux
    port map (
            O => \N__48050\,
            I => \N__47966\
        );

    \I__11300\ : InMux
    port map (
            O => \N__48047\,
            I => \N__47966\
        );

    \I__11299\ : InMux
    port map (
            O => \N__48044\,
            I => \N__47963\
        );

    \I__11298\ : CascadeMux
    port map (
            O => \N__48043\,
            I => \N__47960\
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__48042\,
            I => \N__47957\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__48041\,
            I => \N__47954\
        );

    \I__11295\ : CascadeMux
    port map (
            O => \N__48040\,
            I => \N__47951\
        );

    \I__11294\ : Span4Mux_h
    port map (
            O => \N__48037\,
            I => \N__47948\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__48032\,
            I => \N__47943\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__48023\,
            I => \N__47943\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48020\,
            I => \N__47936\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48017\,
            I => \N__47936\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48014\,
            I => \N__47936\
        );

    \I__11288\ : Span4Mux_v
    port map (
            O => \N__48011\,
            I => \N__47929\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__48006\,
            I => \N__47929\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__48003\,
            I => \N__47929\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48000\,
            I => \N__47926\
        );

    \I__11284\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47923\
        );

    \I__11283\ : InMux
    port map (
            O => \N__47994\,
            I => \N__47918\
        );

    \I__11282\ : InMux
    port map (
            O => \N__47991\,
            I => \N__47918\
        );

    \I__11281\ : InMux
    port map (
            O => \N__47990\,
            I => \N__47915\
        );

    \I__11280\ : InMux
    port map (
            O => \N__47989\,
            I => \N__47912\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__47982\,
            I => \N__47907\
        );

    \I__11278\ : Span4Mux_h
    port map (
            O => \N__47979\,
            I => \N__47907\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__47976\,
            I => \N__47900\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__47971\,
            I => \N__47900\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__47966\,
            I => \N__47900\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__47963\,
            I => \N__47897\
        );

    \I__11273\ : InMux
    port map (
            O => \N__47960\,
            I => \N__47894\
        );

    \I__11272\ : InMux
    port map (
            O => \N__47957\,
            I => \N__47891\
        );

    \I__11271\ : InMux
    port map (
            O => \N__47954\,
            I => \N__47886\
        );

    \I__11270\ : InMux
    port map (
            O => \N__47951\,
            I => \N__47886\
        );

    \I__11269\ : Span4Mux_v
    port map (
            O => \N__47948\,
            I => \N__47880\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__47943\,
            I => \N__47875\
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__47936\,
            I => \N__47875\
        );

    \I__11266\ : Span4Mux_v
    port map (
            O => \N__47929\,
            I => \N__47872\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__47926\,
            I => \N__47865\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__47923\,
            I => \N__47865\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__47918\,
            I => \N__47865\
        );

    \I__11262\ : LocalMux
    port map (
            O => \N__47915\,
            I => \N__47860\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__47912\,
            I => \N__47860\
        );

    \I__11260\ : Span4Mux_h
    port map (
            O => \N__47907\,
            I => \N__47853\
        );

    \I__11259\ : Span4Mux_v
    port map (
            O => \N__47900\,
            I => \N__47853\
        );

    \I__11258\ : Span4Mux_v
    port map (
            O => \N__47897\,
            I => \N__47853\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__47894\,
            I => \N__47846\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__47891\,
            I => \N__47846\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__47886\,
            I => \N__47846\
        );

    \I__11254\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47843\
        );

    \I__11253\ : CascadeMux
    port map (
            O => \N__47884\,
            I => \N__47839\
        );

    \I__11252\ : CascadeMux
    port map (
            O => \N__47883\,
            I => \N__47836\
        );

    \I__11251\ : Span4Mux_v
    port map (
            O => \N__47880\,
            I => \N__47833\
        );

    \I__11250\ : Span4Mux_v
    port map (
            O => \N__47875\,
            I => \N__47830\
        );

    \I__11249\ : Span4Mux_h
    port map (
            O => \N__47872\,
            I => \N__47823\
        );

    \I__11248\ : Span4Mux_v
    port map (
            O => \N__47865\,
            I => \N__47823\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__47860\,
            I => \N__47823\
        );

    \I__11246\ : Span4Mux_h
    port map (
            O => \N__47853\,
            I => \N__47816\
        );

    \I__11245\ : Span4Mux_v
    port map (
            O => \N__47846\,
            I => \N__47816\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__47843\,
            I => \N__47816\
        );

    \I__11243\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47809\
        );

    \I__11242\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47809\
        );

    \I__11241\ : InMux
    port map (
            O => \N__47836\,
            I => \N__47809\
        );

    \I__11240\ : Odrv4
    port map (
            O => \N__47833\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11239\ : Odrv4
    port map (
            O => \N__47830\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11238\ : Odrv4
    port map (
            O => \N__47823\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11237\ : Odrv4
    port map (
            O => \N__47816\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47809\,
            I => \CONSTANT_ONE_NET\
        );

    \I__11235\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47795\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__47795\,
            I => \N__47792\
        );

    \I__11233\ : Span4Mux_h
    port map (
            O => \N__47792\,
            I => \N__47789\
        );

    \I__11232\ : Odrv4
    port map (
            O => \N__47789\,
            I => \pid_front.un1_pid_prereg_cry_11_THRU_CO\
        );

    \I__11231\ : InMux
    port map (
            O => \N__47786\,
            I => \pid_front.un1_pid_prereg_cry_11\
        );

    \I__11230\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47780\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__47780\,
            I => \N__47777\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__47777\,
            I => \N__47774\
        );

    \I__11227\ : Odrv4
    port map (
            O => \N__47774\,
            I => \pid_front.un1_pid_prereg_cry_12_THRU_CO\
        );

    \I__11226\ : InMux
    port map (
            O => \N__47771\,
            I => \pid_front.un1_pid_prereg_cry_12\
        );

    \I__11225\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47765\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__47765\,
            I => \N__47762\
        );

    \I__11223\ : Span4Mux_v
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__11222\ : Odrv4
    port map (
            O => \N__47759\,
            I => \pid_front.un1_pid_prereg_cry_13_THRU_CO\
        );

    \I__11221\ : InMux
    port map (
            O => \N__47756\,
            I => \pid_front.un1_pid_prereg_cry_13\
        );

    \I__11220\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47750\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__47750\,
            I => \N__47747\
        );

    \I__11218\ : Odrv4
    port map (
            O => \N__47747\,
            I => \pid_front.un1_pid_prereg_cry_14_THRU_CO\
        );

    \I__11217\ : InMux
    port map (
            O => \N__47744\,
            I => \pid_front.un1_pid_prereg_cry_14\
        );

    \I__11216\ : InMux
    port map (
            O => \N__47741\,
            I => \N__47738\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__47738\,
            I => \N__47735\
        );

    \I__11214\ : Odrv4
    port map (
            O => \N__47735\,
            I => \pid_front.un1_pid_prereg_cry_15_THRU_CO\
        );

    \I__11213\ : InMux
    port map (
            O => \N__47732\,
            I => \pid_front.un1_pid_prereg_cry_15\
        );

    \I__11212\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47726\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__47726\,
            I => \N__47723\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__47723\,
            I => \N__47720\
        );

    \I__11209\ : Odrv4
    port map (
            O => \N__47720\,
            I => \pid_front.un1_pid_prereg_cry_16_THRU_CO\
        );

    \I__11208\ : InMux
    port map (
            O => \N__47717\,
            I => \bfn_18_24_0_\
        );

    \I__11207\ : SRMux
    port map (
            O => \N__47714\,
            I => \N__47705\
        );

    \I__11206\ : SRMux
    port map (
            O => \N__47713\,
            I => \N__47705\
        );

    \I__11205\ : SRMux
    port map (
            O => \N__47712\,
            I => \N__47705\
        );

    \I__11204\ : GlobalMux
    port map (
            O => \N__47705\,
            I => \N__47702\
        );

    \I__11203\ : gio2CtrlBuf
    port map (
            O => \N__47702\,
            I => \ppm_encoder_1.N_661_g\
        );

    \I__11202\ : CascadeMux
    port map (
            O => \N__47699\,
            I => \N__47696\
        );

    \I__11201\ : InMux
    port map (
            O => \N__47696\,
            I => \N__47693\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__47693\,
            I => \N__47690\
        );

    \I__11199\ : Span4Mux_h
    port map (
            O => \N__47690\,
            I => \N__47687\
        );

    \I__11198\ : Odrv4
    port map (
            O => \N__47687\,
            I => \pid_front.un1_pid_prereg_cry_1_THRU_CO\
        );

    \I__11197\ : InMux
    port map (
            O => \N__47684\,
            I => \pid_front.un1_pid_prereg_cry_1\
        );

    \I__11196\ : CascadeMux
    port map (
            O => \N__47681\,
            I => \N__47678\
        );

    \I__11195\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47675\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47672\
        );

    \I__11193\ : Span4Mux_h
    port map (
            O => \N__47672\,
            I => \N__47669\
        );

    \I__11192\ : Odrv4
    port map (
            O => \N__47669\,
            I => \pid_front.un1_pid_prereg_cry_2_THRU_CO\
        );

    \I__11191\ : InMux
    port map (
            O => \N__47666\,
            I => \pid_front.un1_pid_prereg_cry_2\
        );

    \I__11190\ : CascadeMux
    port map (
            O => \N__47663\,
            I => \N__47660\
        );

    \I__11189\ : InMux
    port map (
            O => \N__47660\,
            I => \N__47657\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__47657\,
            I => \N__47654\
        );

    \I__11187\ : Span4Mux_v
    port map (
            O => \N__47654\,
            I => \N__47651\
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__47651\,
            I => \pid_front.un1_pid_prereg_cry_3_THRU_CO\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47648\,
            I => \pid_front.un1_pid_prereg_cry_3\
        );

    \I__11184\ : CascadeMux
    port map (
            O => \N__47645\,
            I => \N__47642\
        );

    \I__11183\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47639\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47639\,
            I => \N__47636\
        );

    \I__11181\ : Span4Mux_h
    port map (
            O => \N__47636\,
            I => \N__47633\
        );

    \I__11180\ : Odrv4
    port map (
            O => \N__47633\,
            I => \pid_front.un1_pid_prereg_cry_4_THRU_CO\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47630\,
            I => \pid_front.un1_pid_prereg_cry_4\
        );

    \I__11178\ : InMux
    port map (
            O => \N__47627\,
            I => \N__47624\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__47624\,
            I => \N__47621\
        );

    \I__11176\ : Span4Mux_h
    port map (
            O => \N__47621\,
            I => \N__47618\
        );

    \I__11175\ : Odrv4
    port map (
            O => \N__47618\,
            I => \pid_front.un1_pid_prereg_cry_5_THRU_CO\
        );

    \I__11174\ : InMux
    port map (
            O => \N__47615\,
            I => \pid_front.un1_pid_prereg_cry_5\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47609\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__47609\,
            I => \N__47606\
        );

    \I__11171\ : Odrv12
    port map (
            O => \N__47606\,
            I => \pid_front.un1_pid_prereg_cry_6_THRU_CO\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47603\,
            I => \pid_front.un1_pid_prereg_cry_6\
        );

    \I__11169\ : InMux
    port map (
            O => \N__47600\,
            I => \N__47597\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__47597\,
            I => \pid_front.un1_pid_prereg_cry_7_THRU_CO\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47594\,
            I => \pid_front.un1_pid_prereg_cry_7\
        );

    \I__11166\ : InMux
    port map (
            O => \N__47591\,
            I => \N__47588\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__47588\,
            I => \N__47585\
        );

    \I__11164\ : Span4Mux_h
    port map (
            O => \N__47585\,
            I => \N__47582\
        );

    \I__11163\ : Odrv4
    port map (
            O => \N__47582\,
            I => \pid_front.un1_pid_prereg_cry_8_THRU_CO\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47579\,
            I => \bfn_18_23_0_\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47576\,
            I => \N__47571\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47575\,
            I => \N__47568\
        );

    \I__11159\ : InMux
    port map (
            O => \N__47574\,
            I => \N__47565\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__47571\,
            I => \N__47562\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47568\,
            I => \N__47559\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__47565\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47562\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__47559\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__11153\ : InMux
    port map (
            O => \N__47552\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47549\,
            I => \N__47544\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47548\,
            I => \N__47541\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47547\,
            I => \N__47538\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47544\,
            I => \N__47535\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__47541\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47538\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__11146\ : Odrv4
    port map (
            O => \N__47535\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__11145\ : InMux
    port map (
            O => \N__47528\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47520\
        );

    \I__11143\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47517\
        );

    \I__11142\ : InMux
    port map (
            O => \N__47523\,
            I => \N__47514\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__47520\,
            I => \N__47511\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__47517\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__47514\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__11138\ : Odrv4
    port map (
            O => \N__47511\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47504\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47498\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__47498\,
            I => \N__47493\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47497\,
            I => \N__47490\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47487\
        );

    \I__11132\ : Span4Mux_v
    port map (
            O => \N__47493\,
            I => \N__47484\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__47490\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47487\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__11129\ : Odrv4
    port map (
            O => \N__47484\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__11128\ : InMux
    port map (
            O => \N__47477\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__11127\ : CascadeMux
    port map (
            O => \N__47474\,
            I => \N__47471\
        );

    \I__11126\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47468\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__47468\,
            I => \N__47463\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47467\,
            I => \N__47460\
        );

    \I__11123\ : InMux
    port map (
            O => \N__47466\,
            I => \N__47457\
        );

    \I__11122\ : Span4Mux_v
    port map (
            O => \N__47463\,
            I => \N__47454\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47460\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47457\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__11119\ : Odrv4
    port map (
            O => \N__47454\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47447\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47444\,
            I => \N__47439\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47443\,
            I => \N__47436\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47442\,
            I => \N__47433\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__47439\,
            I => \N__47430\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__47436\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47433\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__11111\ : Odrv12
    port map (
            O => \N__47430\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47423\,
            I => \bfn_18_21_0_\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47420\,
            I => \N__47415\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47419\,
            I => \N__47412\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47409\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47415\,
            I => \N__47406\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47412\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47409\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__11103\ : Odrv12
    port map (
            O => \N__47406\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47399\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47396\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__47393\,
            I => \N__47388\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47392\,
            I => \N__47385\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47382\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47388\,
            I => \N__47379\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__47385\,
            I => \N__47376\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__47382\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47379\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__11093\ : Odrv12
    port map (
            O => \N__47376\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47369\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47366\,
            I => \N__47360\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47355\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47355\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47352\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47360\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__47355\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47352\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47345\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__11083\ : InMux
    port map (
            O => \N__47342\,
            I => \N__47337\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47341\,
            I => \N__47334\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47331\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47337\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47334\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__47331\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47324\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47321\,
            I => \N__47316\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47313\
        );

    \I__11074\ : InMux
    port map (
            O => \N__47319\,
            I => \N__47310\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__47316\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47313\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__47310\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__11070\ : InMux
    port map (
            O => \N__47303\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47295\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47299\,
            I => \N__47292\
        );

    \I__11067\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47289\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47295\,
            I => \N__47286\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__47292\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__47289\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__11063\ : Odrv12
    port map (
            O => \N__47286\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47279\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47272\
        );

    \I__11060\ : CascadeMux
    port map (
            O => \N__47275\,
            I => \N__47268\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__47272\,
            I => \N__47265\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47262\
        );

    \I__11057\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47259\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__47265\,
            I => \N__47256\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47262\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47259\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__11053\ : Odrv4
    port map (
            O => \N__47256\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__11052\ : InMux
    port map (
            O => \N__47249\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__11051\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47241\
        );

    \I__11050\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47238\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47235\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47232\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__47238\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__47235\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__11045\ : Odrv4
    port map (
            O => \N__47232\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__11044\ : InMux
    port map (
            O => \N__47225\,
            I => \bfn_18_20_0_\
        );

    \I__11043\ : InMux
    port map (
            O => \N__47222\,
            I => \N__47215\
        );

    \I__11042\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47215\
        );

    \I__11041\ : InMux
    port map (
            O => \N__47220\,
            I => \N__47212\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47215\,
            I => \N__47209\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47212\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__11038\ : Odrv4
    port map (
            O => \N__47209\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__11037\ : InMux
    port map (
            O => \N__47204\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__11036\ : CascadeMux
    port map (
            O => \N__47201\,
            I => \N__47198\
        );

    \I__11035\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47191\
        );

    \I__11034\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47191\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47188\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47185\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47188\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__11030\ : Odrv4
    port map (
            O => \N__47185\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__11029\ : InMux
    port map (
            O => \N__47180\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__11028\ : InMux
    port map (
            O => \N__47177\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47167\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47167\
        );

    \I__11025\ : CascadeMux
    port map (
            O => \N__47172\,
            I => \N__47164\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47167\,
            I => \N__47160\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47155\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47155\
        );

    \I__11021\ : Odrv4
    port map (
            O => \N__47160\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__47155\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47147\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__47147\,
            I => \N__47144\
        );

    \I__11017\ : Odrv12
    port map (
            O => \N__47144\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__11016\ : CascadeMux
    port map (
            O => \N__47141\,
            I => \N__47138\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47135\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__47135\,
            I => \N__47132\
        );

    \I__11013\ : Span4Mux_v
    port map (
            O => \N__47132\,
            I => \N__47129\
        );

    \I__11012\ : Odrv4
    port map (
            O => \N__47129\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47123\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__47123\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__11009\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47117\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__47117\,
            I => \N__47114\
        );

    \I__11007\ : Span4Mux_v
    port map (
            O => \N__47114\,
            I => \N__47111\
        );

    \I__11006\ : Odrv4
    port map (
            O => \N__47111\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__11005\ : CascadeMux
    port map (
            O => \N__47108\,
            I => \N__47105\
        );

    \I__11004\ : InMux
    port map (
            O => \N__47105\,
            I => \N__47102\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__47099\
        );

    \I__11002\ : Span4Mux_v
    port map (
            O => \N__47099\,
            I => \N__47096\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__47096\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47093\,
            I => \N__47090\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__47090\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47087\,
            I => \N__47081\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47086\,
            I => \N__47081\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47081\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47078\,
            I => \N__47075\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__47075\,
            I => \N__47072\
        );

    \I__10993\ : Odrv12
    port map (
            O => \N__47072\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__10992\ : CascadeMux
    port map (
            O => \N__47069\,
            I => \N__47066\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47066\,
            I => \N__47063\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__47063\,
            I => \N__47060\
        );

    \I__10989\ : Span4Mux_h
    port map (
            O => \N__47060\,
            I => \N__47057\
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__47057\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47054\,
            I => \N__47051\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__47051\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__10985\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47045\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47045\,
            I => \N__47042\
        );

    \I__10983\ : Span4Mux_v
    port map (
            O => \N__47042\,
            I => \N__47039\
        );

    \I__10982\ : Odrv4
    port map (
            O => \N__47039\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__10981\ : CascadeMux
    port map (
            O => \N__47036\,
            I => \N__47033\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47030\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47027\
        );

    \I__10978\ : Span4Mux_v
    port map (
            O => \N__47027\,
            I => \N__47024\
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__47024\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__10976\ : InMux
    port map (
            O => \N__47021\,
            I => \N__47018\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__47018\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__10974\ : InMux
    port map (
            O => \N__47015\,
            I => \N__47011\
        );

    \I__10973\ : CascadeMux
    port map (
            O => \N__47014\,
            I => \N__47008\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__47011\,
            I => \N__47005\
        );

    \I__10971\ : InMux
    port map (
            O => \N__47008\,
            I => \N__47002\
        );

    \I__10970\ : Odrv4
    port map (
            O => \N__47005\,
            I => \ppm_encoder_1.N_1818_i\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47002\,
            I => \ppm_encoder_1.N_1818_i\
        );

    \I__10968\ : InMux
    port map (
            O => \N__46997\,
            I => \N__46992\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46989\
        );

    \I__10966\ : InMux
    port map (
            O => \N__46995\,
            I => \N__46986\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__46992\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__46989\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__46986\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__10962\ : InMux
    port map (
            O => \N__46979\,
            I => \N__46973\
        );

    \I__10961\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46966\
        );

    \I__10960\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46966\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46966\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__46973\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__46966\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__10956\ : InMux
    port map (
            O => \N__46961\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__10955\ : CascadeMux
    port map (
            O => \N__46958\,
            I => \N__46955\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46955\,
            I => \N__46950\
        );

    \I__10953\ : CascadeMux
    port map (
            O => \N__46954\,
            I => \N__46947\
        );

    \I__10952\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46943\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46940\
        );

    \I__10950\ : InMux
    port map (
            O => \N__46947\,
            I => \N__46935\
        );

    \I__10949\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46935\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46943\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__10947\ : Odrv4
    port map (
            O => \N__46940\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__46935\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46925\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__46925\,
            I => \N__46922\
        );

    \I__10943\ : Odrv12
    port map (
            O => \N__46922\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__10942\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46916\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__46916\,
            I => \N__46913\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__46913\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__10939\ : InMux
    port map (
            O => \N__46910\,
            I => \N__46907\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__46907\,
            I => \N__46904\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__46904\,
            I => \N__46901\
        );

    \I__10936\ : Odrv4
    port map (
            O => \N__46901\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46895\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46892\
        );

    \I__10933\ : Odrv12
    port map (
            O => \N__46892\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46889\,
            I => \N__46886\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46886\,
            I => \N__46883\
        );

    \I__10930\ : Odrv12
    port map (
            O => \N__46883\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4\
        );

    \I__10929\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46877\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__46877\,
            I => \N__46874\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__46874\,
            I => \N__46871\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__46871\,
            I => \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46868\,
            I => \N__46864\
        );

    \I__10924\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46861\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46858\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46853\
        );

    \I__10921\ : Span4Mux_v
    port map (
            O => \N__46858\,
            I => \N__46853\
        );

    \I__10920\ : Odrv4
    port map (
            O => \N__46853\,
            I => side_order_4
        );

    \I__10919\ : CascadeMux
    port map (
            O => \N__46850\,
            I => \N__46847\
        );

    \I__10918\ : InMux
    port map (
            O => \N__46847\,
            I => \N__46844\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__46844\,
            I => \N__46841\
        );

    \I__10916\ : Span4Mux_h
    port map (
            O => \N__46841\,
            I => \N__46838\
        );

    \I__10915\ : Odrv4
    port map (
            O => \N__46838\,
            I => \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\
        );

    \I__10914\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46832\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__46832\,
            I => \N__46828\
        );

    \I__10912\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46825\
        );

    \I__10911\ : Span4Mux_v
    port map (
            O => \N__46828\,
            I => \N__46820\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46820\
        );

    \I__10909\ : Span4Mux_h
    port map (
            O => \N__46820\,
            I => \N__46817\
        );

    \I__10908\ : Odrv4
    port map (
            O => \N__46817\,
            I => front_order_4
        );

    \I__10907\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46808\
        );

    \I__10906\ : CascadeMux
    port map (
            O => \N__46813\,
            I => \N__46802\
        );

    \I__10905\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46799\
        );

    \I__10904\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46796\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46792\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46807\,
            I => \N__46789\
        );

    \I__10901\ : InMux
    port map (
            O => \N__46806\,
            I => \N__46783\
        );

    \I__10900\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46779\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46776\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46799\,
            I => \N__46771\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__46796\,
            I => \N__46771\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46768\
        );

    \I__10895\ : Span4Mux_v
    port map (
            O => \N__46792\,
            I => \N__46760\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46789\,
            I => \N__46760\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46755\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46755\
        );

    \I__10891\ : InMux
    port map (
            O => \N__46786\,
            I => \N__46749\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46746\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46742\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__46779\,
            I => \N__46733\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46733\
        );

    \I__10886\ : Span4Mux_v
    port map (
            O => \N__46771\,
            I => \N__46733\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__46768\,
            I => \N__46733\
        );

    \I__10884\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46730\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46725\
        );

    \I__10882\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46725\
        );

    \I__10881\ : Span4Mux_h
    port map (
            O => \N__46760\,
            I => \N__46720\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__46755\,
            I => \N__46720\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46713\
        );

    \I__10878\ : InMux
    port map (
            O => \N__46753\,
            I => \N__46713\
        );

    \I__10877\ : InMux
    port map (
            O => \N__46752\,
            I => \N__46713\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46708\
        );

    \I__10875\ : Span4Mux_v
    port map (
            O => \N__46746\,
            I => \N__46708\
        );

    \I__10874\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46705\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46700\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__46733\,
            I => \N__46700\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46730\,
            I => \N__46693\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46725\,
            I => \N__46693\
        );

    \I__10869\ : Sp12to4
    port map (
            O => \N__46720\,
            I => \N__46693\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46690\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__46708\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__46705\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__46700\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10864\ : Odrv12
    port map (
            O => \N__46693\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10863\ : Odrv12
    port map (
            O => \N__46690\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__10862\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46670\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46670\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46677\,
            I => \N__46670\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__46670\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46667\,
            I => \N__46659\
        );

    \I__10857\ : CascadeMux
    port map (
            O => \N__46666\,
            I => \N__46656\
        );

    \I__10856\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46652\
        );

    \I__10855\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46649\
        );

    \I__10854\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46646\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__46662\,
            I => \N__46639\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46659\,
            I => \N__46636\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46656\,
            I => \N__46633\
        );

    \I__10850\ : CascadeMux
    port map (
            O => \N__46655\,
            I => \N__46627\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46652\,
            I => \N__46624\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46649\,
            I => \N__46619\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__46646\,
            I => \N__46619\
        );

    \I__10846\ : CascadeMux
    port map (
            O => \N__46645\,
            I => \N__46616\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46644\,
            I => \N__46613\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46643\,
            I => \N__46610\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46605\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46605\
        );

    \I__10841\ : Span4Mux_v
    port map (
            O => \N__46636\,
            I => \N__46602\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46633\,
            I => \N__46598\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46632\,
            I => \N__46593\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46631\,
            I => \N__46593\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46630\,
            I => \N__46590\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46586\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__46624\,
            I => \N__46577\
        );

    \I__10834\ : Span4Mux_v
    port map (
            O => \N__46619\,
            I => \N__46577\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46616\,
            I => \N__46574\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46613\,
            I => \N__46567\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46567\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46567\
        );

    \I__10829\ : Span4Mux_h
    port map (
            O => \N__46602\,
            I => \N__46564\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46561\
        );

    \I__10827\ : Span4Mux_v
    port map (
            O => \N__46598\,
            I => \N__46554\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__46593\,
            I => \N__46554\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__46590\,
            I => \N__46554\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46551\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46586\,
            I => \N__46548\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46585\,
            I => \N__46545\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46542\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46539\
        );

    \I__10819\ : CascadeMux
    port map (
            O => \N__46582\,
            I => \N__46535\
        );

    \I__10818\ : Span4Mux_h
    port map (
            O => \N__46577\,
            I => \N__46532\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46574\,
            I => \N__46523\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__46567\,
            I => \N__46523\
        );

    \I__10815\ : Span4Mux_h
    port map (
            O => \N__46564\,
            I => \N__46523\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46523\
        );

    \I__10813\ : Span4Mux_v
    port map (
            O => \N__46554\,
            I => \N__46518\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46518\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__46548\,
            I => \N__46509\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46545\,
            I => \N__46509\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46542\,
            I => \N__46509\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__46539\,
            I => \N__46509\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46538\,
            I => \N__46506\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46535\,
            I => \N__46503\
        );

    \I__10805\ : Span4Mux_v
    port map (
            O => \N__46532\,
            I => \N__46500\
        );

    \I__10804\ : Span4Mux_v
    port map (
            O => \N__46523\,
            I => \N__46497\
        );

    \I__10803\ : Span4Mux_h
    port map (
            O => \N__46518\,
            I => \N__46490\
        );

    \I__10802\ : Span4Mux_v
    port map (
            O => \N__46509\,
            I => \N__46490\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46506\,
            I => \N__46490\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__46503\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__46500\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__10798\ : Odrv4
    port map (
            O => \N__46497\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__10797\ : Odrv4
    port map (
            O => \N__46490\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__10796\ : CascadeMux
    port map (
            O => \N__46481\,
            I => \ppm_encoder_1.N_290_cascade_\
        );

    \I__10795\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46469\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46469\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46469\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__46469\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46463\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46463\,
            I => \N__46460\
        );

    \I__10789\ : Odrv12
    port map (
            O => \N__46460\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46457\,
            I => \N__46454\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46454\,
            I => \N__46451\
        );

    \I__10786\ : Span4Mux_v
    port map (
            O => \N__46451\,
            I => \N__46448\
        );

    \I__10785\ : Span4Mux_h
    port map (
            O => \N__46448\,
            I => \N__46445\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__46445\,
            I => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46442\,
            I => \N__46439\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46439\,
            I => \N__46435\
        );

    \I__10781\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46432\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__46435\,
            I => \N__46429\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__46432\,
            I => \N__46426\
        );

    \I__10778\ : Span4Mux_h
    port map (
            O => \N__46429\,
            I => \N__46423\
        );

    \I__10777\ : Span4Mux_v
    port map (
            O => \N__46426\,
            I => \N__46420\
        );

    \I__10776\ : Odrv4
    port map (
            O => \N__46423\,
            I => throttle_order_4
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__46420\,
            I => throttle_order_4
        );

    \I__10774\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46410\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46405\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46405\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__46410\,
            I => \N__46402\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46405\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__46402\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__10768\ : CascadeMux
    port map (
            O => \N__46397\,
            I => \N__46391\
        );

    \I__10767\ : CascadeMux
    port map (
            O => \N__46396\,
            I => \N__46383\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__46395\,
            I => \N__46380\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__46394\,
            I => \N__46377\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46371\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__46390\,
            I => \N__46368\
        );

    \I__10762\ : CascadeMux
    port map (
            O => \N__46389\,
            I => \N__46362\
        );

    \I__10761\ : CascadeMux
    port map (
            O => \N__46388\,
            I => \N__46359\
        );

    \I__10760\ : CascadeMux
    port map (
            O => \N__46387\,
            I => \N__46356\
        );

    \I__10759\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46351\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46351\
        );

    \I__10757\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46348\
        );

    \I__10756\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46343\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46343\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__46375\,
            I => \N__46337\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__46374\,
            I => \N__46334\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__46371\,
            I => \N__46329\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46368\,
            I => \N__46325\
        );

    \I__10750\ : CascadeMux
    port map (
            O => \N__46367\,
            I => \N__46322\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46366\,
            I => \N__46312\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46365\,
            I => \N__46312\
        );

    \I__10747\ : InMux
    port map (
            O => \N__46362\,
            I => \N__46312\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46312\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46301\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__46351\,
            I => \N__46294\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46348\,
            I => \N__46294\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__46343\,
            I => \N__46294\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46279\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46279\
        );

    \I__10739\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46279\
        );

    \I__10738\ : InMux
    port map (
            O => \N__46337\,
            I => \N__46279\
        );

    \I__10737\ : InMux
    port map (
            O => \N__46334\,
            I => \N__46279\
        );

    \I__10736\ : InMux
    port map (
            O => \N__46333\,
            I => \N__46279\
        );

    \I__10735\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46279\
        );

    \I__10734\ : Span4Mux_h
    port map (
            O => \N__46329\,
            I => \N__46276\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46328\,
            I => \N__46273\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__46325\,
            I => \N__46270\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46265\
        );

    \I__10730\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46265\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46312\,
            I => \N__46262\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46311\,
            I => \N__46257\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46257\
        );

    \I__10726\ : CascadeMux
    port map (
            O => \N__46309\,
            I => \N__46252\
        );

    \I__10725\ : CascadeMux
    port map (
            O => \N__46308\,
            I => \N__46249\
        );

    \I__10724\ : CascadeMux
    port map (
            O => \N__46307\,
            I => \N__46245\
        );

    \I__10723\ : CascadeMux
    port map (
            O => \N__46306\,
            I => \N__46239\
        );

    \I__10722\ : CascadeMux
    port map (
            O => \N__46305\,
            I => \N__46236\
        );

    \I__10721\ : CascadeMux
    port map (
            O => \N__46304\,
            I => \N__46233\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__46301\,
            I => \N__46230\
        );

    \I__10719\ : Span4Mux_v
    port map (
            O => \N__46294\,
            I => \N__46221\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__46279\,
            I => \N__46221\
        );

    \I__10717\ : Span4Mux_v
    port map (
            O => \N__46276\,
            I => \N__46221\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46273\,
            I => \N__46221\
        );

    \I__10715\ : Span4Mux_h
    port map (
            O => \N__46270\,
            I => \N__46212\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__46265\,
            I => \N__46212\
        );

    \I__10713\ : Span4Mux_h
    port map (
            O => \N__46262\,
            I => \N__46212\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__46257\,
            I => \N__46212\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46209\
        );

    \I__10710\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46200\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46200\
        );

    \I__10708\ : InMux
    port map (
            O => \N__46249\,
            I => \N__46200\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46200\
        );

    \I__10706\ : InMux
    port map (
            O => \N__46245\,
            I => \N__46195\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46195\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46243\,
            I => \N__46176\
        );

    \I__10703\ : InMux
    port map (
            O => \N__46242\,
            I => \N__46176\
        );

    \I__10702\ : InMux
    port map (
            O => \N__46239\,
            I => \N__46176\
        );

    \I__10701\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46176\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46176\
        );

    \I__10699\ : Span4Mux_v
    port map (
            O => \N__46230\,
            I => \N__46171\
        );

    \I__10698\ : Span4Mux_v
    port map (
            O => \N__46221\,
            I => \N__46171\
        );

    \I__10697\ : Span4Mux_v
    port map (
            O => \N__46212\,
            I => \N__46161\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__46209\,
            I => \N__46161\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__46200\,
            I => \N__46161\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__46195\,
            I => \N__46161\
        );

    \I__10693\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46158\
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__46193\,
            I => \N__46152\
        );

    \I__10691\ : CascadeMux
    port map (
            O => \N__46192\,
            I => \N__46148\
        );

    \I__10690\ : CascadeMux
    port map (
            O => \N__46191\,
            I => \N__46145\
        );

    \I__10689\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46141\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__46189\,
            I => \N__46137\
        );

    \I__10687\ : CascadeMux
    port map (
            O => \N__46188\,
            I => \N__46134\
        );

    \I__10686\ : CascadeMux
    port map (
            O => \N__46187\,
            I => \N__46131\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__46176\,
            I => \N__46128\
        );

    \I__10684\ : Span4Mux_h
    port map (
            O => \N__46171\,
            I => \N__46125\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__46170\,
            I => \N__46122\
        );

    \I__10682\ : Span4Mux_v
    port map (
            O => \N__46161\,
            I => \N__46119\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__46158\,
            I => \N__46116\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46157\,
            I => \N__46113\
        );

    \I__10679\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46106\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46106\
        );

    \I__10677\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46106\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46097\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46097\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46145\,
            I => \N__46097\
        );

    \I__10673\ : InMux
    port map (
            O => \N__46144\,
            I => \N__46097\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46141\,
            I => \N__46094\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46140\,
            I => \N__46085\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46085\
        );

    \I__10669\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46085\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46131\,
            I => \N__46085\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__46128\,
            I => \N__46082\
        );

    \I__10666\ : Span4Mux_h
    port map (
            O => \N__46125\,
            I => \N__46079\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46122\,
            I => \N__46076\
        );

    \I__10664\ : Span4Mux_h
    port map (
            O => \N__46119\,
            I => \N__46069\
        );

    \I__10663\ : Span4Mux_v
    port map (
            O => \N__46116\,
            I => \N__46069\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__46113\,
            I => \N__46069\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__46106\,
            I => \N__46062\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46097\,
            I => \N__46062\
        );

    \I__10659\ : Sp12to4
    port map (
            O => \N__46094\,
            I => \N__46062\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__46085\,
            I => \N__46059\
        );

    \I__10657\ : Span4Mux_h
    port map (
            O => \N__46082\,
            I => \N__46054\
        );

    \I__10656\ : Span4Mux_v
    port map (
            O => \N__46079\,
            I => \N__46054\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46076\,
            I => \N__46049\
        );

    \I__10654\ : Span4Mux_v
    port map (
            O => \N__46069\,
            I => \N__46049\
        );

    \I__10653\ : Span12Mux_v
    port map (
            O => \N__46062\,
            I => \N__46046\
        );

    \I__10652\ : Span4Mux_v
    port map (
            O => \N__46059\,
            I => \N__46041\
        );

    \I__10651\ : Span4Mux_v
    port map (
            O => \N__46054\,
            I => \N__46041\
        );

    \I__10650\ : Span4Mux_v
    port map (
            O => \N__46049\,
            I => \N__46038\
        );

    \I__10649\ : Odrv12
    port map (
            O => \N__46046\,
            I => pid_altitude_dv
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__46041\,
            I => pid_altitude_dv
        );

    \I__10647\ : Odrv4
    port map (
            O => \N__46038\,
            I => pid_altitude_dv
        );

    \I__10646\ : InMux
    port map (
            O => \N__46031\,
            I => \N__46027\
        );

    \I__10645\ : CascadeMux
    port map (
            O => \N__46030\,
            I => \N__46023\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__46020\
        );

    \I__10643\ : InMux
    port map (
            O => \N__46026\,
            I => \N__46017\
        );

    \I__10642\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46014\
        );

    \I__10641\ : Span4Mux_v
    port map (
            O => \N__46020\,
            I => \N__46011\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__46008\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46014\,
            I => side_order_0
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__46011\,
            I => side_order_0
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__46008\,
            I => side_order_0
        );

    \I__10636\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45998\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__45998\,
            I => \N__45994\
        );

    \I__10634\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45990\
        );

    \I__10633\ : Span4Mux_v
    port map (
            O => \N__45994\,
            I => \N__45987\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45984\
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__45990\,
            I => \ppm_encoder_1.aileronZ0Z_0\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__45987\,
            I => \ppm_encoder_1.aileronZ0Z_0\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__45984\,
            I => \ppm_encoder_1.aileronZ0Z_0\
        );

    \I__10628\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45974\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__45974\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__10626\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45968\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__45968\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45965\,
            I => \N__45961\
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__45964\,
            I => \N__45958\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__45961\,
            I => \N__45955\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45951\
        );

    \I__10620\ : Span4Mux_v
    port map (
            O => \N__45955\,
            I => \N__45948\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45945\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__45951\,
            I => \N__45940\
        );

    \I__10617\ : Span4Mux_h
    port map (
            O => \N__45948\,
            I => \N__45940\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__45945\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__10615\ : Odrv4
    port map (
            O => \N__45940\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__10614\ : CascadeMux
    port map (
            O => \N__45935\,
            I => \N__45929\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__45934\,
            I => \N__45926\
        );

    \I__10612\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45921\
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__45932\,
            I => \N__45918\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45929\,
            I => \N__45915\
        );

    \I__10609\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45912\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45925\,
            I => \N__45909\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45906\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__45921\,
            I => \N__45902\
        );

    \I__10605\ : InMux
    port map (
            O => \N__45918\,
            I => \N__45899\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__45915\,
            I => \N__45894\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45891\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45884\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__45906\,
            I => \N__45884\
        );

    \I__10600\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45881\
        );

    \I__10599\ : Span4Mux_h
    port map (
            O => \N__45902\,
            I => \N__45876\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__45899\,
            I => \N__45876\
        );

    \I__10597\ : InMux
    port map (
            O => \N__45898\,
            I => \N__45873\
        );

    \I__10596\ : InMux
    port map (
            O => \N__45897\,
            I => \N__45870\
        );

    \I__10595\ : Span4Mux_v
    port map (
            O => \N__45894\,
            I => \N__45865\
        );

    \I__10594\ : Span4Mux_v
    port map (
            O => \N__45891\,
            I => \N__45865\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45862\
        );

    \I__10592\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45859\
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__45884\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45881\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__45876\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__45873\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__45870\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10586\ : Odrv4
    port map (
            O => \N__45865\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__45862\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__45859\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__10583\ : CascadeMux
    port map (
            O => \N__45842\,
            I => \N__45836\
        );

    \I__10582\ : CascadeMux
    port map (
            O => \N__45841\,
            I => \N__45833\
        );

    \I__10581\ : CascadeMux
    port map (
            O => \N__45840\,
            I => \N__45826\
        );

    \I__10580\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45823\
        );

    \I__10579\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45820\
        );

    \I__10578\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45817\
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__45832\,
            I => \N__45814\
        );

    \I__10576\ : CascadeMux
    port map (
            O => \N__45831\,
            I => \N__45810\
        );

    \I__10575\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45807\
        );

    \I__10574\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45804\
        );

    \I__10573\ : InMux
    port map (
            O => \N__45826\,
            I => \N__45799\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__45823\,
            I => \N__45796\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__45820\,
            I => \N__45793\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45790\
        );

    \I__10569\ : InMux
    port map (
            O => \N__45814\,
            I => \N__45787\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__45813\,
            I => \N__45782\
        );

    \I__10567\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45779\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__45807\,
            I => \N__45774\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45804\,
            I => \N__45774\
        );

    \I__10564\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45771\
        );

    \I__10563\ : InMux
    port map (
            O => \N__45802\,
            I => \N__45768\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__45799\,
            I => \N__45765\
        );

    \I__10561\ : Span4Mux_v
    port map (
            O => \N__45796\,
            I => \N__45756\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__45793\,
            I => \N__45756\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__45790\,
            I => \N__45756\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__45787\,
            I => \N__45756\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45753\
        );

    \I__10556\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45748\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45748\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__45779\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10553\ : Odrv4
    port map (
            O => \N__45774\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45771\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__45768\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__45765\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10549\ : Odrv4
    port map (
            O => \N__45756\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__45753\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__45748\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__10546\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45728\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__45728\,
            I => \N__45724\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45721\
        );

    \I__10543\ : Span4Mux_v
    port map (
            O => \N__45724\,
            I => \N__45718\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45721\,
            I => \N__45715\
        );

    \I__10541\ : Odrv4
    port map (
            O => \N__45718\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__10540\ : Odrv4
    port map (
            O => \N__45715\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__45710\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\
        );

    \I__10538\ : CascadeMux
    port map (
            O => \N__45707\,
            I => \N__45704\
        );

    \I__10537\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45701\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__45701\,
            I => \N__45698\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__45698\,
            I => \N__45695\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__45695\,
            I => \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45689\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__45689\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7\
        );

    \I__10531\ : CascadeMux
    port map (
            O => \N__45686\,
            I => \ppm_encoder_1.N_293_cascade_\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45683\,
            I => \N__45680\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__45680\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__45674\,
            I => \N__45671\
        );

    \I__10526\ : Span4Mux_h
    port map (
            O => \N__45671\,
            I => \N__45668\
        );

    \I__10525\ : Span4Mux_h
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10524\ : Odrv4
    port map (
            O => \N__45665\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45655\
        );

    \I__10521\ : CascadeMux
    port map (
            O => \N__45658\,
            I => \N__45651\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__45655\,
            I => \N__45648\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45645\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45651\,
            I => \N__45642\
        );

    \I__10517\ : Span12Mux_s11_h
    port map (
            O => \N__45648\,
            I => \N__45639\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__45645\,
            I => \N__45636\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45642\,
            I => side_order_7
        );

    \I__10514\ : Odrv12
    port map (
            O => \N__45639\,
            I => side_order_7
        );

    \I__10513\ : Odrv4
    port map (
            O => \N__45636\,
            I => side_order_7
        );

    \I__10512\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45620\
        );

    \I__10511\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45620\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45620\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__45620\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45614\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45614\,
            I => \N__45611\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__45611\,
            I => \N__45608\
        );

    \I__10505\ : Odrv4
    port map (
            O => \N__45608\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45602\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45602\,
            I => \N__45598\
        );

    \I__10502\ : CascadeMux
    port map (
            O => \N__45601\,
            I => \N__45594\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__45598\,
            I => \N__45591\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45588\
        );

    \I__10499\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45585\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__45591\,
            I => \N__45582\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45588\,
            I => \N__45579\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45585\,
            I => front_order_7
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__45582\,
            I => front_order_7
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__45579\,
            I => front_order_7
        );

    \I__10493\ : InMux
    port map (
            O => \N__45572\,
            I => \N__45563\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45571\,
            I => \N__45563\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45563\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45563\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45557\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45557\,
            I => \N__45554\
        );

    \I__10487\ : Span4Mux_v
    port map (
            O => \N__45554\,
            I => \N__45551\
        );

    \I__10486\ : Span4Mux_h
    port map (
            O => \N__45551\,
            I => \N__45548\
        );

    \I__10485\ : Odrv4
    port map (
            O => \N__45548\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__10484\ : CascadeMux
    port map (
            O => \N__45545\,
            I => \N__45541\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45544\,
            I => \N__45538\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45535\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45531\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45528\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45525\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45520\
        );

    \I__10477\ : Span4Mux_h
    port map (
            O => \N__45528\,
            I => \N__45520\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45525\,
            I => \N__45517\
        );

    \I__10475\ : Odrv4
    port map (
            O => \N__45520\,
            I => throttle_order_7
        );

    \I__10474\ : Odrv12
    port map (
            O => \N__45517\,
            I => throttle_order_7
        );

    \I__10473\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45503\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45503\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45503\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__45503\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45495\
        );

    \I__10468\ : CascadeMux
    port map (
            O => \N__45499\,
            I => \N__45491\
        );

    \I__10467\ : CascadeMux
    port map (
            O => \N__45498\,
            I => \N__45488\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45495\,
            I => \N__45485\
        );

    \I__10465\ : CascadeMux
    port map (
            O => \N__45494\,
            I => \N__45482\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45479\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45473\
        );

    \I__10462\ : Span4Mux_h
    port map (
            O => \N__45485\,
            I => \N__45470\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45482\,
            I => \N__45467\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45479\,
            I => \N__45464\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45461\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45458\
        );

    \I__10457\ : InMux
    port map (
            O => \N__45476\,
            I => \N__45455\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45473\,
            I => \N__45449\
        );

    \I__10455\ : Span4Mux_v
    port map (
            O => \N__45470\,
            I => \N__45444\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45467\,
            I => \N__45441\
        );

    \I__10453\ : Span4Mux_v
    port map (
            O => \N__45464\,
            I => \N__45435\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__45461\,
            I => \N__45435\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45458\,
            I => \N__45430\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__45455\,
            I => \N__45430\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45425\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45425\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__45452\,
            I => \N__45419\
        );

    \I__10446\ : Span4Mux_h
    port map (
            O => \N__45449\,
            I => \N__45416\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45411\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45447\,
            I => \N__45411\
        );

    \I__10443\ : Span4Mux_h
    port map (
            O => \N__45444\,
            I => \N__45406\
        );

    \I__10442\ : Span4Mux_h
    port map (
            O => \N__45441\,
            I => \N__45406\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45403\
        );

    \I__10440\ : Span4Mux_h
    port map (
            O => \N__45435\,
            I => \N__45396\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__45430\,
            I => \N__45396\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45396\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45393\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45388\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45388\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45385\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__45416\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45411\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10431\ : Odrv4
    port map (
            O => \N__45406\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45403\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10429\ : Odrv4
    port map (
            O => \N__45396\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45393\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45388\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45385\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__45368\,
            I => \N__45363\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45367\,
            I => \N__45357\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45354\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45349\
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__45362\,
            I => \N__45346\
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__45361\,
            I => \N__45343\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__45360\,
            I => \N__45340\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45357\,
            I => \N__45333\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45333\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45330\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45327\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__45349\,
            I => \N__45324\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45321\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45343\,
            I => \N__45318\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45315\
        );

    \I__10410\ : CascadeMux
    port map (
            O => \N__45339\,
            I => \N__45311\
        );

    \I__10409\ : CascadeMux
    port map (
            O => \N__45338\,
            I => \N__45305\
        );

    \I__10408\ : Span4Mux_v
    port map (
            O => \N__45333\,
            I => \N__45299\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__45330\,
            I => \N__45299\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__45327\,
            I => \N__45288\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__45324\,
            I => \N__45288\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45321\,
            I => \N__45288\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45318\,
            I => \N__45288\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__45315\,
            I => \N__45288\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45285\
        );

    \I__10400\ : InMux
    port map (
            O => \N__45311\,
            I => \N__45282\
        );

    \I__10399\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45277\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45309\,
            I => \N__45277\
        );

    \I__10397\ : InMux
    port map (
            O => \N__45308\,
            I => \N__45274\
        );

    \I__10396\ : InMux
    port map (
            O => \N__45305\,
            I => \N__45269\
        );

    \I__10395\ : InMux
    port map (
            O => \N__45304\,
            I => \N__45269\
        );

    \I__10394\ : Odrv4
    port map (
            O => \N__45299\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__45288\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__45285\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__45282\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45277\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45274\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45269\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45250\
        );

    \I__10386\ : CascadeMux
    port map (
            O => \N__45253\,
            I => \N__45247\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__45250\,
            I => \N__45244\
        );

    \I__10384\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45241\
        );

    \I__10383\ : Span4Mux_h
    port map (
            O => \N__45244\,
            I => \N__45237\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__45241\,
            I => \N__45234\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45240\,
            I => \N__45231\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__45237\,
            I => \N__45226\
        );

    \I__10379\ : Span4Mux_h
    port map (
            O => \N__45234\,
            I => \N__45226\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45231\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__10377\ : Odrv4
    port map (
            O => \N__45226\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__10376\ : CascadeMux
    port map (
            O => \N__45221\,
            I => \N__45215\
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__45220\,
            I => \N__45212\
        );

    \I__10374\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45202\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45202\
        );

    \I__10372\ : InMux
    port map (
            O => \N__45215\,
            I => \N__45202\
        );

    \I__10371\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45202\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45199\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__45202\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_153_d\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__45199\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_153_d\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__45194\,
            I => \N__45191\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45185\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45185\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__45185\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__10363\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45175\
        );

    \I__10362\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45175\
        );

    \I__10361\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45172\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__45175\,
            I => \N__45169\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45172\,
            I => \N__45164\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__45169\,
            I => \N__45164\
        );

    \I__10357\ : Odrv4
    port map (
            O => \N__45164\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__10356\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45153\
        );

    \I__10355\ : CascadeMux
    port map (
            O => \N__45160\,
            I => \N__45149\
        );

    \I__10354\ : CascadeMux
    port map (
            O => \N__45159\,
            I => \N__45145\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__45158\,
            I => \N__45141\
        );

    \I__10352\ : CascadeMux
    port map (
            O => \N__45157\,
            I => \N__45137\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45128\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45153\,
            I => \N__45118\
        );

    \I__10349\ : InMux
    port map (
            O => \N__45152\,
            I => \N__45111\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45149\,
            I => \N__45111\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45148\,
            I => \N__45111\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45145\,
            I => \N__45106\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45144\,
            I => \N__45106\
        );

    \I__10344\ : InMux
    port map (
            O => \N__45141\,
            I => \N__45101\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45140\,
            I => \N__45101\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45092\
        );

    \I__10341\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45092\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45092\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45092\
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__45133\,
            I => \N__45086\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45082\
        );

    \I__10336\ : CascadeMux
    port map (
            O => \N__45131\,
            I => \N__45079\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__45128\,
            I => \N__45075\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45127\,
            I => \N__45066\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45066\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45125\,
            I => \N__45066\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45124\,
            I => \N__45066\
        );

    \I__10330\ : CascadeMux
    port map (
            O => \N__45123\,
            I => \N__45063\
        );

    \I__10329\ : CascadeMux
    port map (
            O => \N__45122\,
            I => \N__45057\
        );

    \I__10328\ : CascadeMux
    port map (
            O => \N__45121\,
            I => \N__45053\
        );

    \I__10327\ : Span4Mux_h
    port map (
            O => \N__45118\,
            I => \N__45046\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45111\,
            I => \N__45046\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__45106\,
            I => \N__45043\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45101\,
            I => \N__45038\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__45092\,
            I => \N__45038\
        );

    \I__10322\ : CascadeMux
    port map (
            O => \N__45091\,
            I => \N__45035\
        );

    \I__10321\ : CascadeMux
    port map (
            O => \N__45090\,
            I => \N__45032\
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__45089\,
            I => \N__45025\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45086\,
            I => \N__45020\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45085\,
            I => \N__45017\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__45082\,
            I => \N__45014\
        );

    \I__10316\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45009\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45009\
        );

    \I__10314\ : Span4Mux_v
    port map (
            O => \N__45075\,
            I => \N__45004\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45066\,
            I => \N__45004\
        );

    \I__10312\ : InMux
    port map (
            O => \N__45063\,
            I => \N__44995\
        );

    \I__10311\ : InMux
    port map (
            O => \N__45062\,
            I => \N__44995\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45061\,
            I => \N__44995\
        );

    \I__10309\ : InMux
    port map (
            O => \N__45060\,
            I => \N__44995\
        );

    \I__10308\ : InMux
    port map (
            O => \N__45057\,
            I => \N__44984\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45056\,
            I => \N__44984\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45053\,
            I => \N__44984\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45052\,
            I => \N__44984\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45051\,
            I => \N__44984\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__45046\,
            I => \N__44977\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__45043\,
            I => \N__44977\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__45038\,
            I => \N__44977\
        );

    \I__10300\ : InMux
    port map (
            O => \N__45035\,
            I => \N__44968\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45032\,
            I => \N__44968\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45031\,
            I => \N__44968\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45030\,
            I => \N__44968\
        );

    \I__10296\ : InMux
    port map (
            O => \N__45029\,
            I => \N__44959\
        );

    \I__10295\ : InMux
    port map (
            O => \N__45028\,
            I => \N__44959\
        );

    \I__10294\ : InMux
    port map (
            O => \N__45025\,
            I => \N__44959\
        );

    \I__10293\ : InMux
    port map (
            O => \N__45024\,
            I => \N__44959\
        );

    \I__10292\ : InMux
    port map (
            O => \N__45023\,
            I => \N__44956\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__45020\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__45017\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__45014\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45009\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__45004\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__44995\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44984\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__44977\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44968\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44959\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__44956\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__10280\ : CascadeMux
    port map (
            O => \N__44933\,
            I => \N__44927\
        );

    \I__10279\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44904\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44904\
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__44930\,
            I => \N__44901\
        );

    \I__10276\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44893\
        );

    \I__10275\ : InMux
    port map (
            O => \N__44926\,
            I => \N__44888\
        );

    \I__10274\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44888\
        );

    \I__10273\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44879\
        );

    \I__10272\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44879\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44879\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44921\,
            I => \N__44879\
        );

    \I__10269\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44874\
        );

    \I__10268\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44874\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44918\,
            I => \N__44865\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44865\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44865\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44865\
        );

    \I__10263\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44862\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__44913\,
            I => \N__44854\
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__44912\,
            I => \N__44836\
        );

    \I__10260\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44819\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44910\,
            I => \N__44819\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44819\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__44904\,
            I => \N__44816\
        );

    \I__10256\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44811\
        );

    \I__10255\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44811\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44806\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44806\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44801\
        );

    \I__10251\ : InMux
    port map (
            O => \N__44896\,
            I => \N__44801\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__44893\,
            I => \N__44796\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__44888\,
            I => \N__44796\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44793\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44874\,
            I => \N__44788\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44865\,
            I => \N__44788\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__44862\,
            I => \N__44783\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44861\,
            I => \N__44772\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44860\,
            I => \N__44772\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44772\
        );

    \I__10241\ : InMux
    port map (
            O => \N__44858\,
            I => \N__44772\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44857\,
            I => \N__44772\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44757\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44757\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44757\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44851\,
            I => \N__44757\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44757\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44757\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44757\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44748\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44846\,
            I => \N__44748\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44845\,
            I => \N__44748\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44748\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44739\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44739\
        );

    \I__10226\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44739\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44739\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44839\,
            I => \N__44726\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44836\,
            I => \N__44726\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44726\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44726\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44726\
        );

    \I__10219\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44726\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44711\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44711\
        );

    \I__10216\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44711\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44828\,
            I => \N__44711\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44711\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44826\,
            I => \N__44708\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44819\,
            I => \N__44703\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__44816\,
            I => \N__44703\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44811\,
            I => \N__44700\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__44806\,
            I => \N__44689\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__44801\,
            I => \N__44689\
        );

    \I__10207\ : Span4Mux_v
    port map (
            O => \N__44796\,
            I => \N__44689\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__44793\,
            I => \N__44689\
        );

    \I__10205\ : Span4Mux_h
    port map (
            O => \N__44788\,
            I => \N__44689\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44684\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44786\,
            I => \N__44684\
        );

    \I__10202\ : Span4Mux_v
    port map (
            O => \N__44783\,
            I => \N__44679\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__44772\,
            I => \N__44679\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44757\,
            I => \N__44670\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44670\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__44739\,
            I => \N__44670\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44726\,
            I => \N__44670\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__44725\,
            I => \N__44663\
        );

    \I__10195\ : CascadeMux
    port map (
            O => \N__44724\,
            I => \N__44660\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44655\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44655\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44711\,
            I => \N__44652\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__44708\,
            I => \N__44649\
        );

    \I__10190\ : Span4Mux_v
    port map (
            O => \N__44703\,
            I => \N__44646\
        );

    \I__10189\ : Span4Mux_h
    port map (
            O => \N__44700\,
            I => \N__44641\
        );

    \I__10188\ : Span4Mux_v
    port map (
            O => \N__44689\,
            I => \N__44641\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__44684\,
            I => \N__44634\
        );

    \I__10186\ : Span4Mux_h
    port map (
            O => \N__44679\,
            I => \N__44634\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44670\,
            I => \N__44634\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44669\,
            I => \N__44627\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44627\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44627\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44624\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44621\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44660\,
            I => \N__44618\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__44655\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10177\ : Odrv4
    port map (
            O => \N__44652\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10176\ : Odrv4
    port map (
            O => \N__44649\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10175\ : Odrv4
    port map (
            O => \N__44646\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10174\ : Odrv4
    port map (
            O => \N__44641\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10173\ : Odrv4
    port map (
            O => \N__44634\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__44627\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44624\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44621\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44618\,
            I => \ppm_encoder_1.PPM_STATE_53_d\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44594\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__44594\,
            I => \N__44591\
        );

    \I__10166\ : Odrv4
    port map (
            O => \N__44591\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44585\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44582\
        );

    \I__10163\ : Odrv12
    port map (
            O => \N__44582\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44579\,
            I => \N__44576\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44576\,
            I => \N__44573\
        );

    \I__10160\ : Span4Mux_v
    port map (
            O => \N__44573\,
            I => \N__44570\
        );

    \I__10159\ : Span4Mux_h
    port map (
            O => \N__44570\,
            I => \N__44567\
        );

    \I__10158\ : Odrv4
    port map (
            O => \N__44567\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44561\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44558\,
            I => \N__44555\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44555\,
            I => \N__44552\
        );

    \I__10153\ : Span4Mux_v
    port map (
            O => \N__44552\,
            I => \N__44549\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44549\,
            I => \N__44546\
        );

    \I__10151\ : Odrv4
    port map (
            O => \N__44546\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__44543\,
            I => \N__44540\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44537\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__44537\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44534\,
            I => \N__44531\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44528\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__44528\,
            I => \N__44525\
        );

    \I__10144\ : Odrv4
    port map (
            O => \N__44525\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44519\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__44519\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44513\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44510\
        );

    \I__10139\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44507\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__44507\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\
        );

    \I__10137\ : CascadeMux
    port map (
            O => \N__44504\,
            I => \N__44495\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44503\,
            I => \N__44477\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44502\,
            I => \N__44477\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44501\,
            I => \N__44477\
        );

    \I__10133\ : InMux
    port map (
            O => \N__44500\,
            I => \N__44477\
        );

    \I__10132\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44477\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44474\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44464\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44494\,
            I => \N__44464\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44464\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44464\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44455\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44455\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44455\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44455\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44477\,
            I => \N__44452\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44474\,
            I => \N__44449\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44446\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44464\,
            I => \N__44443\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44455\,
            I => \N__44440\
        );

    \I__10117\ : Span4Mux_v
    port map (
            O => \N__44452\,
            I => \N__44437\
        );

    \I__10116\ : Span12Mux_v
    port map (
            O => \N__44449\,
            I => \N__44434\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44446\,
            I => \N__44427\
        );

    \I__10114\ : Span12Mux_s8_h
    port map (
            O => \N__44443\,
            I => \N__44427\
        );

    \I__10113\ : Span12Mux_v
    port map (
            O => \N__44440\,
            I => \N__44427\
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__44437\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__10111\ : Odrv12
    port map (
            O => \N__44434\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__10110\ : Odrv12
    port map (
            O => \N__44427\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44420\,
            I => \N__44417\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44417\,
            I => \N__44414\
        );

    \I__10107\ : Odrv4
    port map (
            O => \N__44414\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__10106\ : CEMux
    port map (
            O => \N__44411\,
            I => \N__44405\
        );

    \I__10105\ : CEMux
    port map (
            O => \N__44410\,
            I => \N__44401\
        );

    \I__10104\ : CEMux
    port map (
            O => \N__44409\,
            I => \N__44398\
        );

    \I__10103\ : CEMux
    port map (
            O => \N__44408\,
            I => \N__44395\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44405\,
            I => \N__44392\
        );

    \I__10101\ : CEMux
    port map (
            O => \N__44404\,
            I => \N__44389\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44386\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44398\,
            I => \N__44383\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44395\,
            I => \N__44378\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__44392\,
            I => \N__44378\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44375\
        );

    \I__10095\ : Span4Mux_h
    port map (
            O => \N__44386\,
            I => \N__44372\
        );

    \I__10094\ : Span4Mux_h
    port map (
            O => \N__44383\,
            I => \N__44369\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__44378\,
            I => \N__44366\
        );

    \I__10092\ : Odrv12
    port map (
            O => \N__44375\,
            I => \ppm_encoder_1.N_1818_0\
        );

    \I__10091\ : Odrv4
    port map (
            O => \N__44372\,
            I => \ppm_encoder_1.N_1818_0\
        );

    \I__10090\ : Odrv4
    port map (
            O => \N__44369\,
            I => \ppm_encoder_1.N_1818_0\
        );

    \I__10089\ : Odrv4
    port map (
            O => \N__44366\,
            I => \ppm_encoder_1.N_1818_0\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44354\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__44351\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44345\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__10083\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44339\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__44339\,
            I => \N__44336\
        );

    \I__10081\ : Span4Mux_h
    port map (
            O => \N__44336\,
            I => \N__44333\
        );

    \I__10080\ : Span4Mux_h
    port map (
            O => \N__44333\,
            I => \N__44330\
        );

    \I__10079\ : Odrv4
    port map (
            O => \N__44330\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44324\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44324\,
            I => \N__44321\
        );

    \I__10076\ : Span4Mux_h
    port map (
            O => \N__44321\,
            I => \N__44318\
        );

    \I__10075\ : Odrv4
    port map (
            O => \N__44318\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44315\,
            I => \N__44312\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__44312\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__10072\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__10070\ : Odrv12
    port map (
            O => \N__44303\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44300\,
            I => \N__44297\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44297\,
            I => \N__44294\
        );

    \I__10067\ : Span4Mux_h
    port map (
            O => \N__44294\,
            I => \N__44291\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__44291\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44282\
        );

    \I__10063\ : Span12Mux_v
    port map (
            O => \N__44282\,
            I => \N__44279\
        );

    \I__10062\ : Odrv12
    port map (
            O => \N__44279\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__10061\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44273\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44270\
        );

    \I__10059\ : Span4Mux_h
    port map (
            O => \N__44270\,
            I => \N__44267\
        );

    \I__10058\ : Span4Mux_h
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__44264\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44261\,
            I => \N__44255\
        );

    \I__10055\ : InMux
    port map (
            O => \N__44260\,
            I => \N__44255\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44255\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44249\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__44249\,
            I => \N__44246\
        );

    \I__10051\ : Span4Mux_h
    port map (
            O => \N__44246\,
            I => \N__44241\
        );

    \I__10050\ : InMux
    port map (
            O => \N__44245\,
            I => \N__44236\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44236\
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__44241\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44236\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__44231\,
            I => \N__44227\
        );

    \I__10045\ : CascadeMux
    port map (
            O => \N__44230\,
            I => \N__44224\
        );

    \I__10044\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44219\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44224\,
            I => \N__44219\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__44219\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44216\,
            I => \N__44212\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44215\,
            I => \N__44209\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__44212\,
            I => \N__44206\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44209\,
            I => \N__44203\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__44206\,
            I => \N__44197\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__44203\,
            I => \N__44197\
        );

    \I__10035\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44194\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__44197\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__44194\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__10032\ : InMux
    port map (
            O => \N__44189\,
            I => \N__44185\
        );

    \I__10031\ : InMux
    port map (
            O => \N__44188\,
            I => \N__44182\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44185\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__44182\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44177\,
            I => \N__44174\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44171\
        );

    \I__10026\ : Span4Mux_v
    port map (
            O => \N__44171\,
            I => \N__44167\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44164\
        );

    \I__10024\ : Span4Mux_v
    port map (
            O => \N__44167\,
            I => \N__44158\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44164\,
            I => \N__44158\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44155\
        );

    \I__10021\ : Odrv4
    port map (
            O => \N__44158\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__44155\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44147\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__44147\,
            I => \N__44143\
        );

    \I__10017\ : InMux
    port map (
            O => \N__44146\,
            I => \N__44140\
        );

    \I__10016\ : Span4Mux_v
    port map (
            O => \N__44143\,
            I => \N__44135\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__44140\,
            I => \N__44135\
        );

    \I__10014\ : Span4Mux_v
    port map (
            O => \N__44135\,
            I => \N__44132\
        );

    \I__10013\ : Span4Mux_h
    port map (
            O => \N__44132\,
            I => \N__44129\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__44129\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__10011\ : InMux
    port map (
            O => \N__44126\,
            I => \N__44123\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__44123\,
            I => \N__44119\
        );

    \I__10009\ : InMux
    port map (
            O => \N__44122\,
            I => \N__44116\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__44119\,
            I => \N__44111\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__44116\,
            I => \N__44111\
        );

    \I__10006\ : Span4Mux_v
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__44108\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44105\,
            I => \N__44102\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44097\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44101\,
            I => \N__44094\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44091\
        );

    \I__10000\ : Span4Mux_v
    port map (
            O => \N__44097\,
            I => \N__44088\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44083\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44083\
        );

    \I__9997\ : Odrv4
    port map (
            O => \N__44088\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9996\ : Odrv12
    port map (
            O => \N__44083\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44074\
        );

    \I__9994\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44071\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__44074\,
            I => \N__44068\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__44071\,
            I => \N__44065\
        );

    \I__9991\ : Span4Mux_v
    port map (
            O => \N__44068\,
            I => \N__44062\
        );

    \I__9990\ : Span4Mux_h
    port map (
            O => \N__44065\,
            I => \N__44059\
        );

    \I__9989\ : Odrv4
    port map (
            O => \N__44062\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__9988\ : Odrv4
    port map (
            O => \N__44059\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44051\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__44051\,
            I => \N__44048\
        );

    \I__9985\ : Span4Mux_h
    port map (
            O => \N__44048\,
            I => \N__44045\
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__44045\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44039\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44035\
        );

    \I__9981\ : CascadeMux
    port map (
            O => \N__44038\,
            I => \N__44031\
        );

    \I__9980\ : Span4Mux_h
    port map (
            O => \N__44035\,
            I => \N__44028\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44034\,
            I => \N__44025\
        );

    \I__9978\ : InMux
    port map (
            O => \N__44031\,
            I => \N__44022\
        );

    \I__9977\ : Span4Mux_h
    port map (
            O => \N__44028\,
            I => \N__44017\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__44017\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__44022\,
            I => throttle_order_0
        );

    \I__9974\ : Odrv4
    port map (
            O => \N__44017\,
            I => throttle_order_0
        );

    \I__9973\ : InMux
    port map (
            O => \N__44012\,
            I => \N__44007\
        );

    \I__9972\ : InMux
    port map (
            O => \N__44011\,
            I => \N__44004\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44000\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__44007\,
            I => \N__43995\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__44004\,
            I => \N__43995\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43992\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__44000\,
            I => \N__43987\
        );

    \I__9966\ : Span4Mux_v
    port map (
            O => \N__43995\,
            I => \N__43987\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43982\
        );

    \I__9964\ : Span4Mux_h
    port map (
            O => \N__43987\,
            I => \N__43982\
        );

    \I__9963\ : Odrv4
    port map (
            O => \N__43982\,
            I => \ppm_encoder_1.elevatorZ0Z_0\
        );

    \I__9962\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43974\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43978\,
            I => \N__43969\
        );

    \I__9960\ : InMux
    port map (
            O => \N__43977\,
            I => \N__43969\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43966\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__43969\,
            I => \N__43961\
        );

    \I__9957\ : Span4Mux_v
    port map (
            O => \N__43966\,
            I => \N__43961\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__43961\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__9955\ : InMux
    port map (
            O => \N__43958\,
            I => \N__43955\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__43955\,
            I => \N__43950\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43947\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43941\
        );

    \I__9951\ : Span4Mux_h
    port map (
            O => \N__43950\,
            I => \N__43936\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__43947\,
            I => \N__43936\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43946\,
            I => \N__43929\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43929\
        );

    \I__9947\ : InMux
    port map (
            O => \N__43944\,
            I => \N__43929\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__43941\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9945\ : Odrv4
    port map (
            O => \N__43936\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__43929\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__43922\,
            I => \ppm_encoder_1.N_286_cascade_\
        );

    \I__9942\ : InMux
    port map (
            O => \N__43919\,
            I => \N__43916\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__43916\,
            I => \N__43913\
        );

    \I__9940\ : Span4Mux_h
    port map (
            O => \N__43913\,
            I => \N__43910\
        );

    \I__9939\ : Span4Mux_v
    port map (
            O => \N__43910\,
            I => \N__43907\
        );

    \I__9938\ : Odrv4
    port map (
            O => \N__43907\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\
        );

    \I__9937\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43899\
        );

    \I__9936\ : InMux
    port map (
            O => \N__43903\,
            I => \N__43896\
        );

    \I__9935\ : InMux
    port map (
            O => \N__43902\,
            I => \N__43893\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__43899\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__43896\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__43893\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__9931\ : CascadeMux
    port map (
            O => \N__43886\,
            I => \N__43883\
        );

    \I__9930\ : InMux
    port map (
            O => \N__43883\,
            I => \N__43875\
        );

    \I__9929\ : InMux
    port map (
            O => \N__43882\,
            I => \N__43875\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43872\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43866\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__43875\,
            I => \N__43861\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__43872\,
            I => \N__43861\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43871\,
            I => \N__43856\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43870\,
            I => \N__43856\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43853\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43849\
        );

    \I__9920\ : Span4Mux_v
    port map (
            O => \N__43861\,
            I => \N__43844\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__43856\,
            I => \N__43844\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__43853\,
            I => \N__43841\
        );

    \I__9917\ : CascadeMux
    port map (
            O => \N__43852\,
            I => \N__43836\
        );

    \I__9916\ : Span12Mux_v
    port map (
            O => \N__43849\,
            I => \N__43828\
        );

    \I__9915\ : Span4Mux_v
    port map (
            O => \N__43844\,
            I => \N__43825\
        );

    \I__9914\ : Span4Mux_h
    port map (
            O => \N__43841\,
            I => \N__43822\
        );

    \I__9913\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43819\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43816\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43811\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43835\,
            I => \N__43811\
        );

    \I__9909\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43806\
        );

    \I__9908\ : InMux
    port map (
            O => \N__43833\,
            I => \N__43806\
        );

    \I__9907\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43801\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43831\,
            I => \N__43801\
        );

    \I__9905\ : Odrv12
    port map (
            O => \N__43828\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__43825\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__43822\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__43819\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43816\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__43811\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__43806\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43801\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__9897\ : CascadeMux
    port map (
            O => \N__43784\,
            I => \N__43779\
        );

    \I__9896\ : CascadeMux
    port map (
            O => \N__43783\,
            I => \N__43773\
        );

    \I__9895\ : InMux
    port map (
            O => \N__43782\,
            I => \N__43767\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43767\
        );

    \I__9893\ : CascadeMux
    port map (
            O => \N__43778\,
            I => \N__43763\
        );

    \I__9892\ : CascadeMux
    port map (
            O => \N__43777\,
            I => \N__43758\
        );

    \I__9891\ : CascadeMux
    port map (
            O => \N__43776\,
            I => \N__43754\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43773\,
            I => \N__43750\
        );

    \I__9889\ : CascadeMux
    port map (
            O => \N__43772\,
            I => \N__43746\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__43767\,
            I => \N__43743\
        );

    \I__9887\ : InMux
    port map (
            O => \N__43766\,
            I => \N__43740\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43736\
        );

    \I__9885\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43729\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43761\,
            I => \N__43729\
        );

    \I__9883\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43729\
        );

    \I__9882\ : InMux
    port map (
            O => \N__43757\,
            I => \N__43723\
        );

    \I__9881\ : InMux
    port map (
            O => \N__43754\,
            I => \N__43723\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43753\,
            I => \N__43720\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__43750\,
            I => \N__43717\
        );

    \I__9878\ : InMux
    port map (
            O => \N__43749\,
            I => \N__43712\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43712\
        );

    \I__9876\ : Span4Mux_v
    port map (
            O => \N__43743\,
            I => \N__43705\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__43740\,
            I => \N__43705\
        );

    \I__9874\ : CascadeMux
    port map (
            O => \N__43739\,
            I => \N__43702\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__43736\,
            I => \N__43696\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43729\,
            I => \N__43696\
        );

    \I__9871\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43693\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43688\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N__43688\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__43717\,
            I => \N__43683\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__43712\,
            I => \N__43683\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43711\,
            I => \N__43678\
        );

    \I__9865\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43678\
        );

    \I__9864\ : Span4Mux_v
    port map (
            O => \N__43705\,
            I => \N__43675\
        );

    \I__9863\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43672\
        );

    \I__9862\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43669\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__43696\,
            I => \N__43662\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__43693\,
            I => \N__43662\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__43688\,
            I => \N__43662\
        );

    \I__9858\ : Span4Mux_v
    port map (
            O => \N__43683\,
            I => \N__43655\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43655\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__43675\,
            I => \N__43655\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43672\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__43669\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__43662\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9852\ : Odrv4
    port map (
            O => \N__43655\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43643\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__43643\,
            I => \N__43639\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43636\
        );

    \I__9848\ : Span4Mux_v
    port map (
            O => \N__43639\,
            I => \N__43633\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43636\,
            I => \N__43630\
        );

    \I__9846\ : Odrv4
    port map (
            O => \N__43633\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__9845\ : Odrv12
    port map (
            O => \N__43630\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43622\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43622\,
            I => \drone_H_disp_front_i_9\
        );

    \I__9842\ : CascadeMux
    port map (
            O => \N__43619\,
            I => \N__43616\
        );

    \I__9841\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43613\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__43613\,
            I => front_command_5
        );

    \I__9839\ : InMux
    port map (
            O => \N__43610\,
            I => \N__43607\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43607\,
            I => \N__43604\
        );

    \I__9837\ : Span12Mux_s8_h
    port map (
            O => \N__43604\,
            I => \N__43601\
        );

    \I__9836\ : Odrv12
    port map (
            O => \N__43601\,
            I => \pid_front.error_9\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43598\,
            I => \pid_front.error_cry_4\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43595\,
            I => \N__43592\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43592\,
            I => \N__43589\
        );

    \I__9832\ : Odrv4
    port map (
            O => \N__43589\,
            I => front_command_6
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__43586\,
            I => \N__43583\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43580\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43580\,
            I => \drone_H_disp_front_i_10\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43574\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43574\,
            I => \N__43571\
        );

    \I__9826\ : Span4Mux_s3_h
    port map (
            O => \N__43571\,
            I => \N__43568\
        );

    \I__9825\ : Span4Mux_h
    port map (
            O => \N__43568\,
            I => \N__43565\
        );

    \I__9824\ : Odrv4
    port map (
            O => \N__43565\,
            I => \pid_front.error_10\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43562\,
            I => \pid_front.error_cry_5\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43556\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__43556\,
            I => \pid_front.error_axbZ0Z_7\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43550\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43547\
        );

    \I__9818\ : Span4Mux_v
    port map (
            O => \N__43547\,
            I => \N__43544\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__43544\,
            I => \N__43541\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__43541\,
            I => \pid_front.error_11\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43538\,
            I => \pid_front.error_cry_6\
        );

    \I__9814\ : InMux
    port map (
            O => \N__43535\,
            I => \N__43532\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43532\,
            I => \pid_front.error_axb_8_l_ofx_0\
        );

    \I__9812\ : CascadeMux
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43522\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43519\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43522\,
            I => \N__43515\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43519\,
            I => \N__43512\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43509\
        );

    \I__9806\ : Span4Mux_h
    port map (
            O => \N__43515\,
            I => \N__43504\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__43512\,
            I => \N__43504\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43509\,
            I => \drone_H_disp_front_12\
        );

    \I__9803\ : Odrv4
    port map (
            O => \N__43504\,
            I => \drone_H_disp_front_12\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43496\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43493\
        );

    \I__9800\ : Span4Mux_v
    port map (
            O => \N__43493\,
            I => \N__43490\
        );

    \I__9799\ : Span4Mux_h
    port map (
            O => \N__43490\,
            I => \N__43487\
        );

    \I__9798\ : Odrv4
    port map (
            O => \N__43487\,
            I => \pid_front.error_12\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43484\,
            I => \pid_front.error_cry_7\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43481\,
            I => \N__43478\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43475\
        );

    \I__9794\ : Odrv12
    port map (
            O => \N__43475\,
            I => \drone_H_disp_front_i_12\
        );

    \I__9793\ : CascadeMux
    port map (
            O => \N__43472\,
            I => \N__43469\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43465\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43462\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43465\,
            I => \N__43459\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43456\
        );

    \I__9788\ : Odrv4
    port map (
            O => \N__43459\,
            I => \drone_H_disp_front_13\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__43456\,
            I => \drone_H_disp_front_13\
        );

    \I__9786\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43448\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__43448\,
            I => \N__43445\
        );

    \I__9784\ : Span4Mux_v
    port map (
            O => \N__43445\,
            I => \N__43442\
        );

    \I__9783\ : Span4Mux_h
    port map (
            O => \N__43442\,
            I => \N__43439\
        );

    \I__9782\ : Odrv4
    port map (
            O => \N__43439\,
            I => \pid_front.error_13\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43436\,
            I => \pid_front.error_cry_8\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43433\,
            I => \N__43430\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43430\,
            I => \N__43427\
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__43427\,
            I => \drone_H_disp_front_i_13\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43424\,
            I => \N__43421\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43421\,
            I => \N__43418\
        );

    \I__9775\ : Span4Mux_s3_h
    port map (
            O => \N__43418\,
            I => \N__43415\
        );

    \I__9774\ : Span4Mux_h
    port map (
            O => \N__43415\,
            I => \N__43412\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__43412\,
            I => \pid_front.error_14\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43409\,
            I => \pid_front.error_cry_9\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43403\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__43403\,
            I => \N__43400\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__43400\,
            I => \N__43397\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__43397\,
            I => \drone_H_disp_front_15\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43394\,
            I => \pid_front.error_cry_10\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43388\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43385\
        );

    \I__9764\ : Span4Mux_s3_h
    port map (
            O => \N__43385\,
            I => \N__43382\
        );

    \I__9763\ : Span4Mux_h
    port map (
            O => \N__43382\,
            I => \N__43379\
        );

    \I__9762\ : Odrv4
    port map (
            O => \N__43379\,
            I => \pid_front.error_15\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43376\,
            I => \N__43367\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43367\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__43374\,
            I => \N__43363\
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__43373\,
            I => \N__43355\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43347\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43367\,
            I => \N__43344\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43341\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43363\,
            I => \N__43338\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43362\,
            I => \N__43331\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43361\,
            I => \N__43331\
        );

    \I__9751\ : InMux
    port map (
            O => \N__43360\,
            I => \N__43331\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43326\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43326\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43323\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43354\,
            I => \N__43318\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43318\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43311\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43311\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43311\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43347\,
            I => \N__43305\
        );

    \I__9741\ : Span4Mux_v
    port map (
            O => \N__43344\,
            I => \N__43300\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__43341\,
            I => \N__43300\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__43338\,
            I => \N__43287\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__43331\,
            I => \N__43287\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43326\,
            I => \N__43287\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43323\,
            I => \N__43287\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43318\,
            I => \N__43287\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N__43287\
        );

    \I__9733\ : InMux
    port map (
            O => \N__43310\,
            I => \N__43280\
        );

    \I__9732\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43280\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43308\,
            I => \N__43280\
        );

    \I__9730\ : Span4Mux_v
    port map (
            O => \N__43305\,
            I => \N__43275\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__43300\,
            I => \N__43275\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__43287\,
            I => \N__43272\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43269\
        );

    \I__9726\ : Span4Mux_v
    port map (
            O => \N__43275\,
            I => \N__43266\
        );

    \I__9725\ : Span4Mux_v
    port map (
            O => \N__43272\,
            I => \N__43263\
        );

    \I__9724\ : Odrv12
    port map (
            O => \N__43269\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__43266\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43263\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43256\,
            I => \N__43253\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43253\,
            I => \N__43250\
        );

    \I__9719\ : Span4Mux_h
    port map (
            O => \N__43250\,
            I => \N__43247\
        );

    \I__9718\ : Odrv4
    port map (
            O => \N__43247\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__43244\,
            I => \N__43233\
        );

    \I__9716\ : CascadeMux
    port map (
            O => \N__43243\,
            I => \N__43230\
        );

    \I__9715\ : CascadeMux
    port map (
            O => \N__43242\,
            I => \N__43227\
        );

    \I__9714\ : CascadeMux
    port map (
            O => \N__43241\,
            I => \N__43224\
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__43240\,
            I => \N__43215\
        );

    \I__9712\ : CascadeMux
    port map (
            O => \N__43239\,
            I => \N__43212\
        );

    \I__9711\ : CascadeMux
    port map (
            O => \N__43238\,
            I => \N__43209\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43204\
        );

    \I__9709\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43204\
        );

    \I__9708\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43201\
        );

    \I__9707\ : InMux
    port map (
            O => \N__43230\,
            I => \N__43196\
        );

    \I__9706\ : InMux
    port map (
            O => \N__43227\,
            I => \N__43196\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43224\,
            I => \N__43193\
        );

    \I__9704\ : InMux
    port map (
            O => \N__43223\,
            I => \N__43190\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43185\
        );

    \I__9702\ : InMux
    port map (
            O => \N__43221\,
            I => \N__43185\
        );

    \I__9701\ : CascadeMux
    port map (
            O => \N__43220\,
            I => \N__43182\
        );

    \I__9700\ : CascadeMux
    port map (
            O => \N__43219\,
            I => \N__43179\
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__43218\,
            I => \N__43172\
        );

    \I__9698\ : InMux
    port map (
            O => \N__43215\,
            I => \N__43167\
        );

    \I__9697\ : InMux
    port map (
            O => \N__43212\,
            I => \N__43167\
        );

    \I__9696\ : InMux
    port map (
            O => \N__43209\,
            I => \N__43164\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__43204\,
            I => \N__43161\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__43201\,
            I => \N__43156\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__43196\,
            I => \N__43156\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__43193\,
            I => \N__43149\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43190\,
            I => \N__43149\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43185\,
            I => \N__43149\
        );

    \I__9689\ : InMux
    port map (
            O => \N__43182\,
            I => \N__43146\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43141\
        );

    \I__9687\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43141\
        );

    \I__9686\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43136\
        );

    \I__9685\ : InMux
    port map (
            O => \N__43176\,
            I => \N__43136\
        );

    \I__9684\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43133\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43172\,
            I => \N__43130\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43125\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43164\,
            I => \N__43125\
        );

    \I__9680\ : Span4Mux_h
    port map (
            O => \N__43161\,
            I => \N__43122\
        );

    \I__9679\ : Span4Mux_h
    port map (
            O => \N__43156\,
            I => \N__43117\
        );

    \I__9678\ : Span4Mux_h
    port map (
            O => \N__43149\,
            I => \N__43117\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43146\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__43141\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__43136\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43133\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__43130\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9672\ : Odrv12
    port map (
            O => \N__43125\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__43122\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9670\ : Odrv4
    port map (
            O => \N__43117\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__9669\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43097\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__43097\,
            I => \N__43094\
        );

    \I__9667\ : Span4Mux_h
    port map (
            O => \N__43094\,
            I => \N__43091\
        );

    \I__9666\ : Odrv4
    port map (
            O => \N__43091\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__9665\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43085\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__43085\,
            I => \N__43082\
        );

    \I__9663\ : Span12Mux_s9_v
    port map (
            O => \N__43082\,
            I => \N__43079\
        );

    \I__9662\ : Odrv12
    port map (
            O => \N__43079\,
            I => \pid_front.error_axbZ0Z_2\
        );

    \I__9661\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43073\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__43073\,
            I => \N__43070\
        );

    \I__9659\ : Span12Mux_s8_h
    port map (
            O => \N__43070\,
            I => \N__43067\
        );

    \I__9658\ : Odrv12
    port map (
            O => \N__43067\,
            I => \pid_front.error_2\
        );

    \I__9657\ : InMux
    port map (
            O => \N__43064\,
            I => \pid_front.error_cry_1\
        );

    \I__9656\ : InMux
    port map (
            O => \N__43061\,
            I => \N__43058\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__43058\,
            I => \N__43055\
        );

    \I__9654\ : Span4Mux_h
    port map (
            O => \N__43055\,
            I => \N__43052\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__43052\,
            I => \N__43049\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__43049\,
            I => \pid_front.error_axbZ0Z_3\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43046\,
            I => \N__43043\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__43043\,
            I => \N__43040\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9648\ : Span4Mux_h
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9647\ : Odrv4
    port map (
            O => \N__43034\,
            I => \pid_front.error_3\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43031\,
            I => \pid_front.error_cry_2\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43028\,
            I => \N__43025\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__43025\,
            I => front_command_0
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__43022\,
            I => \N__43019\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43016\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__43016\,
            I => \drone_H_disp_front_i_4\
        );

    \I__9640\ : InMux
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__9638\ : Span4Mux_v
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__9637\ : Span4Mux_h
    port map (
            O => \N__43004\,
            I => \N__43001\
        );

    \I__9636\ : Odrv4
    port map (
            O => \N__43001\,
            I => \pid_front.error_4\
        );

    \I__9635\ : InMux
    port map (
            O => \N__42998\,
            I => \pid_front.error_cry_3\
        );

    \I__9634\ : InMux
    port map (
            O => \N__42995\,
            I => \N__42992\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__42992\,
            I => \drone_H_disp_front_i_5\
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__42989\,
            I => \N__42986\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42986\,
            I => \N__42983\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__42983\,
            I => front_command_1
        );

    \I__9629\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42977\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__42977\,
            I => \N__42974\
        );

    \I__9627\ : Span4Mux_s3_h
    port map (
            O => \N__42974\,
            I => \N__42971\
        );

    \I__9626\ : Span4Mux_h
    port map (
            O => \N__42971\,
            I => \N__42968\
        );

    \I__9625\ : Odrv4
    port map (
            O => \N__42968\,
            I => \pid_front.error_5\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42965\,
            I => \pid_front.error_cry_0_0\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__42959\,
            I => \drone_H_disp_front_i_6\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__42956\,
            I => \N__42953\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42950\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__42950\,
            I => front_command_2
        );

    \I__9618\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42944\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__42944\,
            I => \N__42941\
        );

    \I__9616\ : Span4Mux_s3_h
    port map (
            O => \N__42941\,
            I => \N__42938\
        );

    \I__9615\ : Span4Mux_h
    port map (
            O => \N__42938\,
            I => \N__42935\
        );

    \I__9614\ : Odrv4
    port map (
            O => \N__42935\,
            I => \pid_front.error_6\
        );

    \I__9613\ : InMux
    port map (
            O => \N__42932\,
            I => \pid_front.error_cry_1_0\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42926\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__42926\,
            I => \drone_H_disp_front_i_7\
        );

    \I__9610\ : CascadeMux
    port map (
            O => \N__42923\,
            I => \N__42920\
        );

    \I__9609\ : InMux
    port map (
            O => \N__42920\,
            I => \N__42917\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__42917\,
            I => front_command_3
        );

    \I__9607\ : InMux
    port map (
            O => \N__42914\,
            I => \N__42911\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__42911\,
            I => \N__42908\
        );

    \I__9605\ : Span4Mux_s3_h
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__9604\ : Span4Mux_h
    port map (
            O => \N__42905\,
            I => \N__42902\
        );

    \I__9603\ : Odrv4
    port map (
            O => \N__42902\,
            I => \pid_front.error_7\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42899\,
            I => \pid_front.error_cry_2_0\
        );

    \I__9601\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__42893\,
            I => front_command_4
        );

    \I__9599\ : CascadeMux
    port map (
            O => \N__42890\,
            I => \N__42887\
        );

    \I__9598\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42884\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__42881\,
            I => \N__42878\
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__42878\,
            I => \drone_H_disp_front_i_8\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42875\,
            I => \N__42872\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9592\ : Span4Mux_s3_h
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__9591\ : Span4Mux_h
    port map (
            O => \N__42866\,
            I => \N__42863\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__42863\,
            I => \pid_front.error_8\
        );

    \I__9589\ : InMux
    port map (
            O => \N__42860\,
            I => \bfn_17_24_0_\
        );

    \I__9588\ : CascadeMux
    port map (
            O => \N__42857\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\
        );

    \I__9587\ : CascadeMux
    port map (
            O => \N__42854\,
            I => \N__42850\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42853\,
            I => \N__42847\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42844\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42839\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__42844\,
            I => \N__42839\
        );

    \I__9582\ : Odrv4
    port map (
            O => \N__42839\,
            I => \ppm_encoder_1.N_139_17\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42836\,
            I => \N__42833\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__42833\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42824\
        );

    \I__9578\ : InMux
    port map (
            O => \N__42829\,
            I => \N__42824\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__42824\,
            I => \N__42821\
        );

    \I__9576\ : Odrv12
    port map (
            O => \N__42821\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__42818\,
            I => \N__42811\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__42817\,
            I => \N__42806\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__42816\,
            I => \N__42795\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__42815\,
            I => \N__42792\
        );

    \I__9571\ : InMux
    port map (
            O => \N__42814\,
            I => \N__42788\
        );

    \I__9570\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42785\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42810\,
            I => \N__42780\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42780\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42806\,
            I => \N__42777\
        );

    \I__9566\ : CascadeMux
    port map (
            O => \N__42805\,
            I => \N__42772\
        );

    \I__9565\ : CascadeMux
    port map (
            O => \N__42804\,
            I => \N__42768\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__42803\,
            I => \N__42765\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42802\,
            I => \N__42761\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42801\,
            I => \N__42756\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42756\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42751\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42751\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42744\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42744\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42744\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__42788\,
            I => \N__42737\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42737\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__42780\,
            I => \N__42737\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__42777\,
            I => \N__42734\
        );

    \I__9551\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42727\
        );

    \I__9550\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42727\
        );

    \I__9549\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42727\
        );

    \I__9548\ : CascadeMux
    port map (
            O => \N__42771\,
            I => \N__42723\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42716\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42716\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42716\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42761\,
            I => \N__42713\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42704\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__42751\,
            I => \N__42704\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__42744\,
            I => \N__42704\
        );

    \I__9540\ : Span4Mux_v
    port map (
            O => \N__42737\,
            I => \N__42704\
        );

    \I__9539\ : Span4Mux_v
    port map (
            O => \N__42734\,
            I => \N__42699\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42727\,
            I => \N__42699\
        );

    \I__9537\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42696\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42691\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__42716\,
            I => \N__42688\
        );

    \I__9534\ : Span4Mux_h
    port map (
            O => \N__42713\,
            I => \N__42683\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__42704\,
            I => \N__42683\
        );

    \I__9532\ : Sp12to4
    port map (
            O => \N__42699\,
            I => \N__42678\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42696\,
            I => \N__42678\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42695\,
            I => \N__42675\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42694\,
            I => \N__42672\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__42691\,
            I => \N__42662\
        );

    \I__9527\ : Span12Mux_h
    port map (
            O => \N__42688\,
            I => \N__42662\
        );

    \I__9526\ : Sp12to4
    port map (
            O => \N__42683\,
            I => \N__42662\
        );

    \I__9525\ : Span12Mux_h
    port map (
            O => \N__42678\,
            I => \N__42662\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42675\,
            I => \N__42657\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__42672\,
            I => \N__42657\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42654\
        );

    \I__9521\ : Span12Mux_v
    port map (
            O => \N__42662\,
            I => \N__42651\
        );

    \I__9520\ : Span4Mux_v
    port map (
            O => \N__42657\,
            I => \N__42648\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42654\,
            I => \pid_front.stateZ0Z_0\
        );

    \I__9518\ : Odrv12
    port map (
            O => \N__42651\,
            I => \pid_front.stateZ0Z_0\
        );

    \I__9517\ : Odrv4
    port map (
            O => \N__42648\,
            I => \pid_front.stateZ0Z_0\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42634\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42634\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42631\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42634\,
            I => \N__42627\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42631\,
            I => \N__42624\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42621\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__42627\,
            I => \N__42616\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__42624\,
            I => \N__42616\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42621\,
            I => \pid_front.pid_preregZ0Z_8\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__42616\,
            I => \pid_front.pid_preregZ0Z_8\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42607\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42602\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42607\,
            I => \N__42598\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42595\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42592\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42602\,
            I => \N__42589\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42586\
        );

    \I__9499\ : Span4Mux_h
    port map (
            O => \N__42598\,
            I => \N__42581\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42595\,
            I => \N__42581\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__42592\,
            I => \N__42578\
        );

    \I__9496\ : Span4Mux_v
    port map (
            O => \N__42589\,
            I => \N__42575\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42586\,
            I => \N__42572\
        );

    \I__9494\ : Span4Mux_v
    port map (
            O => \N__42581\,
            I => \N__42567\
        );

    \I__9493\ : Span4Mux_v
    port map (
            O => \N__42578\,
            I => \N__42564\
        );

    \I__9492\ : Span4Mux_h
    port map (
            O => \N__42575\,
            I => \N__42559\
        );

    \I__9491\ : Span4Mux_v
    port map (
            O => \N__42572\,
            I => \N__42559\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42556\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42553\
        );

    \I__9488\ : Span4Mux_h
    port map (
            O => \N__42567\,
            I => \N__42548\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__42564\,
            I => \N__42548\
        );

    \I__9486\ : Span4Mux_v
    port map (
            O => \N__42559\,
            I => \N__42543\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42556\,
            I => \N__42543\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42553\,
            I => \N__42540\
        );

    \I__9483\ : Span4Mux_v
    port map (
            O => \N__42548\,
            I => \N__42535\
        );

    \I__9482\ : Span4Mux_v
    port map (
            O => \N__42543\,
            I => \N__42535\
        );

    \I__9481\ : Span4Mux_h
    port map (
            O => \N__42540\,
            I => \N__42532\
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__42535\,
            I => uart_drone_data_0
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__42532\,
            I => uart_drone_data_0
        );

    \I__9478\ : CEMux
    port map (
            O => \N__42527\,
            I => \N__42523\
        );

    \I__9477\ : CEMux
    port map (
            O => \N__42526\,
            I => \N__42520\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42523\,
            I => \N__42516\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42520\,
            I => \N__42513\
        );

    \I__9474\ : CEMux
    port map (
            O => \N__42519\,
            I => \N__42510\
        );

    \I__9473\ : Span4Mux_h
    port map (
            O => \N__42516\,
            I => \N__42506\
        );

    \I__9472\ : Span4Mux_h
    port map (
            O => \N__42513\,
            I => \N__42501\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42510\,
            I => \N__42501\
        );

    \I__9470\ : CEMux
    port map (
            O => \N__42509\,
            I => \N__42498\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__42506\,
            I => \N__42495\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__42501\,
            I => \N__42492\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__42498\,
            I => \N__42489\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42495\,
            I => \dron_frame_decoder_1.N_731_0\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__42492\,
            I => \dron_frame_decoder_1.N_731_0\
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__42489\,
            I => \dron_frame_decoder_1.N_731_0\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42482\,
            I => \N__42479\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42479\,
            I => \N__42476\
        );

    \I__9461\ : Span4Mux_s3_h
    port map (
            O => \N__42476\,
            I => \N__42473\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__42473\,
            I => \N__42469\
        );

    \I__9459\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42466\
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__42469\,
            I => \drone_H_disp_front_0\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42466\,
            I => \drone_H_disp_front_0\
        );

    \I__9456\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42458\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42458\,
            I => \pid_front.error_axb_0\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42452\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42452\,
            I => \N__42449\
        );

    \I__9452\ : Span4Mux_v
    port map (
            O => \N__42449\,
            I => \N__42446\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__42446\,
            I => \pid_front.error_axbZ0Z_1\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42440\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42440\,
            I => \N__42437\
        );

    \I__9448\ : Span4Mux_v
    port map (
            O => \N__42437\,
            I => \N__42434\
        );

    \I__9447\ : Span4Mux_h
    port map (
            O => \N__42434\,
            I => \N__42431\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__42431\,
            I => \pid_front.error_1\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42428\,
            I => \pid_front.error_cry_0\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42412\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42424\,
            I => \N__42412\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42412\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42409\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42402\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42402\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42419\,
            I => \N__42402\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__42412\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__42409\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42402\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__9434\ : CascadeMux
    port map (
            O => \N__42395\,
            I => \N__42392\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42392\,
            I => \N__42389\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__42389\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42383\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42383\,
            I => \N__42380\
        );

    \I__9429\ : Span4Mux_v
    port map (
            O => \N__42380\,
            I => \N__42377\
        );

    \I__9428\ : Span4Mux_h
    port map (
            O => \N__42377\,
            I => \N__42374\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__42374\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42371\,
            I => \N__42368\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__42368\,
            I => \N__42365\
        );

    \I__9424\ : Span4Mux_v
    port map (
            O => \N__42365\,
            I => \N__42362\
        );

    \I__9423\ : Odrv4
    port map (
            O => \N__42362\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42359\,
            I => \N__42356\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42356\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42350\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__42350\,
            I => \N__42347\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__42347\,
            I => \N__42344\
        );

    \I__9417\ : Odrv4
    port map (
            O => \N__42344\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__9416\ : CascadeMux
    port map (
            O => \N__42341\,
            I => \N__42338\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42338\,
            I => \N__42335\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42335\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__9413\ : InMux
    port map (
            O => \N__42332\,
            I => \N__42329\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__42329\,
            I => \N__42326\
        );

    \I__9411\ : Span4Mux_v
    port map (
            O => \N__42326\,
            I => \N__42323\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__42323\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42320\,
            I => \N__42317\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42317\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__9407\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42311\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__42311\,
            I => \N__42308\
        );

    \I__9405\ : Span4Mux_v
    port map (
            O => \N__42308\,
            I => \N__42305\
        );

    \I__9404\ : Odrv4
    port map (
            O => \N__42305\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42302\,
            I => \N__42299\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__42299\,
            I => \N__42296\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__42296\,
            I => \N__42293\
        );

    \I__9400\ : Span4Mux_v
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__42290\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\
        );

    \I__9398\ : CascadeMux
    port map (
            O => \N__42287\,
            I => \N__42284\
        );

    \I__9397\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__42281\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__9395\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42273\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42270\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42267\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__42273\,
            I => \N__42264\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42270\,
            I => \ppm_encoder_1.aileronZ0Z_3\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__42267\,
            I => \ppm_encoder_1.aileronZ0Z_3\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__42264\,
            I => \ppm_encoder_1.aileronZ0Z_3\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42254\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__42254\,
            I => \N__42251\
        );

    \I__9386\ : Span4Mux_v
    port map (
            O => \N__42251\,
            I => \N__42248\
        );

    \I__9385\ : Span4Mux_h
    port map (
            O => \N__42248\,
            I => \N__42245\
        );

    \I__9384\ : Odrv4
    port map (
            O => \N__42245\,
            I => \ppm_encoder_1.N_289\
        );

    \I__9383\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42239\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__42239\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\
        );

    \I__9381\ : CascadeMux
    port map (
            O => \N__42236\,
            I => \ppm_encoder_1.PPM_STATE_53_d_cascade_\
        );

    \I__9380\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42230\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42230\,
            I => \N__42227\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__42227\,
            I => \N__42224\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__42224\,
            I => \ppm_encoder_1.N_134_0\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42214\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42209\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42209\
        );

    \I__9373\ : CascadeMux
    port map (
            O => \N__42218\,
            I => \N__42206\
        );

    \I__9372\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42201\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42214\,
            I => \N__42196\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42196\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42189\
        );

    \I__9368\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42189\
        );

    \I__9367\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42189\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__42201\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9365\ : Odrv12
    port map (
            O => \N__42196\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__42189\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42179\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42176\
        );

    \I__9361\ : Span12Mux_v
    port map (
            O => \N__42176\,
            I => \N__42168\
        );

    \I__9360\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42165\
        );

    \I__9359\ : InMux
    port map (
            O => \N__42174\,
            I => \N__42162\
        );

    \I__9358\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42155\
        );

    \I__9357\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42155\
        );

    \I__9356\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42155\
        );

    \I__9355\ : Odrv12
    port map (
            O => \N__42168\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__42165\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__42162\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42155\,
            I => \ppm_encoder_1.N_221\
        );

    \I__9351\ : CascadeMux
    port map (
            O => \N__42146\,
            I => \ppm_encoder_1.N_232_cascade_\
        );

    \I__9350\ : IoInMux
    port map (
            O => \N__42143\,
            I => \N__42140\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42140\,
            I => \N__42137\
        );

    \I__9348\ : Span12Mux_s1_v
    port map (
            O => \N__42137\,
            I => \N__42134\
        );

    \I__9347\ : Span12Mux_v
    port map (
            O => \N__42134\,
            I => \N__42131\
        );

    \I__9346\ : Odrv12
    port map (
            O => \N__42131\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__9345\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42125\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__42122\
        );

    \I__9343\ : Span4Mux_h
    port map (
            O => \N__42122\,
            I => \N__42119\
        );

    \I__9342\ : Span4Mux_h
    port map (
            O => \N__42119\,
            I => \N__42116\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__42116\,
            I => \ppm_encoder_1.N_139\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42107\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42112\,
            I => \N__42107\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42107\,
            I => \ppm_encoder_1.N_232\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42101\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__42101\,
            I => \N__42098\
        );

    \I__9335\ : Span4Mux_h
    port map (
            O => \N__42098\,
            I => \N__42094\
        );

    \I__9334\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42091\
        );

    \I__9333\ : Span4Mux_v
    port map (
            O => \N__42094\,
            I => \N__42088\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__42091\,
            I => \N__42081\
        );

    \I__9331\ : Span4Mux_h
    port map (
            O => \N__42088\,
            I => \N__42081\
        );

    \I__9330\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42078\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42086\,
            I => \N__42075\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__42081\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__42078\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42075\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42065\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__42065\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__42062\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__42059\,
            I => \N__42055\
        );

    \I__9321\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42052\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42055\,
            I => \N__42049\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__42052\,
            I => \N__42046\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__42049\,
            I => \N__42040\
        );

    \I__9317\ : Span4Mux_v
    port map (
            O => \N__42046\,
            I => \N__42040\
        );

    \I__9316\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42037\
        );

    \I__9315\ : Odrv4
    port map (
            O => \N__42040\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__42037\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__9313\ : InMux
    port map (
            O => \N__42032\,
            I => \N__42029\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__42026\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__42026\,
            I => \N__42023\
        );

    \I__9310\ : Odrv4
    port map (
            O => \N__42023\,
            I => \ppm_encoder_1.un1_init_pulses_10_0\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42020\,
            I => \N__42017\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__42017\,
            I => \N__42012\
        );

    \I__9307\ : InMux
    port map (
            O => \N__42016\,
            I => \N__42009\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42006\
        );

    \I__9305\ : Span4Mux_v
    port map (
            O => \N__42012\,
            I => \N__42003\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__42009\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42006\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__9302\ : Odrv4
    port map (
            O => \N__42003\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41992\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41989\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41986\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__41989\,
            I => \N__41983\
        );

    \I__9297\ : Span4Mux_h
    port map (
            O => \N__41986\,
            I => \N__41980\
        );

    \I__9296\ : Odrv12
    port map (
            O => \N__41983\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__9295\ : Odrv4
    port map (
            O => \N__41980\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41975\,
            I => \N__41972\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__41972\,
            I => \N__41967\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__41971\,
            I => \N__41964\
        );

    \I__9291\ : InMux
    port map (
            O => \N__41970\,
            I => \N__41961\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__41967\,
            I => \N__41958\
        );

    \I__9289\ : InMux
    port map (
            O => \N__41964\,
            I => \N__41955\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__41961\,
            I => \N__41952\
        );

    \I__9287\ : Span4Mux_h
    port map (
            O => \N__41958\,
            I => \N__41949\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__41955\,
            I => \ppm_encoder_1.elevatorZ0Z_3\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__41952\,
            I => \ppm_encoder_1.elevatorZ0Z_3\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__41949\,
            I => \ppm_encoder_1.elevatorZ0Z_3\
        );

    \I__9283\ : CascadeMux
    port map (
            O => \N__41942\,
            I => \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__41939\,
            I => \N__41936\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41933\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__41933\,
            I => \N__41930\
        );

    \I__9279\ : Span4Mux_h
    port map (
            O => \N__41930\,
            I => \N__41927\
        );

    \I__9278\ : Span4Mux_v
    port map (
            O => \N__41927\,
            I => \N__41924\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__41924\,
            I => \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\
        );

    \I__9276\ : InMux
    port map (
            O => \N__41921\,
            I => \N__41916\
        );

    \I__9275\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41913\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41910\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41905\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41913\,
            I => \N__41905\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41910\,
            I => \N__41902\
        );

    \I__9270\ : Span4Mux_v
    port map (
            O => \N__41905\,
            I => \N__41899\
        );

    \I__9269\ : Span4Mux_h
    port map (
            O => \N__41902\,
            I => \N__41896\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__41899\,
            I => \pid_side.pid_preregZ0Z_0\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__41896\,
            I => \pid_side.pid_preregZ0Z_0\
        );

    \I__9266\ : CEMux
    port map (
            O => \N__41891\,
            I => \N__41887\
        );

    \I__9265\ : CEMux
    port map (
            O => \N__41890\,
            I => \N__41884\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__41887\,
            I => \N__41881\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41884\,
            I => \N__41878\
        );

    \I__9262\ : Span4Mux_h
    port map (
            O => \N__41881\,
            I => \N__41875\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__41878\,
            I => \N__41872\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__41875\,
            I => \N__41869\
        );

    \I__9259\ : Span4Mux_h
    port map (
            O => \N__41872\,
            I => \N__41866\
        );

    \I__9258\ : Odrv4
    port map (
            O => \N__41869\,
            I => \pid_side.state_0_0\
        );

    \I__9257\ : Odrv4
    port map (
            O => \N__41866\,
            I => \pid_side.state_0_0\
        );

    \I__9256\ : CascadeMux
    port map (
            O => \N__41861\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\
        );

    \I__9255\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41855\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__41855\,
            I => \N__41852\
        );

    \I__9253\ : Span4Mux_h
    port map (
            O => \N__41852\,
            I => \N__41848\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41845\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__41848\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__41845\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__9249\ : CascadeMux
    port map (
            O => \N__41840\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__41837\,
            I => \N__41834\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41831\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41828\
        );

    \I__9245\ : Span4Mux_h
    port map (
            O => \N__41828\,
            I => \N__41825\
        );

    \I__9244\ : Odrv4
    port map (
            O => \N__41825\,
            I => \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\
        );

    \I__9243\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41819\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__41819\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41810\
        );

    \I__9240\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41810\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41810\,
            I => \N__41807\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__41807\,
            I => \N__41804\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__41804\,
            I => \N__41801\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__41801\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41792\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41792\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41792\,
            I => \N__41789\
        );

    \I__9232\ : Span12Mux_v
    port map (
            O => \N__41789\,
            I => \N__41786\
        );

    \I__9231\ : Odrv12
    port map (
            O => \N__41786\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__41783\,
            I => \ppm_encoder_1.N_300_cascade_\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41780\,
            I => \N__41774\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41779\,
            I => \N__41774\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41774\,
            I => \N__41771\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__41771\,
            I => \N__41768\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__41768\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__9224\ : CascadeMux
    port map (
            O => \N__41765\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_\
        );

    \I__9223\ : InMux
    port map (
            O => \N__41762\,
            I => \N__41759\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41759\,
            I => \N__41756\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__41756\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__9220\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41750\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41750\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__9218\ : CascadeMux
    port map (
            O => \N__41747\,
            I => \N__41742\
        );

    \I__9217\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41738\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41735\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41742\,
            I => \N__41730\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41741\,
            I => \N__41730\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__41738\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41735\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41730\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41717\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41714\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41709\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41720\,
            I => \N__41709\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41717\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41714\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41709\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__9203\ : CascadeMux
    port map (
            O => \N__41702\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41696\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41696\,
            I => \ppm_encoder_1.un2_throttle_iv_0_0\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41693\,
            I => \N__41688\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41685\
        );

    \I__9198\ : CascadeMux
    port map (
            O => \N__41691\,
            I => \N__41682\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41688\,
            I => \N__41679\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41685\,
            I => \N__41676\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41673\
        );

    \I__9194\ : Span4Mux_v
    port map (
            O => \N__41679\,
            I => \N__41668\
        );

    \I__9193\ : Span4Mux_v
    port map (
            O => \N__41676\,
            I => \N__41668\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41673\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__41668\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41660\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__41660\,
            I => \N__41656\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41659\,
            I => \N__41653\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__41656\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__41653\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__9185\ : CascadeMux
    port map (
            O => \N__41648\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__41645\,
            I => \N__41642\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41639\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41639\,
            I => \N__41636\
        );

    \I__9181\ : Span4Mux_v
    port map (
            O => \N__41636\,
            I => \N__41633\
        );

    \I__9180\ : Odrv4
    port map (
            O => \N__41633\,
            I => \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41627\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__41627\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13\
        );

    \I__9177\ : CascadeMux
    port map (
            O => \N__41624\,
            I => \ppm_encoder_1.N_299_cascade_\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__41621\,
            I => \N__41617\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__41620\,
            I => \N__41614\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41611\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41608\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__41611\,
            I => \N__41605\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41608\,
            I => \N__41602\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__41605\,
            I => \N__41599\
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__41602\,
            I => side_order_13
        );

    \I__9168\ : Odrv4
    port map (
            O => \N__41599\,
            I => side_order_13
        );

    \I__9167\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41591\,
            I => \N__41588\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__41588\,
            I => \N__41585\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__41585\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41573\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41581\,
            I => \N__41573\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41580\,
            I => \N__41573\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41573\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41570\,
            I => \N__41567\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41567\,
            I => \N__41564\
        );

    \I__9157\ : Span4Mux_v
    port map (
            O => \N__41564\,
            I => \N__41561\
        );

    \I__9156\ : Span4Mux_v
    port map (
            O => \N__41561\,
            I => \N__41557\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41560\,
            I => \N__41554\
        );

    \I__9154\ : Sp12to4
    port map (
            O => \N__41557\,
            I => \N__41549\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__41554\,
            I => \N__41549\
        );

    \I__9152\ : Odrv12
    port map (
            O => \N__41549\,
            I => front_order_13
        );

    \I__9151\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41543\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__41543\,
            I => \N__41540\
        );

    \I__9149\ : Span4Mux_h
    port map (
            O => \N__41540\,
            I => \N__41537\
        );

    \I__9148\ : Span4Mux_v
    port map (
            O => \N__41537\,
            I => \N__41534\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__41534\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41522\
        );

    \I__9145\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41522\
        );

    \I__9144\ : InMux
    port map (
            O => \N__41529\,
            I => \N__41522\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41522\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41516\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41516\,
            I => \N__41513\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__41513\,
            I => \N__41509\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__41512\,
            I => \N__41506\
        );

    \I__9138\ : Span4Mux_h
    port map (
            O => \N__41509\,
            I => \N__41503\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41500\
        );

    \I__9136\ : Odrv4
    port map (
            O => \N__41503\,
            I => throttle_order_13
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41500\,
            I => throttle_order_13
        );

    \I__9134\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__41492\,
            I => \N__41489\
        );

    \I__9132\ : Odrv12
    port map (
            O => \N__41489\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__41486\,
            I => \N__41481\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41476\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41476\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41473\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__41476\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__41473\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41464\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41461\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__41464\,
            I => \N__41458\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41461\,
            I => \N__41453\
        );

    \I__9121\ : Span4Mux_v
    port map (
            O => \N__41458\,
            I => \N__41453\
        );

    \I__9120\ : Span4Mux_h
    port map (
            O => \N__41453\,
            I => \N__41450\
        );

    \I__9119\ : Odrv4
    port map (
            O => \N__41450\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41444\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41444\,
            I => \N__41436\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41443\,
            I => \N__41433\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41424\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41441\,
            I => \N__41424\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41440\,
            I => \N__41424\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41424\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__41436\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41433\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41424\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__41417\,
            I => \N__41413\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41416\,
            I => \N__41410\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41406\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41410\,
            I => \N__41402\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41399\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__41406\,
            I => \N__41396\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41393\
        );

    \I__9101\ : Span4Mux_v
    port map (
            O => \N__41402\,
            I => \N__41388\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41399\,
            I => \N__41388\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__41396\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41393\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__41388\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__9096\ : CascadeMux
    port map (
            O => \N__41381\,
            I => \N__41378\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41375\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41375\,
            I => \ppm_encoder_1.un1_init_pulses_11_0\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41372\,
            I => \N__41369\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__41369\,
            I => \N__41364\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41368\,
            I => \N__41361\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__41367\,
            I => \N__41358\
        );

    \I__9089\ : Span4Mux_v
    port map (
            O => \N__41364\,
            I => \N__41353\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41361\,
            I => \N__41353\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41350\
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__41353\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_6\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__41350\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_6\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41341\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__41344\,
            I => \N__41338\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41341\,
            I => \N__41334\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41329\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41329\
        );

    \I__9079\ : Span4Mux_v
    port map (
            O => \N__41334\,
            I => \N__41318\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41329\,
            I => \N__41318\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41328\,
            I => \N__41309\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41309\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41326\,
            I => \N__41309\
        );

    \I__9074\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41309\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41306\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41323\,
            I => \N__41303\
        );

    \I__9071\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41298\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41298\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__41306\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__41303\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__9067\ : Odrv4
    port map (
            O => \N__41298\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\
        );

    \I__9066\ : CascadeMux
    port map (
            O => \N__41291\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__41285\,
            I => \N__41282\
        );

    \I__9063\ : Span4Mux_h
    port map (
            O => \N__41282\,
            I => \N__41279\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__41279\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__41276\,
            I => \N__41271\
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__41275\,
            I => \N__41267\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__41274\,
            I => \N__41264\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41256\
        );

    \I__9057\ : InMux
    port map (
            O => \N__41270\,
            I => \N__41256\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41267\,
            I => \N__41251\
        );

    \I__9055\ : InMux
    port map (
            O => \N__41264\,
            I => \N__41251\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41248\
        );

    \I__9053\ : InMux
    port map (
            O => \N__41262\,
            I => \N__41243\
        );

    \I__9052\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41243\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41256\,
            I => \N__41240\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41251\,
            I => \N__41237\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41234\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__41243\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__9047\ : Odrv4
    port map (
            O => \N__41240\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__41237\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__9045\ : Odrv12
    port map (
            O => \N__41234\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41225\,
            I => \N__41222\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41222\,
            I => \N__41217\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41221\,
            I => \N__41212\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41220\,
            I => \N__41212\
        );

    \I__9040\ : Odrv12
    port map (
            O => \N__41217\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__41212\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41204\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41204\,
            I => \N__41199\
        );

    \I__9036\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41196\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__41202\,
            I => \N__41193\
        );

    \I__9034\ : Span4Mux_v
    port map (
            O => \N__41199\,
            I => \N__41189\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__41196\,
            I => \N__41186\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41193\,
            I => \N__41183\
        );

    \I__9031\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41180\
        );

    \I__9030\ : Span4Mux_h
    port map (
            O => \N__41189\,
            I => \N__41175\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__41186\,
            I => \N__41175\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__41183\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41180\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__9026\ : Odrv4
    port map (
            O => \N__41175\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41163\
        );

    \I__9024\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41160\
        );

    \I__9023\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41157\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__41163\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__41160\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41157\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__9019\ : InMux
    port map (
            O => \N__41150\,
            I => \N__41145\
        );

    \I__9018\ : InMux
    port map (
            O => \N__41149\,
            I => \N__41142\
        );

    \I__9017\ : CascadeMux
    port map (
            O => \N__41148\,
            I => \N__41139\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__41145\,
            I => \N__41136\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__41142\,
            I => \N__41133\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41130\
        );

    \I__9013\ : Span4Mux_h
    port map (
            O => \N__41136\,
            I => \N__41127\
        );

    \I__9012\ : Span4Mux_v
    port map (
            O => \N__41133\,
            I => \N__41124\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41130\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__41127\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__41124\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__41117\,
            I => \N__41114\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41114\,
            I => \N__41108\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41113\,
            I => \N__41108\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41104\
        );

    \I__9004\ : CascadeMux
    port map (
            O => \N__41107\,
            I => \N__41101\
        );

    \I__9003\ : Span4Mux_h
    port map (
            O => \N__41104\,
            I => \N__41098\
        );

    \I__9002\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41095\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__41098\,
            I => \N__41092\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41095\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__41092\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__41084\,
            I => \N__41078\
        );

    \I__8996\ : InMux
    port map (
            O => \N__41083\,
            I => \N__41074\
        );

    \I__8995\ : InMux
    port map (
            O => \N__41082\,
            I => \N__41069\
        );

    \I__8994\ : InMux
    port map (
            O => \N__41081\,
            I => \N__41069\
        );

    \I__8993\ : Span4Mux_v
    port map (
            O => \N__41078\,
            I => \N__41066\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41077\,
            I => \N__41063\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__41074\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__41069\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__41066\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__41063\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41045\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41045\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41045\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__41045\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41042\,
            I => \N__41038\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41035\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__41038\,
            I => \N__41032\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__41035\,
            I => \N__41029\
        );

    \I__8979\ : Span4Mux_v
    port map (
            O => \N__41032\,
            I => \N__41026\
        );

    \I__8978\ : Span12Mux_v
    port map (
            O => \N__41029\,
            I => \N__41023\
        );

    \I__8977\ : Odrv4
    port map (
            O => \N__41026\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__8976\ : Odrv12
    port map (
            O => \N__41023\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41018\,
            I => \N__41015\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__41012\
        );

    \I__8973\ : Span4Mux_h
    port map (
            O => \N__41012\,
            I => \N__41009\
        );

    \I__8972\ : Odrv4
    port map (
            O => \N__41009\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__41006\,
            I => \N__41003\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41003\,
            I => \N__41000\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41000\,
            I => \N__40997\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__40997\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__8967\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40990\
        );

    \I__8966\ : CascadeMux
    port map (
            O => \N__40993\,
            I => \N__40987\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__40990\,
            I => \N__40984\
        );

    \I__8964\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40980\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__40984\,
            I => \N__40977\
        );

    \I__8962\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40974\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__40980\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__40977\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__40974\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__8958\ : InMux
    port map (
            O => \N__40967\,
            I => \N__40964\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__40964\,
            I => \N__40959\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40963\,
            I => \N__40954\
        );

    \I__8955\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40954\
        );

    \I__8954\ : Span4Mux_h
    port map (
            O => \N__40959\,
            I => \N__40951\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__40954\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__40951\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__40946\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40943\,
            I => \N__40938\
        );

    \I__8949\ : InMux
    port map (
            O => \N__40942\,
            I => \N__40933\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40941\,
            I => \N__40933\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40938\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__40933\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__40928\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\
        );

    \I__8944\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40921\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40924\,
            I => \N__40918\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__40921\,
            I => \N__40915\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__40918\,
            I => \N__40912\
        );

    \I__8940\ : Span4Mux_h
    port map (
            O => \N__40915\,
            I => \N__40908\
        );

    \I__8939\ : Span4Mux_h
    port map (
            O => \N__40912\,
            I => \N__40905\
        );

    \I__8938\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40902\
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__40908\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8936\ : Odrv4
    port map (
            O => \N__40905\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__40902\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40892\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__40892\,
            I => \N__40889\
        );

    \I__8932\ : Sp12to4
    port map (
            O => \N__40889\,
            I => \N__40884\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40881\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40878\
        );

    \I__8929\ : Span12Mux_v
    port map (
            O => \N__40884\,
            I => \N__40873\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40873\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40870\
        );

    \I__8926\ : Odrv12
    port map (
            O => \N__40873\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__8925\ : Odrv12
    port map (
            O => \N__40870\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40865\,
            I => \N__40862\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__40862\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40856\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__40856\,
            I => \N__40853\
        );

    \I__8920\ : Span4Mux_v
    port map (
            O => \N__40853\,
            I => \N__40850\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__40850\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40844\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__40844\,
            I => \N__40841\
        );

    \I__8916\ : Odrv4
    port map (
            O => \N__40841\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40838\,
            I => \N__40835\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__40835\,
            I => \N__40832\
        );

    \I__8913\ : Span4Mux_h
    port map (
            O => \N__40832\,
            I => \N__40829\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__40829\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__8911\ : CascadeMux
    port map (
            O => \N__40826\,
            I => \N__40823\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40820\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__40820\,
            I => \N__40817\
        );

    \I__8908\ : Odrv4
    port map (
            O => \N__40817\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40811\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__40811\,
            I => \N__40808\
        );

    \I__8905\ : Span4Mux_h
    port map (
            O => \N__40808\,
            I => \N__40805\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__40805\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40799\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40799\,
            I => \N__40796\
        );

    \I__8901\ : Odrv4
    port map (
            O => \N__40796\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40790\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40786\
        );

    \I__8898\ : InMux
    port map (
            O => \N__40789\,
            I => \N__40783\
        );

    \I__8897\ : Span4Mux_v
    port map (
            O => \N__40786\,
            I => \N__40778\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__40783\,
            I => \N__40778\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__40778\,
            I => \N__40775\
        );

    \I__8894\ : Sp12to4
    port map (
            O => \N__40775\,
            I => \N__40772\
        );

    \I__8893\ : Odrv12
    port map (
            O => \N__40772\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__8892\ : InMux
    port map (
            O => \N__40769\,
            I => \N__40766\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40766\,
            I => \N__40763\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__40763\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__8889\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40752\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40752\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40743\
        );

    \I__8886\ : InMux
    port map (
            O => \N__40757\,
            I => \N__40743\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40752\,
            I => \N__40740\
        );

    \I__8884\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40731\
        );

    \I__8883\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40731\
        );

    \I__8882\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40731\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40748\,
            I => \N__40731\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40728\
        );

    \I__8879\ : Span4Mux_h
    port map (
            O => \N__40740\,
            I => \N__40725\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40731\,
            I => \N__40722\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__40728\,
            I => \N__40719\
        );

    \I__8876\ : Odrv4
    port map (
            O => \N__40725\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__40722\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__40719\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8873\ : CascadeMux
    port map (
            O => \N__40712\,
            I => \N__40708\
        );

    \I__8872\ : CascadeMux
    port map (
            O => \N__40711\,
            I => \N__40701\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40695\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40695\
        );

    \I__8869\ : IoInMux
    port map (
            O => \N__40706\,
            I => \N__40688\
        );

    \I__8868\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40685\
        );

    \I__8867\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40682\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40677\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40700\,
            I => \N__40677\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__40695\,
            I => \N__40673\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40694\,
            I => \N__40670\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40663\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40663\
        );

    \I__8860\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40663\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__40688\,
            I => \N__40660\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40685\,
            I => \N__40657\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__40682\,
            I => \N__40654\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__40677\,
            I => \N__40651\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__40676\,
            I => \N__40647\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__40673\,
            I => \N__40644\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__40670\,
            I => \N__40638\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40663\,
            I => \N__40638\
        );

    \I__8851\ : Span4Mux_s2_v
    port map (
            O => \N__40660\,
            I => \N__40635\
        );

    \I__8850\ : Span4Mux_h
    port map (
            O => \N__40657\,
            I => \N__40630\
        );

    \I__8849\ : Span4Mux_v
    port map (
            O => \N__40654\,
            I => \N__40630\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__40651\,
            I => \N__40627\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40624\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40647\,
            I => \N__40621\
        );

    \I__8845\ : Sp12to4
    port map (
            O => \N__40644\,
            I => \N__40618\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40643\,
            I => \N__40615\
        );

    \I__8843\ : Span4Mux_v
    port map (
            O => \N__40638\,
            I => \N__40612\
        );

    \I__8842\ : Span4Mux_h
    port map (
            O => \N__40635\,
            I => \N__40605\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__40630\,
            I => \N__40605\
        );

    \I__8840\ : Span4Mux_v
    port map (
            O => \N__40627\,
            I => \N__40605\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__40624\,
            I => \N__40596\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__40621\,
            I => \N__40596\
        );

    \I__8837\ : Span12Mux_h
    port map (
            O => \N__40618\,
            I => \N__40596\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40615\,
            I => \N__40596\
        );

    \I__8835\ : Odrv4
    port map (
            O => \N__40612\,
            I => \debug_CH2_18A_c\
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__40605\,
            I => \debug_CH2_18A_c\
        );

    \I__8833\ : Odrv12
    port map (
            O => \N__40596\,
            I => \debug_CH2_18A_c\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40589\,
            I => \N__40586\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40586\,
            I => \N__40582\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40579\
        );

    \I__8829\ : Span4Mux_h
    port map (
            O => \N__40582\,
            I => \N__40576\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40579\,
            I => \N__40570\
        );

    \I__8827\ : Span4Mux_h
    port map (
            O => \N__40576\,
            I => \N__40570\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40567\
        );

    \I__8825\ : Odrv4
    port map (
            O => \N__40570\,
            I => \uart_pc.N_152\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40567\,
            I => \uart_pc.N_152\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__40562\,
            I => \N__40559\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40556\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40556\,
            I => \N__40553\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__40553\,
            I => \N__40550\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__40550\,
            I => \N__40547\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__40547\,
            I => \N__40544\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40544\,
            I => \N__40540\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40537\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__40540\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40537\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__8813\ : SRMux
    port map (
            O => \N__40532\,
            I => \N__40529\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__40529\,
            I => \N__40525\
        );

    \I__8811\ : SRMux
    port map (
            O => \N__40528\,
            I => \N__40521\
        );

    \I__8810\ : Span4Mux_h
    port map (
            O => \N__40525\,
            I => \N__40518\
        );

    \I__8809\ : SRMux
    port map (
            O => \N__40524\,
            I => \N__40515\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40512\
        );

    \I__8807\ : Span4Mux_h
    port map (
            O => \N__40518\,
            I => \N__40509\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40506\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__40512\,
            I => \N__40503\
        );

    \I__8804\ : Odrv4
    port map (
            O => \N__40509\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8803\ : Odrv4
    port map (
            O => \N__40506\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__40503\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40493\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__40493\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40487\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__40487\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40481\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__40481\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40475\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40475\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__40472\,
            I => \N__40469\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40466\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__40466\,
            I => \N__40461\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40456\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40456\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__40461\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__40456\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__40451\,
            I => \N__40448\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40448\,
            I => \N__40445\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40445\,
            I => \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__40442\,
            I => \N__40439\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40439\,
            I => \N__40436\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40436\,
            I => \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__40427\,
            I => \N__40422\
        );

    \I__8777\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40417\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40417\
        );

    \I__8775\ : Odrv4
    port map (
            O => \N__40422\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__40417\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__8773\ : CascadeMux
    port map (
            O => \N__40412\,
            I => \N__40409\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40406\,
            I => \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40397\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40392\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40389\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40386\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__40397\,
            I => \N__40383\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40396\,
            I => \N__40380\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40395\,
            I => \N__40375\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40370\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__40389\,
            I => \N__40370\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40386\,
            I => \N__40366\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__40383\,
            I => \N__40363\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40380\,
            I => \N__40360\
        );

    \I__8758\ : InMux
    port map (
            O => \N__40379\,
            I => \N__40356\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40353\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40375\,
            I => \N__40350\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__40370\,
            I => \N__40347\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40369\,
            I => \N__40344\
        );

    \I__8753\ : Span4Mux_h
    port map (
            O => \N__40366\,
            I => \N__40341\
        );

    \I__8752\ : Sp12to4
    port map (
            O => \N__40363\,
            I => \N__40338\
        );

    \I__8751\ : Span4Mux_h
    port map (
            O => \N__40360\,
            I => \N__40335\
        );

    \I__8750\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40332\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__40356\,
            I => \N__40329\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__40353\,
            I => \N__40324\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__40350\,
            I => \N__40324\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__40347\,
            I => \N__40317\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__40344\,
            I => \N__40317\
        );

    \I__8744\ : Span4Mux_h
    port map (
            O => \N__40341\,
            I => \N__40317\
        );

    \I__8743\ : Span12Mux_h
    port map (
            O => \N__40338\,
            I => \N__40312\
        );

    \I__8742\ : Sp12to4
    port map (
            O => \N__40335\,
            I => \N__40312\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40309\
        );

    \I__8740\ : Span4Mux_h
    port map (
            O => \N__40329\,
            I => \N__40306\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__40324\,
            I => \N__40301\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__40317\,
            I => \N__40301\
        );

    \I__8737\ : Span12Mux_v
    port map (
            O => \N__40312\,
            I => \N__40296\
        );

    \I__8736\ : Span4Mux_h
    port map (
            O => \N__40309\,
            I => \N__40291\
        );

    \I__8735\ : Span4Mux_h
    port map (
            O => \N__40306\,
            I => \N__40291\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__40301\,
            I => \N__40288\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40283\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40283\
        );

    \I__8731\ : Odrv12
    port map (
            O => \N__40296\,
            I => uart_pc_data_4
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__40291\,
            I => uart_pc_data_4
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__40288\,
            I => uart_pc_data_4
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__40283\,
            I => uart_pc_data_4
        );

    \I__8727\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40269\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40273\,
            I => \N__40266\
        );

    \I__8725\ : InMux
    port map (
            O => \N__40272\,
            I => \N__40263\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40269\,
            I => \N__40258\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40266\,
            I => \N__40251\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__40263\,
            I => \N__40247\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40243\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40240\
        );

    \I__8719\ : Span4Mux_h
    port map (
            O => \N__40258\,
            I => \N__40235\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40232\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40229\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40226\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40254\,
            I => \N__40223\
        );

    \I__8714\ : Span4Mux_h
    port map (
            O => \N__40251\,
            I => \N__40220\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40217\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__40247\,
            I => \N__40214\
        );

    \I__8711\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40211\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__40243\,
            I => \N__40208\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__40240\,
            I => \N__40205\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40200\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40200\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__40235\,
            I => \N__40195\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__40232\,
            I => \N__40195\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__40229\,
            I => \N__40189\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40226\,
            I => \N__40189\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40223\,
            I => \N__40184\
        );

    \I__8701\ : Span4Mux_h
    port map (
            O => \N__40220\,
            I => \N__40184\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__40217\,
            I => \N__40179\
        );

    \I__8699\ : Sp12to4
    port map (
            O => \N__40214\,
            I => \N__40179\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40211\,
            I => \N__40170\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__40208\,
            I => \N__40170\
        );

    \I__8696\ : Span4Mux_v
    port map (
            O => \N__40205\,
            I => \N__40170\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__40200\,
            I => \N__40170\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__40195\,
            I => \N__40167\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40164\
        );

    \I__8692\ : Span12Mux_v
    port map (
            O => \N__40189\,
            I => \N__40161\
        );

    \I__8691\ : Sp12to4
    port map (
            O => \N__40184\,
            I => \N__40156\
        );

    \I__8690\ : Span12Mux_s8_h
    port map (
            O => \N__40179\,
            I => \N__40156\
        );

    \I__8689\ : Span4Mux_h
    port map (
            O => \N__40170\,
            I => \N__40151\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__40167\,
            I => \N__40151\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__40164\,
            I => uart_pc_data_5
        );

    \I__8686\ : Odrv12
    port map (
            O => \N__40161\,
            I => uart_pc_data_5
        );

    \I__8685\ : Odrv12
    port map (
            O => \N__40156\,
            I => uart_pc_data_5
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__40151\,
            I => uart_pc_data_5
        );

    \I__8683\ : InMux
    port map (
            O => \N__40142\,
            I => \N__40135\
        );

    \I__8682\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40132\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40129\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40126\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40123\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40116\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40116\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__40129\,
            I => \N__40111\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40111\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__40123\,
            I => \N__40107\
        );

    \I__8673\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40103\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40100\
        );

    \I__8671\ : Span4Mux_v
    port map (
            O => \N__40116\,
            I => \N__40097\
        );

    \I__8670\ : Span4Mux_v
    port map (
            O => \N__40111\,
            I => \N__40094\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40110\,
            I => \N__40090\
        );

    \I__8668\ : Span4Mux_h
    port map (
            O => \N__40107\,
            I => \N__40087\
        );

    \I__8667\ : InMux
    port map (
            O => \N__40106\,
            I => \N__40084\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__40103\,
            I => \N__40081\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__40100\,
            I => \N__40078\
        );

    \I__8664\ : Sp12to4
    port map (
            O => \N__40097\,
            I => \N__40075\
        );

    \I__8663\ : Sp12to4
    port map (
            O => \N__40094\,
            I => \N__40072\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40069\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40090\,
            I => \N__40066\
        );

    \I__8660\ : Span4Mux_h
    port map (
            O => \N__40087\,
            I => \N__40063\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__40084\,
            I => \N__40060\
        );

    \I__8658\ : Span4Mux_v
    port map (
            O => \N__40081\,
            I => \N__40057\
        );

    \I__8657\ : Span12Mux_s10_v
    port map (
            O => \N__40078\,
            I => \N__40048\
        );

    \I__8656\ : Span12Mux_s5_h
    port map (
            O => \N__40075\,
            I => \N__40048\
        );

    \I__8655\ : Span12Mux_h
    port map (
            O => \N__40072\,
            I => \N__40048\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40048\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__40066\,
            I => \N__40045\
        );

    \I__8652\ : Span4Mux_v
    port map (
            O => \N__40063\,
            I => \N__40042\
        );

    \I__8651\ : Span4Mux_h
    port map (
            O => \N__40060\,
            I => \N__40037\
        );

    \I__8650\ : Sp12to4
    port map (
            O => \N__40057\,
            I => \N__40032\
        );

    \I__8649\ : Span12Mux_v
    port map (
            O => \N__40048\,
            I => \N__40032\
        );

    \I__8648\ : Span4Mux_h
    port map (
            O => \N__40045\,
            I => \N__40027\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__40042\,
            I => \N__40027\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40041\,
            I => \N__40022\
        );

    \I__8645\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40022\
        );

    \I__8644\ : Odrv4
    port map (
            O => \N__40037\,
            I => uart_pc_data_6
        );

    \I__8643\ : Odrv12
    port map (
            O => \N__40032\,
            I => uart_pc_data_6
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__40027\,
            I => uart_pc_data_6
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40022\,
            I => uart_pc_data_6
        );

    \I__8640\ : InMux
    port map (
            O => \N__40013\,
            I => \N__40007\
        );

    \I__8639\ : InMux
    port map (
            O => \N__40012\,
            I => \N__40002\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40011\,
            I => \N__39998\
        );

    \I__8637\ : InMux
    port map (
            O => \N__40010\,
            I => \N__39995\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__40007\,
            I => \N__39990\
        );

    \I__8635\ : InMux
    port map (
            O => \N__40006\,
            I => \N__39987\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40005\,
            I => \N__39984\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40002\,
            I => \N__39979\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39976\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__39998\,
            I => \N__39969\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__39995\,
            I => \N__39969\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39966\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39963\
        );

    \I__8627\ : Span4Mux_v
    port map (
            O => \N__39990\,
            I => \N__39960\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39987\,
            I => \N__39955\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__39984\,
            I => \N__39955\
        );

    \I__8624\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39952\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39949\
        );

    \I__8622\ : Span4Mux_h
    port map (
            O => \N__39979\,
            I => \N__39944\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__39976\,
            I => \N__39944\
        );

    \I__8620\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39939\
        );

    \I__8619\ : InMux
    port map (
            O => \N__39974\,
            I => \N__39939\
        );

    \I__8618\ : Span4Mux_v
    port map (
            O => \N__39969\,
            I => \N__39934\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39966\,
            I => \N__39934\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__39963\,
            I => \N__39931\
        );

    \I__8615\ : Span4Mux_h
    port map (
            O => \N__39960\,
            I => \N__39925\
        );

    \I__8614\ : Span4Mux_v
    port map (
            O => \N__39955\,
            I => \N__39925\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__39952\,
            I => \N__39918\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__39949\,
            I => \N__39918\
        );

    \I__8611\ : Span4Mux_v
    port map (
            O => \N__39944\,
            I => \N__39918\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39939\,
            I => \N__39915\
        );

    \I__8609\ : Span4Mux_v
    port map (
            O => \N__39934\,
            I => \N__39912\
        );

    \I__8608\ : Span12Mux_h
    port map (
            O => \N__39931\,
            I => \N__39909\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39906\
        );

    \I__8606\ : Span4Mux_v
    port map (
            O => \N__39925\,
            I => \N__39901\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39901\
        );

    \I__8604\ : Span4Mux_h
    port map (
            O => \N__39915\,
            I => \N__39898\
        );

    \I__8603\ : Span4Mux_h
    port map (
            O => \N__39912\,
            I => \N__39895\
        );

    \I__8602\ : Odrv12
    port map (
            O => \N__39909\,
            I => uart_pc_data_7
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__39906\,
            I => uart_pc_data_7
        );

    \I__8600\ : Odrv4
    port map (
            O => \N__39901\,
            I => uart_pc_data_7
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__39898\,
            I => uart_pc_data_7
        );

    \I__8598\ : Odrv4
    port map (
            O => \N__39895\,
            I => uart_pc_data_7
        );

    \I__8597\ : CEMux
    port map (
            O => \N__39884\,
            I => \N__39881\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39881\,
            I => \N__39878\
        );

    \I__8595\ : Span4Mux_v
    port map (
            O => \N__39878\,
            I => \N__39875\
        );

    \I__8594\ : Sp12to4
    port map (
            O => \N__39875\,
            I => \N__39872\
        );

    \I__8593\ : Span12Mux_h
    port map (
            O => \N__39872\,
            I => \N__39869\
        );

    \I__8592\ : Odrv12
    port map (
            O => \N__39869\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39866\,
            I => \N__39863\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__39863\,
            I => \dron_frame_decoder_1.drone_H_disp_front_10\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39857\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__39857\,
            I => \dron_frame_decoder_1.drone_H_disp_front_9\
        );

    \I__8587\ : InMux
    port map (
            O => \N__39854\,
            I => \N__39848\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39848\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__39848\,
            I => front_command_7
        );

    \I__8584\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39839\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39844\,
            I => \N__39839\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__39839\,
            I => \drone_H_disp_front_11\
        );

    \I__8581\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39833\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__39833\,
            I => \N__39830\
        );

    \I__8579\ : Span4Mux_h
    port map (
            O => \N__39830\,
            I => \N__39827\
        );

    \I__8578\ : Span4Mux_h
    port map (
            O => \N__39827\,
            I => \N__39824\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__39824\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__8576\ : CascadeMux
    port map (
            O => \N__39821\,
            I => \N__39818\
        );

    \I__8575\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39815\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39812\
        );

    \I__8573\ : Span4Mux_h
    port map (
            O => \N__39812\,
            I => \N__39808\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__8571\ : Span4Mux_h
    port map (
            O => \N__39808\,
            I => \N__39802\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39805\,
            I => \N__39799\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__39802\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39799\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__8567\ : InMux
    port map (
            O => \N__39794\,
            I => \N__39791\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__39791\,
            I => \dron_frame_decoder_1.drone_H_disp_front_4\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39788\,
            I => \N__39785\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__39785\,
            I => \dron_frame_decoder_1.drone_H_disp_front_5\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39779\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__39779\,
            I => \dron_frame_decoder_1.drone_H_disp_front_6\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39776\,
            I => \N__39773\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39773\,
            I => \dron_frame_decoder_1.drone_H_disp_front_7\
        );

    \I__8559\ : InMux
    port map (
            O => \N__39770\,
            I => \N__39765\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39762\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39756\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__39765\,
            I => \N__39750\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39762\,
            I => \N__39746\
        );

    \I__8554\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39743\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39760\,
            I => \N__39739\
        );

    \I__8552\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39736\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__39756\,
            I => \N__39733\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39730\
        );

    \I__8549\ : InMux
    port map (
            O => \N__39754\,
            I => \N__39727\
        );

    \I__8548\ : InMux
    port map (
            O => \N__39753\,
            I => \N__39724\
        );

    \I__8547\ : Span4Mux_v
    port map (
            O => \N__39750\,
            I => \N__39721\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39749\,
            I => \N__39718\
        );

    \I__8545\ : Span4Mux_v
    port map (
            O => \N__39746\,
            I => \N__39713\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39743\,
            I => \N__39713\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39710\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39739\,
            I => \N__39707\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39736\,
            I => \N__39699\
        );

    \I__8540\ : Sp12to4
    port map (
            O => \N__39733\,
            I => \N__39699\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__39730\,
            I => \N__39699\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39727\,
            I => \N__39692\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39724\,
            I => \N__39692\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__39721\,
            I => \N__39683\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39718\,
            I => \N__39683\
        );

    \I__8534\ : Span4Mux_h
    port map (
            O => \N__39713\,
            I => \N__39683\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__39710\,
            I => \N__39683\
        );

    \I__8532\ : Span12Mux_v
    port map (
            O => \N__39707\,
            I => \N__39680\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39706\,
            I => \N__39677\
        );

    \I__8530\ : Span12Mux_v
    port map (
            O => \N__39699\,
            I => \N__39674\
        );

    \I__8529\ : InMux
    port map (
            O => \N__39698\,
            I => \N__39669\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39697\,
            I => \N__39669\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__39692\,
            I => \N__39664\
        );

    \I__8526\ : Span4Mux_v
    port map (
            O => \N__39683\,
            I => \N__39664\
        );

    \I__8525\ : Odrv12
    port map (
            O => \N__39680\,
            I => uart_pc_data_0
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__39677\,
            I => uart_pc_data_0
        );

    \I__8523\ : Odrv12
    port map (
            O => \N__39674\,
            I => uart_pc_data_0
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39669\,
            I => uart_pc_data_0
        );

    \I__8521\ : Odrv4
    port map (
            O => \N__39664\,
            I => uart_pc_data_0
        );

    \I__8520\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39648\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39645\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39642\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__39648\,
            I => \N__39638\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39635\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39630\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39627\
        );

    \I__8513\ : Span4Mux_h
    port map (
            O => \N__39638\,
            I => \N__39620\
        );

    \I__8512\ : Span4Mux_v
    port map (
            O => \N__39635\,
            I => \N__39620\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39615\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39615\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__39630\,
            I => \N__39612\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__39627\,
            I => \N__39609\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39626\,
            I => \N__39606\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39603\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__39620\,
            I => \N__39598\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39615\,
            I => \N__39598\
        );

    \I__8503\ : Span4Mux_v
    port map (
            O => \N__39612\,
            I => \N__39595\
        );

    \I__8502\ : Span4Mux_v
    port map (
            O => \N__39609\,
            I => \N__39591\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39606\,
            I => \N__39588\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39603\,
            I => \N__39585\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__39598\,
            I => \N__39582\
        );

    \I__8498\ : Sp12to4
    port map (
            O => \N__39595\,
            I => \N__39578\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39594\,
            I => \N__39573\
        );

    \I__8496\ : Span4Mux_v
    port map (
            O => \N__39591\,
            I => \N__39570\
        );

    \I__8495\ : Span4Mux_v
    port map (
            O => \N__39588\,
            I => \N__39565\
        );

    \I__8494\ : Span4Mux_s3_h
    port map (
            O => \N__39585\,
            I => \N__39565\
        );

    \I__8493\ : Span4Mux_h
    port map (
            O => \N__39582\,
            I => \N__39562\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39559\
        );

    \I__8491\ : Span12Mux_h
    port map (
            O => \N__39578\,
            I => \N__39556\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39553\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39550\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39573\,
            I => \N__39541\
        );

    \I__8487\ : Span4Mux_v
    port map (
            O => \N__39570\,
            I => \N__39541\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__39565\,
            I => \N__39541\
        );

    \I__8485\ : Span4Mux_v
    port map (
            O => \N__39562\,
            I => \N__39541\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39559\,
            I => \N__39538\
        );

    \I__8483\ : Odrv12
    port map (
            O => \N__39556\,
            I => uart_pc_data_1
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39553\,
            I => uart_pc_data_1
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39550\,
            I => uart_pc_data_1
        );

    \I__8480\ : Odrv4
    port map (
            O => \N__39541\,
            I => uart_pc_data_1
        );

    \I__8479\ : Odrv4
    port map (
            O => \N__39538\,
            I => uart_pc_data_1
        );

    \I__8478\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39522\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39519\
        );

    \I__8476\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39516\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39522\,
            I => \N__39513\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__39519\,
            I => \N__39509\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__39516\,
            I => \N__39504\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__39513\,
            I => \N__39504\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39501\
        );

    \I__8470\ : Span4Mux_v
    port map (
            O => \N__39509\,
            I => \N__39492\
        );

    \I__8469\ : Span4Mux_h
    port map (
            O => \N__39504\,
            I => \N__39492\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39501\,
            I => \N__39489\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39500\,
            I => \N__39484\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39478\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39478\
        );

    \I__8464\ : CascadeMux
    port map (
            O => \N__39497\,
            I => \N__39475\
        );

    \I__8463\ : Span4Mux_v
    port map (
            O => \N__39492\,
            I => \N__39471\
        );

    \I__8462\ : Sp12to4
    port map (
            O => \N__39489\,
            I => \N__39468\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39488\,
            I => \N__39463\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39487\,
            I => \N__39460\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39484\,
            I => \N__39457\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39483\,
            I => \N__39454\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39478\,
            I => \N__39451\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39448\
        );

    \I__8455\ : CascadeMux
    port map (
            O => \N__39474\,
            I => \N__39445\
        );

    \I__8454\ : Sp12to4
    port map (
            O => \N__39471\,
            I => \N__39440\
        );

    \I__8453\ : Span12Mux_v
    port map (
            O => \N__39468\,
            I => \N__39440\
        );

    \I__8452\ : CascadeMux
    port map (
            O => \N__39467\,
            I => \N__39436\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39466\,
            I => \N__39433\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__39463\,
            I => \N__39430\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39460\,
            I => \N__39427\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__39457\,
            I => \N__39422\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39454\,
            I => \N__39422\
        );

    \I__8446\ : Span4Mux_v
    port map (
            O => \N__39451\,
            I => \N__39419\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39448\,
            I => \N__39416\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39445\,
            I => \N__39413\
        );

    \I__8443\ : Span12Mux_h
    port map (
            O => \N__39440\,
            I => \N__39410\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39439\,
            I => \N__39405\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39405\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39433\,
            I => \N__39394\
        );

    \I__8439\ : Span4Mux_h
    port map (
            O => \N__39430\,
            I => \N__39394\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__39427\,
            I => \N__39394\
        );

    \I__8437\ : Span4Mux_v
    port map (
            O => \N__39422\,
            I => \N__39394\
        );

    \I__8436\ : Span4Mux_v
    port map (
            O => \N__39419\,
            I => \N__39394\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__39416\,
            I => \N__39391\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__39413\,
            I => uart_pc_data_2
        );

    \I__8433\ : Odrv12
    port map (
            O => \N__39410\,
            I => uart_pc_data_2
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39405\,
            I => uart_pc_data_2
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__39394\,
            I => uart_pc_data_2
        );

    \I__8430\ : Odrv4
    port map (
            O => \N__39391\,
            I => uart_pc_data_2
        );

    \I__8429\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39377\,
            I => \N__39374\
        );

    \I__8427\ : Span4Mux_v
    port map (
            O => \N__39374\,
            I => \N__39370\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39367\
        );

    \I__8425\ : Span4Mux_h
    port map (
            O => \N__39370\,
            I => \N__39359\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39367\,
            I => \N__39356\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39353\
        );

    \I__8422\ : InMux
    port map (
            O => \N__39365\,
            I => \N__39348\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39348\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39345\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39362\,
            I => \N__39340\
        );

    \I__8418\ : Span4Mux_h
    port map (
            O => \N__39359\,
            I => \N__39335\
        );

    \I__8417\ : Span4Mux_v
    port map (
            O => \N__39356\,
            I => \N__39335\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39353\,
            I => \N__39331\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39348\,
            I => \N__39328\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39345\,
            I => \N__39325\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39322\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39319\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39340\,
            I => \N__39316\
        );

    \I__8410\ : Span4Mux_v
    port map (
            O => \N__39335\,
            I => \N__39313\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39310\
        );

    \I__8408\ : Span4Mux_v
    port map (
            O => \N__39331\,
            I => \N__39305\
        );

    \I__8407\ : Span4Mux_h
    port map (
            O => \N__39328\,
            I => \N__39305\
        );

    \I__8406\ : Span12Mux_s10_v
    port map (
            O => \N__39325\,
            I => \N__39302\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39322\,
            I => \N__39299\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__39319\,
            I => \N__39294\
        );

    \I__8403\ : Span4Mux_h
    port map (
            O => \N__39316\,
            I => \N__39294\
        );

    \I__8402\ : Sp12to4
    port map (
            O => \N__39313\,
            I => \N__39291\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39288\
        );

    \I__8400\ : Span4Mux_h
    port map (
            O => \N__39305\,
            I => \N__39285\
        );

    \I__8399\ : Span12Mux_v
    port map (
            O => \N__39302\,
            I => \N__39280\
        );

    \I__8398\ : Span4Mux_h
    port map (
            O => \N__39299\,
            I => \N__39277\
        );

    \I__8397\ : Span4Mux_h
    port map (
            O => \N__39294\,
            I => \N__39274\
        );

    \I__8396\ : Span12Mux_h
    port map (
            O => \N__39291\,
            I => \N__39267\
        );

    \I__8395\ : Span12Mux_s9_h
    port map (
            O => \N__39288\,
            I => \N__39267\
        );

    \I__8394\ : Sp12to4
    port map (
            O => \N__39285\,
            I => \N__39267\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39262\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39262\
        );

    \I__8391\ : Odrv12
    port map (
            O => \N__39280\,
            I => uart_pc_data_3
        );

    \I__8390\ : Odrv4
    port map (
            O => \N__39277\,
            I => uart_pc_data_3
        );

    \I__8389\ : Odrv4
    port map (
            O => \N__39274\,
            I => uart_pc_data_3
        );

    \I__8388\ : Odrv12
    port map (
            O => \N__39267\,
            I => uart_pc_data_3
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39262\,
            I => uart_pc_data_3
        );

    \I__8386\ : InMux
    port map (
            O => \N__39251\,
            I => \N__39247\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__39250\,
            I => \N__39243\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39247\,
            I => \N__39240\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39246\,
            I => \N__39237\
        );

    \I__8382\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39234\
        );

    \I__8381\ : Span4Mux_h
    port map (
            O => \N__39240\,
            I => \N__39231\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39237\,
            I => \N__39228\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__39234\,
            I => front_order_2
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__39231\,
            I => front_order_2
        );

    \I__8377\ : Odrv4
    port map (
            O => \N__39228\,
            I => front_order_2
        );

    \I__8376\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39218\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__39218\,
            I => \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\
        );

    \I__8374\ : CascadeMux
    port map (
            O => \N__39215\,
            I => \N__39211\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39208\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39211\,
            I => \N__39204\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39208\,
            I => \N__39201\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39198\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__39204\,
            I => \N__39193\
        );

    \I__8368\ : Span4Mux_h
    port map (
            O => \N__39201\,
            I => \N__39193\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__39198\,
            I => \N__39190\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__39193\,
            I => \ppm_encoder_1.elevatorZ0Z_2\
        );

    \I__8365\ : Odrv12
    port map (
            O => \N__39190\,
            I => \ppm_encoder_1.elevatorZ0Z_2\
        );

    \I__8364\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39182\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__39182\,
            I => \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\
        );

    \I__8362\ : CascadeMux
    port map (
            O => \N__39179\,
            I => \N__39176\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39176\,
            I => \N__39173\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39173\,
            I => \N__39168\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39172\,
            I => \N__39165\
        );

    \I__8358\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39162\
        );

    \I__8357\ : Span4Mux_h
    port map (
            O => \N__39168\,
            I => \N__39157\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39165\,
            I => \N__39157\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39162\,
            I => front_order_6
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__39157\,
            I => front_order_6
        );

    \I__8353\ : InMux
    port map (
            O => \N__39152\,
            I => \N__39149\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39145\
        );

    \I__8351\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39141\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__39145\,
            I => \N__39138\
        );

    \I__8349\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39135\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__39141\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__8347\ : Odrv4
    port map (
            O => \N__39138\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39135\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__8345\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39124\
        );

    \I__8344\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39121\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39118\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__39121\,
            I => \N__39115\
        );

    \I__8341\ : Span4Mux_v
    port map (
            O => \N__39118\,
            I => \N__39112\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__39115\,
            I => \N__39109\
        );

    \I__8339\ : Odrv4
    port map (
            O => \N__39112\,
            I => front_order_5
        );

    \I__8338\ : Odrv4
    port map (
            O => \N__39109\,
            I => front_order_5
        );

    \I__8337\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39101\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__39101\,
            I => \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\
        );

    \I__8335\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39094\
        );

    \I__8334\ : CascadeMux
    port map (
            O => \N__39097\,
            I => \N__39091\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39094\,
            I => \N__39088\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39084\
        );

    \I__8331\ : Span4Mux_h
    port map (
            O => \N__39088\,
            I => \N__39081\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39078\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__39084\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__39081\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__39078\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39068\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__39068\,
            I => \N__39064\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39067\,
            I => \N__39061\
        );

    \I__8323\ : Span4Mux_v
    port map (
            O => \N__39064\,
            I => \N__39058\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39061\,
            I => \N__39055\
        );

    \I__8321\ : Span4Mux_h
    port map (
            O => \N__39058\,
            I => \N__39052\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__39055\,
            I => \N__39049\
        );

    \I__8319\ : Span4Mux_h
    port map (
            O => \N__39052\,
            I => \N__39046\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__39049\,
            I => \N__39043\
        );

    \I__8317\ : Span4Mux_h
    port map (
            O => \N__39046\,
            I => \N__39040\
        );

    \I__8316\ : Span4Mux_h
    port map (
            O => \N__39043\,
            I => \N__39037\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__39040\,
            I => xy_kp_5
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__39037\,
            I => xy_kp_5
        );

    \I__8313\ : CEMux
    port map (
            O => \N__39032\,
            I => \N__39028\
        );

    \I__8312\ : CEMux
    port map (
            O => \N__39031\,
            I => \N__39023\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__39028\,
            I => \N__39020\
        );

    \I__8310\ : CEMux
    port map (
            O => \N__39027\,
            I => \N__39017\
        );

    \I__8309\ : CEMux
    port map (
            O => \N__39026\,
            I => \N__39014\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__39023\,
            I => \N__39011\
        );

    \I__8307\ : Span4Mux_v
    port map (
            O => \N__39020\,
            I => \N__39008\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39017\,
            I => \N__39005\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__39014\,
            I => \N__39002\
        );

    \I__8304\ : Span4Mux_h
    port map (
            O => \N__39011\,
            I => \N__38999\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__39008\,
            I => \N__38994\
        );

    \I__8302\ : Span4Mux_v
    port map (
            O => \N__39005\,
            I => \N__38994\
        );

    \I__8301\ : Span4Mux_h
    port map (
            O => \N__39002\,
            I => \N__38991\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__38999\,
            I => \N__38988\
        );

    \I__8299\ : Span4Mux_h
    port map (
            O => \N__38994\,
            I => \N__38985\
        );

    \I__8298\ : Span4Mux_v
    port map (
            O => \N__38991\,
            I => \N__38982\
        );

    \I__8297\ : Odrv4
    port map (
            O => \N__38988\,
            I => \Commands_frame_decoder.state_RNIG48SZ0Z_7\
        );

    \I__8296\ : Odrv4
    port map (
            O => \N__38985\,
            I => \Commands_frame_decoder.state_RNIG48SZ0Z_7\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__38982\,
            I => \Commands_frame_decoder.state_RNIG48SZ0Z_7\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__38975\,
            I => \N__38970\
        );

    \I__8293\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38967\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38962\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38970\,
            I => \N__38962\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38967\,
            I => \N__38956\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38956\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38952\
        );

    \I__8287\ : Span4Mux_h
    port map (
            O => \N__38956\,
            I => \N__38949\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38955\,
            I => \N__38946\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__38952\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__8284\ : Odrv4
    port map (
            O => \N__38949\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__38946\,
            I => \pid_front.pid_preregZ0Z_4\
        );

    \I__8282\ : InMux
    port map (
            O => \N__38939\,
            I => \N__38931\
        );

    \I__8281\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38931\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38926\
        );

    \I__8279\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38926\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__38931\,
            I => \N__38919\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38919\
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__38925\,
            I => \N__38916\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38913\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__38919\,
            I => \N__38910\
        );

    \I__8273\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38907\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__38913\,
            I => \pid_front.pid_preregZ0Z_5\
        );

    \I__8271\ : Odrv4
    port map (
            O => \N__38910\,
            I => \pid_front.pid_preregZ0Z_5\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38907\,
            I => \pid_front.pid_preregZ0Z_5\
        );

    \I__8269\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38896\
        );

    \I__8268\ : InMux
    port map (
            O => \N__38899\,
            I => \N__38893\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__38896\,
            I => \N__38887\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38887\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38883\
        );

    \I__8264\ : Span4Mux_v
    port map (
            O => \N__38887\,
            I => \N__38880\
        );

    \I__8263\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38877\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__38883\,
            I => \pid_front.pid_preregZ0Z_3\
        );

    \I__8261\ : Odrv4
    port map (
            O => \N__38880\,
            I => \pid_front.pid_preregZ0Z_3\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38877\,
            I => \pid_front.pid_preregZ0Z_3\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38867\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38867\,
            I => \N__38864\
        );

    \I__8257\ : Span12Mux_v
    port map (
            O => \N__38864\,
            I => \N__38861\
        );

    \I__8256\ : Span12Mux_h
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__8255\ : Odrv12
    port map (
            O => \N__38858\,
            I => alt_ki_6
        );

    \I__8254\ : CEMux
    port map (
            O => \N__38855\,
            I => \N__38852\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__38852\,
            I => \N__38849\
        );

    \I__8252\ : Span4Mux_h
    port map (
            O => \N__38849\,
            I => \N__38845\
        );

    \I__8251\ : CEMux
    port map (
            O => \N__38848\,
            I => \N__38842\
        );

    \I__8250\ : Span4Mux_h
    port map (
            O => \N__38845\,
            I => \N__38836\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38842\,
            I => \N__38836\
        );

    \I__8248\ : CEMux
    port map (
            O => \N__38841\,
            I => \N__38833\
        );

    \I__8247\ : Span4Mux_h
    port map (
            O => \N__38836\,
            I => \N__38829\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38833\,
            I => \N__38826\
        );

    \I__8245\ : CEMux
    port map (
            O => \N__38832\,
            I => \N__38823\
        );

    \I__8244\ : Span4Mux_v
    port map (
            O => \N__38829\,
            I => \N__38820\
        );

    \I__8243\ : Span4Mux_v
    port map (
            O => \N__38826\,
            I => \N__38815\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__38823\,
            I => \N__38815\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__38820\,
            I => \N__38810\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__38815\,
            I => \N__38810\
        );

    \I__8239\ : Odrv4
    port map (
            O => \N__38810\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38803\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38806\,
            I => \N__38799\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__38803\,
            I => \N__38796\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38793\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38790\
        );

    \I__8233\ : Span4Mux_v
    port map (
            O => \N__38796\,
            I => \N__38787\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38793\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__38790\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__8230\ : Odrv4
    port map (
            O => \N__38787\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38777\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38777\,
            I => \N__38772\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38776\,
            I => \N__38769\
        );

    \I__8226\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38766\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__38772\,
            I => \N__38763\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__38769\,
            I => \N__38760\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38753\
        );

    \I__8222\ : Span4Mux_v
    port map (
            O => \N__38763\,
            I => \N__38753\
        );

    \I__8221\ : Span4Mux_h
    port map (
            O => \N__38760\,
            I => \N__38753\
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__38753\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38750\,
            I => \N__38747\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__38744\,
            I => \N__38740\
        );

    \I__8216\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38737\
        );

    \I__8215\ : Span4Mux_v
    port map (
            O => \N__38740\,
            I => \N__38734\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__38737\,
            I => \N__38731\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__38734\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__8212\ : Odrv4
    port map (
            O => \N__38731\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__8211\ : CascadeMux
    port map (
            O => \N__38726\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__38723\,
            I => \N__38720\
        );

    \I__8209\ : InMux
    port map (
            O => \N__38720\,
            I => \N__38717\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__38717\,
            I => \N__38714\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__38711\,
            I => \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\
        );

    \I__8205\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__38705\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6\
        );

    \I__8203\ : CascadeMux
    port map (
            O => \N__38702\,
            I => \N__38699\
        );

    \I__8202\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38694\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__38698\,
            I => \N__38691\
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__38697\,
            I => \N__38688\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38685\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38682\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38679\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__38685\,
            I => \N__38674\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__38682\,
            I => \N__38674\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38679\,
            I => side_order_6
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__38674\,
            I => side_order_6
        );

    \I__8192\ : InMux
    port map (
            O => \N__38669\,
            I => \N__38666\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38666\,
            I => \N__38663\
        );

    \I__8190\ : Span4Mux_v
    port map (
            O => \N__38663\,
            I => \N__38660\
        );

    \I__8189\ : Odrv4
    port map (
            O => \N__38660\,
            I => \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38649\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__38653\,
            I => \N__38646\
        );

    \I__8185\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38643\
        );

    \I__8184\ : Span4Mux_h
    port map (
            O => \N__38649\,
            I => \N__38640\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38646\,
            I => \N__38637\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38643\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__38640\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__38637\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38624\
        );

    \I__8177\ : Span4Mux_h
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8176\ : Span4Mux_v
    port map (
            O => \N__38621\,
            I => \N__38618\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__38618\,
            I => \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38615\,
            I => \N__38610\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38614\,
            I => \N__38607\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38604\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38610\,
            I => \N__38601\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38607\,
            I => side_order_3
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__38604\,
            I => side_order_3
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__38601\,
            I => side_order_3
        );

    \I__8167\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38591\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38588\
        );

    \I__8165\ : Span4Mux_h
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__8164\ : Span4Mux_v
    port map (
            O => \N__38585\,
            I => \N__38582\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38582\,
            I => \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38575\
        );

    \I__8161\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38572\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__38575\,
            I => \N__38569\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38572\,
            I => \N__38566\
        );

    \I__8158\ : Span4Mux_v
    port map (
            O => \N__38569\,
            I => \N__38563\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38566\,
            I => side_order_5
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__38563\,
            I => side_order_5
        );

    \I__8155\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38555\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38555\,
            I => \N__38551\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38554\,
            I => \N__38547\
        );

    \I__8152\ : Span4Mux_h
    port map (
            O => \N__38551\,
            I => \N__38544\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__38550\,
            I => \N__38541\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38547\,
            I => \N__38538\
        );

    \I__8149\ : Span4Mux_h
    port map (
            O => \N__38544\,
            I => \N__38535\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38541\,
            I => \N__38532\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38538\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__38535\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__38532\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38521\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__38524\,
            I => \N__38518\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38515\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38511\
        );

    \I__8140\ : Span4Mux_h
    port map (
            O => \N__38515\,
            I => \N__38508\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38505\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38511\,
            I => side_order_9
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__38508\,
            I => side_order_9
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__38505\,
            I => side_order_9
        );

    \I__8135\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38492\
        );

    \I__8133\ : Span4Mux_v
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38489\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38480\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38480\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38480\,
            I => \N__38476\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__8127\ : Span4Mux_h
    port map (
            O => \N__38476\,
            I => \N__38470\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38473\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__38470\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__38465\,
            I => \N__38461\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38457\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38454\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38451\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38457\,
            I => \N__38448\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38454\,
            I => \N__38443\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38451\,
            I => \N__38443\
        );

    \I__8117\ : Span4Mux_v
    port map (
            O => \N__38448\,
            I => \N__38440\
        );

    \I__8116\ : Odrv12
    port map (
            O => \N__38443\,
            I => front_order_10
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__38440\,
            I => front_order_10
        );

    \I__8114\ : InMux
    port map (
            O => \N__38435\,
            I => \N__38432\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38432\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38425\
        );

    \I__8111\ : CascadeMux
    port map (
            O => \N__38428\,
            I => \N__38421\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__38425\,
            I => \N__38418\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38415\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38421\,
            I => \N__38412\
        );

    \I__8107\ : Span4Mux_v
    port map (
            O => \N__38418\,
            I => \N__38409\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__38415\,
            I => \N__38406\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38412\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__38409\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__38406\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38393\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38393\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38390\
        );

    \I__8099\ : Span4Mux_v
    port map (
            O => \N__38390\,
            I => \N__38385\
        );

    \I__8098\ : InMux
    port map (
            O => \N__38389\,
            I => \N__38380\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38380\
        );

    \I__8096\ : Odrv4
    port map (
            O => \N__38385\,
            I => \pid_side.N_563\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__38380\,
            I => \pid_side.N_563\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38372\,
            I => \N__38365\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38365\
        );

    \I__8091\ : CascadeMux
    port map (
            O => \N__38370\,
            I => \N__38362\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38365\,
            I => \N__38357\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38362\,
            I => \N__38354\
        );

    \I__8088\ : InMux
    port map (
            O => \N__38361\,
            I => \N__38351\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38348\
        );

    \I__8086\ : Span4Mux_v
    port map (
            O => \N__38357\,
            I => \N__38345\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38354\,
            I => \N__38340\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38351\,
            I => \N__38340\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__38348\,
            I => \N__38337\
        );

    \I__8082\ : Span4Mux_h
    port map (
            O => \N__38345\,
            I => \N__38332\
        );

    \I__8081\ : Span4Mux_h
    port map (
            O => \N__38340\,
            I => \N__38332\
        );

    \I__8080\ : Span4Mux_h
    port map (
            O => \N__38337\,
            I => \N__38329\
        );

    \I__8079\ : Span4Mux_h
    port map (
            O => \N__38332\,
            I => \N__38326\
        );

    \I__8078\ : Span4Mux_h
    port map (
            O => \N__38329\,
            I => \N__38323\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__38326\,
            I => \pid_side.pid_preregZ0Z_21\
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__38323\,
            I => \pid_side.pid_preregZ0Z_21\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38309\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38309\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38306\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38303\
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__38314\,
            I => \N__38299\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__38309\,
            I => \N__38296\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__38306\,
            I => \N__38293\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__38303\,
            I => \N__38290\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38285\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38285\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__38296\,
            I => \N__38281\
        );

    \I__8064\ : Span4Mux_h
    port map (
            O => \N__38293\,
            I => \N__38274\
        );

    \I__8063\ : Span4Mux_v
    port map (
            O => \N__38290\,
            I => \N__38274\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38274\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38271\
        );

    \I__8060\ : Span4Mux_h
    port map (
            O => \N__38281\,
            I => \N__38268\
        );

    \I__8059\ : Span4Mux_h
    port map (
            O => \N__38274\,
            I => \N__38265\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__38271\,
            I => \pid_side.pid_preregZ0Z_13\
        );

    \I__8057\ : Odrv4
    port map (
            O => \N__38268\,
            I => \pid_side.pid_preregZ0Z_13\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__38265\,
            I => \pid_side.pid_preregZ0Z_13\
        );

    \I__8055\ : CascadeMux
    port map (
            O => \N__38258\,
            I => \N__38253\
        );

    \I__8054\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38250\
        );

    \I__8053\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38247\
        );

    \I__8052\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38243\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__38250\,
            I => \N__38240\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__38247\,
            I => \N__38237\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38234\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__38243\,
            I => \N__38231\
        );

    \I__8047\ : Span4Mux_h
    port map (
            O => \N__38240\,
            I => \N__38227\
        );

    \I__8046\ : Span4Mux_h
    port map (
            O => \N__38237\,
            I => \N__38224\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__38234\,
            I => \N__38219\
        );

    \I__8044\ : Span4Mux_v
    port map (
            O => \N__38231\,
            I => \N__38219\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38216\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__38227\,
            I => \N__38213\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__38224\,
            I => \N__38208\
        );

    \I__8040\ : Span4Mux_h
    port map (
            O => \N__38219\,
            I => \N__38208\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__38216\,
            I => \pid_side.pid_preregZ0Z_4\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__38213\,
            I => \pid_side.pid_preregZ0Z_4\
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__38208\,
            I => \pid_side.pid_preregZ0Z_4\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38195\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38195\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38192\
        );

    \I__8033\ : Span4Mux_h
    port map (
            O => \N__38192\,
            I => \N__38188\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__38188\,
            I => \pid_side.N_534\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__38185\,
            I => \pid_side.N_534\
        );

    \I__8029\ : CascadeMux
    port map (
            O => \N__38180\,
            I => \N__38176\
        );

    \I__8028\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38165\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38165\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38152\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38152\
        );

    \I__8024\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38152\
        );

    \I__8023\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38152\
        );

    \I__8022\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38152\
        );

    \I__8021\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38152\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__38165\,
            I => \pid_side.N_291\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38152\,
            I => \pid_side.N_291\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__38147\,
            I => \N__38144\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38139\
        );

    \I__8016\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38133\
        );

    \I__8015\ : InMux
    port map (
            O => \N__38142\,
            I => \N__38133\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__38139\,
            I => \N__38130\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38127\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__38133\,
            I => \N__38124\
        );

    \I__8011\ : Span4Mux_v
    port map (
            O => \N__38130\,
            I => \N__38118\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38118\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__38124\,
            I => \N__38114\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38111\
        );

    \I__8007\ : Span4Mux_h
    port map (
            O => \N__38118\,
            I => \N__38108\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38105\
        );

    \I__8005\ : Sp12to4
    port map (
            O => \N__38114\,
            I => \N__38100\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__38111\,
            I => \N__38100\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__38108\,
            I => \N__38097\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38105\,
            I => \pid_side.pid_preregZ0Z_5\
        );

    \I__8001\ : Odrv12
    port map (
            O => \N__38100\,
            I => \pid_side.pid_preregZ0Z_5\
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__38097\,
            I => \pid_side.pid_preregZ0Z_5\
        );

    \I__7999\ : CEMux
    port map (
            O => \N__38090\,
            I => \N__38087\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__38087\,
            I => \N__38084\
        );

    \I__7997\ : Span4Mux_h
    port map (
            O => \N__38084\,
            I => \N__38081\
        );

    \I__7996\ : Span4Mux_v
    port map (
            O => \N__38081\,
            I => \N__38078\
        );

    \I__7995\ : Odrv4
    port map (
            O => \N__38078\,
            I => \pid_side.state_0_1\
        );

    \I__7994\ : SRMux
    port map (
            O => \N__38075\,
            I => \N__38070\
        );

    \I__7993\ : SRMux
    port map (
            O => \N__38074\,
            I => \N__38067\
        );

    \I__7992\ : SRMux
    port map (
            O => \N__38073\,
            I => \N__38064\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38070\,
            I => \N__38061\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__38067\,
            I => \N__38057\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38064\,
            I => \N__38054\
        );

    \I__7988\ : Span4Mux_h
    port map (
            O => \N__38061\,
            I => \N__38051\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38060\,
            I => \N__38048\
        );

    \I__7986\ : Odrv4
    port map (
            O => \N__38057\,
            I => \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__38054\,
            I => \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\
        );

    \I__7984\ : Odrv4
    port map (
            O => \N__38051\,
            I => \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__38048\,
            I => \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\
        );

    \I__7982\ : CascadeMux
    port map (
            O => \N__38039\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\
        );

    \I__7981\ : CascadeMux
    port map (
            O => \N__38036\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\
        );

    \I__7980\ : CascadeMux
    port map (
            O => \N__38033\,
            I => \N__38030\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38027\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38027\,
            I => \N__38024\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__38024\,
            I => \N__38021\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__38021\,
            I => \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38018\,
            I => \N__38013\
        );

    \I__7974\ : CascadeMux
    port map (
            O => \N__38017\,
            I => \N__38010\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38016\,
            I => \N__38007\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__38004\
        );

    \I__7971\ : InMux
    port map (
            O => \N__38010\,
            I => \N__38001\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__38007\,
            I => \N__37996\
        );

    \I__7969\ : Span4Mux_h
    port map (
            O => \N__38004\,
            I => \N__37996\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__38001\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__37996\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__7966\ : CascadeMux
    port map (
            O => \N__37991\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37985\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__37985\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5\
        );

    \I__7963\ : CascadeMux
    port map (
            O => \N__37982\,
            I => \N__37979\
        );

    \I__7962\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37976\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__37976\,
            I => \N__37973\
        );

    \I__7960\ : Span4Mux_v
    port map (
            O => \N__37973\,
            I => \N__37970\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__37970\,
            I => \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37960\
        );

    \I__7957\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37960\
        );

    \I__7956\ : InMux
    port map (
            O => \N__37965\,
            I => \N__37957\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__37960\,
            I => \ppm_encoder_1.aileronZ0Z_1\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__37957\,
            I => \ppm_encoder_1.aileronZ0Z_1\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__37952\,
            I => \N__37948\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__37951\,
            I => \N__37944\
        );

    \I__7951\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37941\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37938\
        );

    \I__7949\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37935\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__37941\,
            I => \ppm_encoder_1.elevatorZ0Z_1\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__37938\,
            I => \ppm_encoder_1.elevatorZ0Z_1\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__37935\,
            I => \ppm_encoder_1.elevatorZ0Z_1\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__37928\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__7944\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37922\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__37922\,
            I => \N__37918\
        );

    \I__7942\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37915\
        );

    \I__7941\ : Odrv12
    port map (
            O => \N__37918\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37915\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__37910\,
            I => \N__37907\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__37904\,
            I => \N__37901\
        );

    \I__7936\ : Span4Mux_h
    port map (
            O => \N__37901\,
            I => \N__37898\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__37898\,
            I => \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37890\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37894\,
            I => \N__37887\
        );

    \I__7932\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37884\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__37890\,
            I => \N__37881\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37887\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__37884\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__37881\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__37874\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37871\,
            I => \N__37868\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__37868\,
            I => \ppm_encoder_1.throttle_m_1\
        );

    \I__7924\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37859\
        );

    \I__7923\ : InMux
    port map (
            O => \N__37864\,
            I => \N__37859\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__37859\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37852\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37849\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__37852\,
            I => \N__37844\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__37849\,
            I => \N__37844\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__37844\,
            I => \N__37838\
        );

    \I__7916\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37833\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37833\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37830\
        );

    \I__7913\ : Sp12to4
    port map (
            O => \N__37838\,
            I => \N__37825\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__37833\,
            I => \N__37825\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__37830\,
            I => \pid_side.pid_preregZ0Z_12\
        );

    \I__7910\ : Odrv12
    port map (
            O => \N__37825\,
            I => \pid_side.pid_preregZ0Z_12\
        );

    \I__7909\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37816\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37813\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37810\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37807\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__37810\,
            I => \N__37802\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__37807\,
            I => \N__37802\
        );

    \I__7903\ : Odrv4
    port map (
            O => \N__37802\,
            I => side_order_12
        );

    \I__7902\ : InMux
    port map (
            O => \N__37799\,
            I => \N__37796\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__37796\,
            I => \N__37791\
        );

    \I__7900\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37788\
        );

    \I__7899\ : CascadeMux
    port map (
            O => \N__37794\,
            I => \N__37785\
        );

    \I__7898\ : Span4Mux_h
    port map (
            O => \N__37791\,
            I => \N__37780\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__37788\,
            I => \N__37780\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37777\
        );

    \I__7895\ : Span4Mux_h
    port map (
            O => \N__37780\,
            I => \N__37774\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37777\,
            I => throttle_order_8
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__37774\,
            I => throttle_order_8
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__37769\,
            I => \N__37766\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37763\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37760\
        );

    \I__7889\ : Odrv12
    port map (
            O => \N__37760\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__7888\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37748\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37748\
        );

    \I__7886\ : InMux
    port map (
            O => \N__37755\,
            I => \N__37748\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__37748\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__37745\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\
        );

    \I__7883\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37738\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37734\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37738\,
            I => \N__37731\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37737\,
            I => \N__37728\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37723\
        );

    \I__7878\ : Span4Mux_h
    port map (
            O => \N__37731\,
            I => \N__37723\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37728\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__37723\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__7875\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37715\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__37715\,
            I => \N__37711\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37707\
        );

    \I__7872\ : Span4Mux_h
    port map (
            O => \N__37711\,
            I => \N__37704\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37710\,
            I => \N__37701\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__37707\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__37704\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37701\,
            I => \ppm_encoder_1.aileronZ0Z_2\
        );

    \I__7867\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37688\
        );

    \I__7865\ : Span12Mux_v
    port map (
            O => \N__37688\,
            I => \N__37684\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37681\
        );

    \I__7863\ : Odrv12
    port map (
            O => \N__37684\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__37681\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__7861\ : CascadeMux
    port map (
            O => \N__37676\,
            I => \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\
        );

    \I__7860\ : CascadeMux
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__7859\ : InMux
    port map (
            O => \N__37670\,
            I => \N__37667\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__37667\,
            I => \N__37664\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__37664\,
            I => \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__37658\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__7853\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37649\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__37649\,
            I => \N__37646\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__37646\,
            I => \N__37643\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__37643\,
            I => \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37640\,
            I => \N__37637\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37634\
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__37634\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__37631\,
            I => \N__37628\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37625\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__37625\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37619\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7841\ : Odrv12
    port map (
            O => \N__37616\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__37613\,
            I => \N__37610\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37607\,
            I => \N__37602\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37606\,
            I => \N__37599\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__37605\,
            I => \N__37596\
        );

    \I__7835\ : Span4Mux_h
    port map (
            O => \N__37602\,
            I => \N__37593\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37599\,
            I => \N__37590\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37587\
        );

    \I__7832\ : Span4Mux_v
    port map (
            O => \N__37593\,
            I => \N__37584\
        );

    \I__7831\ : Span4Mux_h
    port map (
            O => \N__37590\,
            I => \N__37581\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__37587\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__37584\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__37581\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__7827\ : CascadeMux
    port map (
            O => \N__37574\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__37571\,
            I => \N__37568\
        );

    \I__7825\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37565\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__37565\,
            I => \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37559\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37559\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__37556\,
            I => \ppm_encoder_1.N_294_cascade_\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37549\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__37552\,
            I => \N__37546\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__37549\,
            I => \N__37543\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37546\,
            I => \N__37539\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__37543\,
            I => \N__37536\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37542\,
            I => \N__37533\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37539\,
            I => side_order_8
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__37536\,
            I => side_order_8
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__37533\,
            I => side_order_8
        );

    \I__7811\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37517\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37505\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37505\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37505\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37505\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__37499\,
            I => \N__37495\
        );

    \I__7801\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37492\
        );

    \I__7800\ : Span4Mux_v
    port map (
            O => \N__37495\,
            I => \N__37488\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37485\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37491\,
            I => \N__37482\
        );

    \I__7797\ : Span4Mux_h
    port map (
            O => \N__37488\,
            I => \N__37477\
        );

    \I__7796\ : Span4Mux_h
    port map (
            O => \N__37485\,
            I => \N__37477\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37482\,
            I => front_order_8
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__37477\,
            I => front_order_8
        );

    \I__7793\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__37463\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37460\,
            I => \N__37455\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37459\,
            I => \N__37450\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37450\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37455\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__37450\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__37442\,
            I => \N__37437\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37432\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37432\
        );

    \I__7780\ : Span4Mux_v
    port map (
            O => \N__37437\,
            I => \N__37429\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37432\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__7778\ : Odrv4
    port map (
            O => \N__37429\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37421\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__37421\,
            I => \N__37418\
        );

    \I__7775\ : Odrv4
    port map (
            O => \N__37418\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37415\,
            I => \N__37412\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__37412\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37406\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37400\,
            I => \N__37397\
        );

    \I__7768\ : Odrv12
    port map (
            O => \N__37397\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37391\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__7763\ : Span4Mux_h
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__37379\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__37373\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__37370\,
            I => \N__37367\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37364\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__7756\ : CascadeMux
    port map (
            O => \N__37361\,
            I => \N__37358\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__37352\,
            I => \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\
        );

    \I__7752\ : CascadeMux
    port map (
            O => \N__37349\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\
        );

    \I__7751\ : CascadeMux
    port map (
            O => \N__37346\,
            I => \N__37343\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37340\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__37337\,
            I => \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7745\ : Odrv4
    port map (
            O => \N__37328\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37322\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__37322\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37316\
        );

    \I__7741\ : LocalMux
    port map (
            O => \N__37316\,
            I => \N__37313\
        );

    \I__7740\ : Odrv4
    port map (
            O => \N__37313\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__7739\ : InMux
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37307\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__7737\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37298\
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__37298\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37295\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__37289\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__7730\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__37280\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__7728\ : InMux
    port map (
            O => \N__37277\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__7726\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37268\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37268\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__7724\ : InMux
    port map (
            O => \N__37265\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__7723\ : InMux
    port map (
            O => \N__37262\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__7722\ : InMux
    port map (
            O => \N__37259\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37256\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37253\,
            I => \N__37250\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37250\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__37244\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__7716\ : InMux
    port map (
            O => \N__37241\,
            I => \bfn_16_10_0_\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37235\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__7713\ : InMux
    port map (
            O => \N__37232\,
            I => \N__37229\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37229\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__7711\ : InMux
    port map (
            O => \N__37226\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__7710\ : InMux
    port map (
            O => \N__37223\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__7709\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__37217\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7706\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37208\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__37208\,
            I => \N__37205\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__37205\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37202\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__7702\ : InMux
    port map (
            O => \N__37199\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__7701\ : InMux
    port map (
            O => \N__37196\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37193\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__7699\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__7697\ : Span4Mux_h
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__37181\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__7695\ : InMux
    port map (
            O => \N__37178\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__7694\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37172\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__7692\ : Span4Mux_h
    port map (
            O => \N__37169\,
            I => \N__37166\
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__37166\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7688\ : Span4Mux_h
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__37154\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37151\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37145\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7682\ : Odrv4
    port map (
            O => \N__37139\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37136\,
            I => \bfn_16_9_0_\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37133\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37125\
        );

    \I__7678\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37122\
        );

    \I__7677\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37119\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37125\,
            I => \N__37115\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__37122\,
            I => \N__37109\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37119\,
            I => \N__37106\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37103\
        );

    \I__7672\ : Span4Mux_h
    port map (
            O => \N__37115\,
            I => \N__37100\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37114\,
            I => \N__37097\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37094\
        );

    \I__7669\ : InMux
    port map (
            O => \N__37112\,
            I => \N__37091\
        );

    \I__7668\ : Span12Mux_h
    port map (
            O => \N__37109\,
            I => \N__37084\
        );

    \I__7667\ : Sp12to4
    port map (
            O => \N__37106\,
            I => \N__37084\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37084\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__37100\,
            I => \N__37081\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37097\,
            I => \N__37078\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__37094\,
            I => \N__37075\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__37091\,
            I => \N__37072\
        );

    \I__7661\ : Span12Mux_v
    port map (
            O => \N__37084\,
            I => \N__37069\
        );

    \I__7660\ : Sp12to4
    port map (
            O => \N__37081\,
            I => \N__37062\
        );

    \I__7659\ : Span12Mux_s10_h
    port map (
            O => \N__37078\,
            I => \N__37062\
        );

    \I__7658\ : Sp12to4
    port map (
            O => \N__37075\,
            I => \N__37062\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__37072\,
            I => \N__37059\
        );

    \I__7656\ : Odrv12
    port map (
            O => \N__37069\,
            I => uart_drone_data_2
        );

    \I__7655\ : Odrv12
    port map (
            O => \N__37062\,
            I => uart_drone_data_2
        );

    \I__7654\ : Odrv4
    port map (
            O => \N__37059\,
            I => uart_drone_data_2
        );

    \I__7653\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37049\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__37045\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37041\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__37045\,
            I => \N__37038\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37044\,
            I => \N__37035\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__37041\,
            I => \N__37031\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__37038\,
            I => \N__37026\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__37035\,
            I => \N__37026\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37023\
        );

    \I__7644\ : Span4Mux_v
    port map (
            O => \N__37031\,
            I => \N__37019\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__37026\,
            I => \N__37014\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__37023\,
            I => \N__37014\
        );

    \I__7641\ : InMux
    port map (
            O => \N__37022\,
            I => \N__37011\
        );

    \I__7640\ : Sp12to4
    port map (
            O => \N__37019\,
            I => \N__37006\
        );

    \I__7639\ : Span4Mux_h
    port map (
            O => \N__37014\,
            I => \N__37003\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37011\,
            I => \N__37000\
        );

    \I__7637\ : InMux
    port map (
            O => \N__37010\,
            I => \N__36997\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37009\,
            I => \N__36993\
        );

    \I__7635\ : Span12Mux_h
    port map (
            O => \N__37006\,
            I => \N__36984\
        );

    \I__7634\ : Sp12to4
    port map (
            O => \N__37003\,
            I => \N__36984\
        );

    \I__7633\ : Sp12to4
    port map (
            O => \N__37000\,
            I => \N__36984\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__36997\,
            I => \N__36984\
        );

    \I__7631\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36981\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36978\
        );

    \I__7629\ : Odrv12
    port map (
            O => \N__36984\,
            I => uart_drone_data_3
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__36981\,
            I => uart_drone_data_3
        );

    \I__7627\ : Odrv4
    port map (
            O => \N__36978\,
            I => uart_drone_data_3
        );

    \I__7626\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36966\
        );

    \I__7625\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36963\
        );

    \I__7624\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36960\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__36966\,
            I => \N__36956\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__36963\,
            I => \N__36953\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36960\,
            I => \N__36950\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36947\
        );

    \I__7619\ : Span4Mux_v
    port map (
            O => \N__36956\,
            I => \N__36943\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__36953\,
            I => \N__36940\
        );

    \I__7617\ : Span4Mux_v
    port map (
            O => \N__36950\,
            I => \N__36935\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__36947\,
            I => \N__36935\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36946\,
            I => \N__36931\
        );

    \I__7614\ : Sp12to4
    port map (
            O => \N__36943\,
            I => \N__36928\
        );

    \I__7613\ : Span4Mux_h
    port map (
            O => \N__36940\,
            I => \N__36923\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__36935\,
            I => \N__36923\
        );

    \I__7611\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36920\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__36931\,
            I => \N__36916\
        );

    \I__7609\ : Span12Mux_h
    port map (
            O => \N__36928\,
            I => \N__36909\
        );

    \I__7608\ : Sp12to4
    port map (
            O => \N__36923\,
            I => \N__36909\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__36920\,
            I => \N__36909\
        );

    \I__7606\ : InMux
    port map (
            O => \N__36919\,
            I => \N__36905\
        );

    \I__7605\ : Span12Mux_v
    port map (
            O => \N__36916\,
            I => \N__36902\
        );

    \I__7604\ : Span12Mux_v
    port map (
            O => \N__36909\,
            I => \N__36899\
        );

    \I__7603\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36896\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36893\
        );

    \I__7601\ : Odrv12
    port map (
            O => \N__36902\,
            I => uart_drone_data_4
        );

    \I__7600\ : Odrv12
    port map (
            O => \N__36899\,
            I => uart_drone_data_4
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__36896\,
            I => uart_drone_data_4
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__36893\,
            I => uart_drone_data_4
        );

    \I__7597\ : InMux
    port map (
            O => \N__36884\,
            I => \N__36881\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36874\
        );

    \I__7595\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36871\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36868\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36865\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36862\
        );

    \I__7591\ : Span4Mux_v
    port map (
            O => \N__36874\,
            I => \N__36857\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36857\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36852\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36852\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36849\
        );

    \I__7586\ : Span4Mux_v
    port map (
            O => \N__36857\,
            I => \N__36845\
        );

    \I__7585\ : Span4Mux_v
    port map (
            O => \N__36852\,
            I => \N__36841\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__36849\,
            I => \N__36838\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36835\
        );

    \I__7582\ : Sp12to4
    port map (
            O => \N__36845\,
            I => \N__36832\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36829\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__36841\,
            I => \N__36822\
        );

    \I__7579\ : Span4Mux_v
    port map (
            O => \N__36838\,
            I => \N__36822\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36835\,
            I => \N__36822\
        );

    \I__7577\ : Span12Mux_h
    port map (
            O => \N__36832\,
            I => \N__36817\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__36829\,
            I => \N__36817\
        );

    \I__7575\ : Span4Mux_v
    port map (
            O => \N__36822\,
            I => \N__36814\
        );

    \I__7574\ : Odrv12
    port map (
            O => \N__36817\,
            I => uart_drone_data_5
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__36814\,
            I => uart_drone_data_5
        );

    \I__7572\ : InMux
    port map (
            O => \N__36809\,
            I => \N__36804\
        );

    \I__7571\ : InMux
    port map (
            O => \N__36808\,
            I => \N__36800\
        );

    \I__7570\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36797\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36793\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36790\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36784\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__36797\,
            I => \N__36784\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36796\,
            I => \N__36781\
        );

    \I__7564\ : Span4Mux_v
    port map (
            O => \N__36793\,
            I => \N__36778\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36790\,
            I => \N__36775\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36772\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__36784\,
            I => \N__36767\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36767\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__36778\,
            I => \N__36760\
        );

    \I__7558\ : Span4Mux_h
    port map (
            O => \N__36775\,
            I => \N__36760\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__36772\,
            I => \N__36760\
        );

    \I__7556\ : Span4Mux_v
    port map (
            O => \N__36767\,
            I => \N__36756\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__36760\,
            I => \N__36753\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36750\
        );

    \I__7553\ : Span4Mux_h
    port map (
            O => \N__36756\,
            I => \N__36746\
        );

    \I__7552\ : Span4Mux_v
    port map (
            O => \N__36753\,
            I => \N__36741\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36741\
        );

    \I__7550\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36738\
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__36746\,
            I => uart_drone_data_1
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__36741\,
            I => uart_drone_data_1
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__36738\,
            I => uart_drone_data_1
        );

    \I__7546\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36727\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__36730\,
            I => \N__36724\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__36727\,
            I => \N__36721\
        );

    \I__7543\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36718\
        );

    \I__7542\ : Odrv12
    port map (
            O => \N__36721\,
            I => scaler_4_data_4
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36718\,
            I => scaler_4_data_4
        );

    \I__7540\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__36710\,
            I => \N__36707\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__36704\,
            I => \N__36701\
        );

    \I__7536\ : Odrv4
    port map (
            O => \N__36701\,
            I => scaler_4_data_5
        );

    \I__7535\ : CEMux
    port map (
            O => \N__36698\,
            I => \N__36694\
        );

    \I__7534\ : CEMux
    port map (
            O => \N__36697\,
            I => \N__36689\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36694\,
            I => \N__36685\
        );

    \I__7532\ : CEMux
    port map (
            O => \N__36693\,
            I => \N__36682\
        );

    \I__7531\ : CEMux
    port map (
            O => \N__36692\,
            I => \N__36679\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36676\
        );

    \I__7529\ : CEMux
    port map (
            O => \N__36688\,
            I => \N__36673\
        );

    \I__7528\ : Span4Mux_v
    port map (
            O => \N__36685\,
            I => \N__36670\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__36682\,
            I => \N__36667\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36664\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__36676\,
            I => \N__36661\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36658\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__36670\,
            I => \N__36653\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__36667\,
            I => \N__36653\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__36664\,
            I => \N__36650\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__36661\,
            I => \N__36647\
        );

    \I__7519\ : Span12Mux_h
    port map (
            O => \N__36658\,
            I => \N__36644\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__36653\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7517\ : Odrv4
    port map (
            O => \N__36650\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__36647\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7515\ : Odrv12
    port map (
            O => \N__36644\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36635\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36629\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__36629\,
            I => \N__36624\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36628\,
            I => \N__36621\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36617\
        );

    \I__7509\ : Span4Mux_h
    port map (
            O => \N__36624\,
            I => \N__36613\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36621\,
            I => \N__36610\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36606\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36617\,
            I => \N__36602\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36599\
        );

    \I__7504\ : Span4Mux_h
    port map (
            O => \N__36613\,
            I => \N__36594\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__36610\,
            I => \N__36594\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36591\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__36606\,
            I => \N__36588\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36585\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__36602\,
            I => \N__36580\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36599\,
            I => \N__36580\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__36594\,
            I => \N__36575\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__36591\,
            I => \N__36575\
        );

    \I__7495\ : Sp12to4
    port map (
            O => \N__36588\,
            I => \N__36570\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36585\,
            I => \N__36570\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__36580\,
            I => \N__36567\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__36575\,
            I => \N__36564\
        );

    \I__7491\ : Span12Mux_v
    port map (
            O => \N__36570\,
            I => \N__36561\
        );

    \I__7490\ : Span4Mux_v
    port map (
            O => \N__36567\,
            I => \N__36558\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__36564\,
            I => \N__36555\
        );

    \I__7488\ : Odrv12
    port map (
            O => \N__36561\,
            I => uart_drone_data_7
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__36558\,
            I => uart_drone_data_7
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__36555\,
            I => uart_drone_data_7
        );

    \I__7485\ : CascadeMux
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36541\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36538\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__36541\,
            I => \pid_front.pid_preregZ0Z_17\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__36538\,
            I => \pid_front.pid_preregZ0Z_17\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36529\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36532\,
            I => \N__36526\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__36529\,
            I => \pid_front.pid_preregZ0Z_20\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36526\,
            I => \pid_front.pid_preregZ0Z_20\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__36521\,
            I => \N__36517\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36520\,
            I => \N__36511\
        );

    \I__7474\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36511\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__36516\,
            I => \N__36507\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36504\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36501\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36498\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__36504\,
            I => \N__36495\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__36501\,
            I => \N__36492\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36498\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__36495\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__36492\,
            I => \pid_front.pid_preregZ0Z_7\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36479\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36474\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36471\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36468\
        );

    \I__7459\ : Span4Mux_h
    port map (
            O => \N__36474\,
            I => \N__36465\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36471\,
            I => \N__36462\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__36468\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__36465\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__36462\,
            I => \pid_front.pid_preregZ0Z_6\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36449\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36454\,
            I => \N__36446\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36441\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36441\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__36449\,
            I => \N__36435\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36446\,
            I => \N__36435\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36441\,
            I => \N__36432\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36429\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__36435\,
            I => \N__36426\
        );

    \I__7445\ : Span4Mux_h
    port map (
            O => \N__36432\,
            I => \N__36423\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36429\,
            I => \pid_front.pid_preregZ0Z_12\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36426\,
            I => \pid_front.pid_preregZ0Z_12\
        );

    \I__7442\ : Odrv4
    port map (
            O => \N__36423\,
            I => \pid_front.pid_preregZ0Z_12\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36412\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36409\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36406\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__36409\,
            I => \pid_front.pid_preregZ0Z_16\
        );

    \I__7437\ : Odrv4
    port map (
            O => \N__36406\,
            I => \pid_front.pid_preregZ0Z_16\
        );

    \I__7436\ : InMux
    port map (
            O => \N__36401\,
            I => \N__36398\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36393\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36390\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36396\,
            I => \N__36387\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__36393\,
            I => \N__36383\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36390\,
            I => \N__36380\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36387\,
            I => \N__36377\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36386\,
            I => \N__36374\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__36383\,
            I => \N__36371\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__36380\,
            I => \N__36368\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__36377\,
            I => \N__36365\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36374\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__36371\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__7423\ : Odrv4
    port map (
            O => \N__36368\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__7422\ : Odrv4
    port map (
            O => \N__36365\,
            I => \pid_front.pid_preregZ0Z_2\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36356\,
            I => \N__36352\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36349\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36349\,
            I => \pid_front.pid_preregZ0Z_15\
        );

    \I__7417\ : Odrv4
    port map (
            O => \N__36346\,
            I => \pid_front.pid_preregZ0Z_15\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36341\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36338\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36330\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36327\
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__36333\,
            I => \N__36324\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__36330\,
            I => \N__36321\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36327\,
            I => \N__36318\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36315\
        );

    \I__7408\ : Span12Mux_h
    port map (
            O => \N__36321\,
            I => \N__36312\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__36318\,
            I => \N__36309\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36315\,
            I => front_order_11
        );

    \I__7405\ : Odrv12
    port map (
            O => \N__36312\,
            I => front_order_11
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__36309\,
            I => front_order_11
        );

    \I__7403\ : CascadeMux
    port map (
            O => \N__36302\,
            I => \N__36299\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36299\,
            I => \N__36296\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__7400\ : Span4Mux_v
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__36290\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36287\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__7397\ : CascadeMux
    port map (
            O => \N__36284\,
            I => \N__36281\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__36278\,
            I => \N__36274\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36271\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__36274\,
            I => \N__36268\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__36271\,
            I => \N__36265\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__36268\,
            I => front_order_12
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__36265\,
            I => front_order_12
        );

    \I__7389\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36257\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__7387\ : Span4Mux_h
    port map (
            O => \N__36254\,
            I => \N__36251\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__36251\,
            I => \N__36248\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__36248\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__7384\ : InMux
    port map (
            O => \N__36245\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36242\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__7382\ : InMux
    port map (
            O => \N__36239\,
            I => \ppm_encoder_1.un1_elevator_cry_13\
        );

    \I__7381\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36232\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36228\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36232\,
            I => \N__36225\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36222\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36219\
        );

    \I__7376\ : Span4Mux_h
    port map (
            O => \N__36225\,
            I => \N__36216\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36213\
        );

    \I__7374\ : Odrv4
    port map (
            O => \N__36219\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__36216\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__7372\ : Odrv4
    port map (
            O => \N__36213\,
            I => \pid_front.pid_preregZ0Z_0\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36203\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__36203\,
            I => \N__36200\
        );

    \I__7369\ : Odrv4
    port map (
            O => \N__36200\,
            I => \pid_front.un1_reset_i_a5_1_7\
        );

    \I__7368\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36193\
        );

    \I__7367\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36189\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36186\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36192\,
            I => \N__36183\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36180\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__36186\,
            I => \N__36177\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36183\,
            I => \N__36174\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__36180\,
            I => front_order_1
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__36177\,
            I => front_order_1
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__36174\,
            I => front_order_1
        );

    \I__7358\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36164\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__7356\ : Odrv12
    port map (
            O => \N__36161\,
            I => \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\
        );

    \I__7355\ : InMux
    port map (
            O => \N__36158\,
            I => \ppm_encoder_1.un1_elevator_cry_0\
        );

    \I__7354\ : InMux
    port map (
            O => \N__36155\,
            I => \ppm_encoder_1.un1_elevator_cry_1\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__36149\,
            I => \N__36144\
        );

    \I__7351\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36141\
        );

    \I__7350\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36138\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__36144\,
            I => \N__36135\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__36141\,
            I => \N__36132\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__36138\,
            I => front_order_3
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__36135\,
            I => front_order_3
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__36132\,
            I => front_order_3
        );

    \I__7344\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36122\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__36122\,
            I => \N__36119\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__36119\,
            I => \N__36116\
        );

    \I__7341\ : Span4Mux_v
    port map (
            O => \N__36116\,
            I => \N__36113\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__36113\,
            I => \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36110\,
            I => \ppm_encoder_1.un1_elevator_cry_2\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36107\,
            I => \ppm_encoder_1.un1_elevator_cry_3\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36104\,
            I => \ppm_encoder_1.un1_elevator_cry_4\
        );

    \I__7336\ : InMux
    port map (
            O => \N__36101\,
            I => \ppm_encoder_1.un1_elevator_cry_5\
        );

    \I__7335\ : InMux
    port map (
            O => \N__36098\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36095\,
            I => \bfn_15_19_0_\
        );

    \I__7333\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36087\
        );

    \I__7332\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36084\
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__36090\,
            I => \N__36081\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36087\,
            I => \N__36078\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36084\,
            I => \N__36075\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36072\
        );

    \I__7327\ : Span4Mux_v
    port map (
            O => \N__36078\,
            I => \N__36067\
        );

    \I__7326\ : Span4Mux_v
    port map (
            O => \N__36075\,
            I => \N__36067\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36072\,
            I => front_order_9
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__36067\,
            I => front_order_9
        );

    \I__7323\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__36056\,
            I => \N__36053\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__36053\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__7319\ : CascadeMux
    port map (
            O => \N__36050\,
            I => \N__36047\
        );

    \I__7318\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36044\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__36041\,
            I => \N__36038\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36033\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36030\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36036\,
            I => \N__36027\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__36033\,
            I => side_order_10
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__36030\,
            I => side_order_10
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__36027\,
            I => side_order_10
        );

    \I__7309\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36011\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36011\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36011\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__36011\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36008\,
            I => \N__36004\
        );

    \I__7304\ : InMux
    port map (
            O => \N__36007\,
            I => \N__36001\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__36004\,
            I => \N__35996\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35996\
        );

    \I__7301\ : Odrv12
    port map (
            O => \N__35996\,
            I => \pid_side.N_531\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__35993\,
            I => \N__35990\
        );

    \I__7299\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35987\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__35987\,
            I => \pid_side.un1_reset_i_a5_0_5\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35981\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__35981\,
            I => \pid_side.un1_reset_i_1\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35973\
        );

    \I__7294\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35970\
        );

    \I__7293\ : InMux
    port map (
            O => \N__35976\,
            I => \N__35967\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__35973\,
            I => \N__35962\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35962\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__35967\,
            I => side_order_1
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__35962\,
            I => side_order_1
        );

    \I__7288\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35953\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35956\,
            I => \N__35950\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__35953\,
            I => \N__35945\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__35950\,
            I => \N__35942\
        );

    \I__7284\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35937\
        );

    \I__7283\ : InMux
    port map (
            O => \N__35948\,
            I => \N__35937\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__35945\,
            I => \pid_side.pid_preregZ0Z_2\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__35942\,
            I => \pid_side.pid_preregZ0Z_2\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__35937\,
            I => \pid_side.pid_preregZ0Z_2\
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__35930\,
            I => \N__35925\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35922\
        );

    \I__7277\ : CascadeMux
    port map (
            O => \N__35928\,
            I => \N__35919\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35916\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35913\
        );

    \I__7274\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35910\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__35916\,
            I => \N__35907\
        );

    \I__7272\ : Span4Mux_h
    port map (
            O => \N__35913\,
            I => \N__35904\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__35910\,
            I => side_order_2
        );

    \I__7270\ : Odrv12
    port map (
            O => \N__35907\,
            I => side_order_2
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__35904\,
            I => side_order_2
        );

    \I__7268\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35882\
        );

    \I__7267\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35879\
        );

    \I__7266\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35868\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35894\,
            I => \N__35868\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35868\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35868\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35852\
        );

    \I__7261\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35852\
        );

    \I__7260\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35852\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35852\
        );

    \I__7258\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35852\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35852\
        );

    \I__7256\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35852\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__35882\,
            I => \N__35849\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__35879\,
            I => \N__35846\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35843\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__35877\,
            I => \N__35840\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__35868\,
            I => \N__35837\
        );

    \I__7250\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35834\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35831\
        );

    \I__7248\ : Span4Mux_h
    port map (
            O => \N__35849\,
            I => \N__35828\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__35846\,
            I => \N__35823\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35823\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35820\
        );

    \I__7244\ : Span4Mux_h
    port map (
            O => \N__35837\,
            I => \N__35817\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35814\
        );

    \I__7242\ : Span4Mux_v
    port map (
            O => \N__35831\,
            I => \N__35809\
        );

    \I__7241\ : Span4Mux_v
    port map (
            O => \N__35828\,
            I => \N__35809\
        );

    \I__7240\ : Span4Mux_h
    port map (
            O => \N__35823\,
            I => \N__35806\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__35820\,
            I => \N__35803\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__35817\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__7237\ : Odrv4
    port map (
            O => \N__35814\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__35809\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__35806\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__7234\ : Odrv12
    port map (
            O => \N__35803\,
            I => \pid_side.stateZ0Z_1\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__35792\,
            I => \N__35789\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35784\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35780\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__35787\,
            I => \N__35777\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__35784\,
            I => \N__35774\
        );

    \I__7228\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35771\
        );

    \I__7227\ : LocalMux
    port map (
            O => \N__35780\,
            I => \N__35768\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35765\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__35774\,
            I => \N__35758\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35758\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__35768\,
            I => \N__35758\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__35765\,
            I => \pid_side.pid_preregZ0Z_3\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__35758\,
            I => \pid_side.pid_preregZ0Z_3\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__35753\,
            I => \pid_side.N_291_cascade_\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35738\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35738\
        );

    \I__7217\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35738\
        );

    \I__7216\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35738\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__35738\,
            I => \pid_side.N_451_1\
        );

    \I__7214\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35732\,
            I => \N__35728\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__35731\,
            I => \N__35724\
        );

    \I__7211\ : Span4Mux_h
    port map (
            O => \N__35728\,
            I => \N__35721\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35727\,
            I => \N__35718\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35715\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__35721\,
            I => \N__35712\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__35718\,
            I => \N__35709\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__35715\,
            I => front_order_0
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__35712\,
            I => front_order_0
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__35709\,
            I => front_order_0
        );

    \I__7203\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35696\
        );

    \I__7202\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35696\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__35696\,
            I => \N__35692\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35689\
        );

    \I__7199\ : Span4Mux_v
    port map (
            O => \N__35692\,
            I => \N__35686\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35689\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__35686\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35678\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__35678\,
            I => \ppm_encoder_1.N_295\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__35675\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35669\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35669\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35666\,
            I => \N__35659\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35665\,
            I => \N__35659\
        );

    \I__7189\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35656\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__35659\,
            I => \N__35653\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__35656\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__7186\ : Odrv12
    port map (
            O => \N__35653\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35648\,
            I => \N__35642\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35642\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35642\,
            I => \N__35638\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35635\
        );

    \I__7181\ : Span4Mux_v
    port map (
            O => \N__35638\,
            I => \N__35632\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35635\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__35632\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35624\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__35624\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35616\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35613\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35610\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__35616\,
            I => \N__35607\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35604\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35610\,
            I => \N__35597\
        );

    \I__7170\ : Span4Mux_v
    port map (
            O => \N__35607\,
            I => \N__35597\
        );

    \I__7169\ : Span4Mux_v
    port map (
            O => \N__35604\,
            I => \N__35597\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__35597\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35588\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__35588\,
            I => \N__35584\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35581\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__35584\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__35581\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__35576\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\
        );

    \I__7160\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35567\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__35567\,
            I => \N__35564\
        );

    \I__7157\ : Odrv12
    port map (
            O => \N__35564\,
            I => \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35558\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35558\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35552\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35552\,
            I => \N__35549\
        );

    \I__7152\ : Odrv12
    port map (
            O => \N__35549\,
            I => \ppm_encoder_1.N_296\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35546\,
            I => \N__35543\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35543\,
            I => \ppm_encoder_1.N_287\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35537\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__35537\,
            I => \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35531\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__35531\,
            I => \N__35528\
        );

    \I__7145\ : Span4Mux_h
    port map (
            O => \N__35528\,
            I => \N__35525\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35525\,
            I => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35518\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35514\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35518\,
            I => \N__35511\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35508\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35514\,
            I => \N__35503\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__35511\,
            I => \N__35503\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__35508\,
            I => \N__35500\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__35503\,
            I => throttle_order_1
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__35500\,
            I => throttle_order_1
        );

    \I__7134\ : InMux
    port map (
            O => \N__35495\,
            I => \N__35492\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__35492\,
            I => \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__35489\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35480\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__35477\,
            I => \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35474\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35468\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__35465\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35462\,
            I => \bfn_15_13_0_\
        );

    \I__7122\ : CascadeMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35453\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__35450\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35444\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35444\,
            I => \N__35441\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__35441\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35438\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35435\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__7113\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__35426\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__7110\ : CascadeMux
    port map (
            O => \N__35423\,
            I => \N__35419\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35416\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35413\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__35416\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35413\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35408\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35402\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35399\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__35396\,
            I => \N__35393\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35390\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__35387\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35384\,
            I => \bfn_15_12_0_\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35381\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35378\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35372\,
            I => \N__35368\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35365\
        );

    \I__7091\ : Sp12to4
    port map (
            O => \N__35368\,
            I => \N__35360\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__35365\,
            I => \N__35360\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__35360\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35351\,
            I => \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\
        );

    \I__7085\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__7083\ : Odrv4
    port map (
            O => \N__35342\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35339\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35333\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35333\,
            I => \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35327\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35327\,
            I => \N__35324\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__35324\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35321\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35318\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35315\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35312\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35306\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__7070\ : InMux
    port map (
            O => \N__35303\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35300\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__7068\ : InMux
    port map (
            O => \N__35297\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__7067\ : InMux
    port map (
            O => \N__35294\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__7066\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35288\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35288\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__7064\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35276\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35276\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35276\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__35276\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35265\
        );

    \I__7058\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35262\
        );

    \I__7057\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35259\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__35265\,
            I => \N__35254\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__35262\,
            I => \N__35254\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__35259\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__35254\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__35249\,
            I => \ppm_encoder_1.N_313_cascade_\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35243\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__35243\,
            I => \reset_module_System.count_1_2\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35236\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35233\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__35236\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__35233\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7045\ : CascadeMux
    port map (
            O => \N__35228\,
            I => \N__35225\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35216\
        );

    \I__7043\ : InMux
    port map (
            O => \N__35224\,
            I => \N__35216\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35223\,
            I => \N__35216\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35216\,
            I => \reset_module_System.reset6_15\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__35213\,
            I => \N__35208\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35204\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35201\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35196\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35196\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35204\,
            I => \reset_module_System.reset6_14\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__35201\,
            I => \reset_module_System.reset6_14\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35196\,
            I => \reset_module_System.reset6_14\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35185\
        );

    \I__7031\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35182\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35185\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35182\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__7028\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35173\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35170\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__35173\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__35170\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__35165\,
            I => \N__35161\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35158\
        );

    \I__7022\ : InMux
    port map (
            O => \N__35161\,
            I => \N__35155\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35158\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__35155\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35146\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35143\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35146\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__35143\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__7015\ : InMux
    port map (
            O => \N__35138\,
            I => \N__35134\
        );

    \I__7014\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35131\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35134\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__35131\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__7011\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35121\
        );

    \I__7010\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35118\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35115\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__35121\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__35118\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__35115\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__7005\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35105\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35105\,
            I => \N__35101\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35098\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__35101\,
            I => \N__35095\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__35098\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__35095\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35086\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35083\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__35086\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__35083\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__6995\ : CascadeMux
    port map (
            O => \N__35078\,
            I => \reset_module_System.reset6_3_cascade_\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35072\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__35072\,
            I => \reset_module_System.reset6_13\
        );

    \I__6992\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35065\
        );

    \I__6991\ : InMux
    port map (
            O => \N__35068\,
            I => \N__35062\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35065\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__35062\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__35051\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35056\,
            I => \N__35048\
        );

    \I__6986\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35045\
        );

    \I__6985\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35042\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35039\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__35048\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35045\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35042\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__35039\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__35030\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__6978\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__35024\,
            I => \N__35021\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__35021\,
            I => \reset_module_System.reset6_11\
        );

    \I__6975\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35012\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35017\,
            I => \N__35005\
        );

    \I__6973\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35005\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35005\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35012\,
            I => \reset_module_System.reset6_19\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35005\,
            I => \reset_module_System.reset6_19\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34997\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__34997\,
            I => \N__34994\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__34994\,
            I => \N__34991\
        );

    \I__6966\ : Span4Mux_h
    port map (
            O => \N__34991\,
            I => \N__34988\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__34988\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__6964\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34982\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__34979\,
            I => \N__34975\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34978\,
            I => \N__34972\
        );

    \I__6960\ : Span4Mux_h
    port map (
            O => \N__34975\,
            I => \N__34969\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34966\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__34969\,
            I => scaler_4_data_9
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__34966\,
            I => scaler_4_data_9
        );

    \I__6956\ : CascadeMux
    port map (
            O => \N__34961\,
            I => \N__34958\
        );

    \I__6955\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34955\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__34955\,
            I => \pid_front.m7_e_4\
        );

    \I__6953\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34948\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34951\,
            I => \N__34945\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34948\,
            I => \pid_front.pid_preregZ0Z_18\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34945\,
            I => \pid_front.pid_preregZ0Z_18\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__34940\,
            I => \N__34936\
        );

    \I__6948\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34933\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34930\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__34933\,
            I => \pid_front.pid_preregZ0Z_19\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__34930\,
            I => \pid_front.pid_preregZ0Z_19\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34918\
        );

    \I__6943\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34918\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__34923\,
            I => \N__34914\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34911\
        );

    \I__6940\ : CascadeMux
    port map (
            O => \N__34917\,
            I => \N__34908\
        );

    \I__6939\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34905\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__34911\,
            I => \N__34902\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34899\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34905\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__34902\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__34899\,
            I => \pid_front.pid_preregZ0Z_9\
        );

    \I__6933\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34888\
        );

    \I__6932\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34885\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34888\,
            I => \N__34881\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34878\
        );

    \I__6929\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34874\
        );

    \I__6928\ : Span4Mux_v
    port map (
            O => \N__34881\,
            I => \N__34871\
        );

    \I__6927\ : Span12Mux_v
    port map (
            O => \N__34878\,
            I => \N__34868\
        );

    \I__6926\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34865\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__34874\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6924\ : Odrv4
    port map (
            O => \N__34871\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6923\ : Odrv12
    port map (
            O => \N__34868\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34865\,
            I => \pid_front.pid_preregZ0Z_11\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34848\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34848\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34842\
        );

    \I__6918\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34842\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34838\
        );

    \I__6916\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34835\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__34842\,
            I => \N__34832\
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__34841\,
            I => \N__34829\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__34838\,
            I => \N__34822\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34835\,
            I => \N__34822\
        );

    \I__6911\ : Span4Mux_h
    port map (
            O => \N__34832\,
            I => \N__34822\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34818\
        );

    \I__6909\ : Span4Mux_v
    port map (
            O => \N__34822\,
            I => \N__34815\
        );

    \I__6908\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34812\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__34818\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__34815\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__34812\,
            I => \pid_front.pid_preregZ0Z_13\
        );

    \I__6904\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34801\
        );

    \I__6903\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34798\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34801\,
            I => \N__34795\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34798\,
            I => \pid_side.pid_preregZ0Z_15\
        );

    \I__6900\ : Odrv12
    port map (
            O => \N__34795\,
            I => \pid_side.pid_preregZ0Z_15\
        );

    \I__6899\ : CascadeMux
    port map (
            O => \N__34790\,
            I => \N__34786\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34783\
        );

    \I__6897\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34780\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34783\,
            I => \N__34777\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34780\,
            I => \pid_side.pid_preregZ0Z_14\
        );

    \I__6894\ : Odrv12
    port map (
            O => \N__34777\,
            I => \pid_side.pid_preregZ0Z_14\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__34772\,
            I => \N__34769\
        );

    \I__6892\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34763\
        );

    \I__6890\ : Span4Mux_h
    port map (
            O => \N__34763\,
            I => \N__34760\
        );

    \I__6889\ : Odrv4
    port map (
            O => \N__34760\,
            I => \pid_side.m7_e_4\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34754\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34750\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34747\
        );

    \I__6885\ : Span4Mux_v
    port map (
            O => \N__34750\,
            I => \N__34744\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__34747\,
            I => \pid_side.pid_preregZ0Z_16\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__34744\,
            I => \pid_side.pid_preregZ0Z_16\
        );

    \I__6882\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__34736\,
            I => \pid_side.un1_reset_i_a5_1_7\
        );

    \I__6880\ : CascadeMux
    port map (
            O => \N__34733\,
            I => \pid_side.N_563_cascade_\
        );

    \I__6879\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__34727\,
            I => \pid_side.un1_reset_i_a5_1_8\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__34724\,
            I => \pid_side.N_311_cascade_\
        );

    \I__6876\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34718\,
            I => \pid_side.un1_reset_i_a5_1_6\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__6872\ : Span4Mux_v
    port map (
            O => \N__34709\,
            I => \N__34705\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34702\
        );

    \I__6870\ : Span4Mux_h
    port map (
            O => \N__34705\,
            I => \N__34698\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34695\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34692\
        );

    \I__6867\ : Sp12to4
    port map (
            O => \N__34698\,
            I => \N__34687\
        );

    \I__6866\ : Span12Mux_v
    port map (
            O => \N__34695\,
            I => \N__34687\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__34692\,
            I => \pid_side.error_p_regZ0Z_2\
        );

    \I__6864\ : Odrv12
    port map (
            O => \N__34687\,
            I => \pid_side.error_p_regZ0Z_2\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__34682\,
            I => \N__34679\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34676\,
            I => \N__34673\
        );

    \I__6860\ : Span4Mux_h
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__34670\,
            I => \N__34667\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__34667\,
            I => \pid_side.un1_pid_prereg_cry_1_THRU_CO\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34661\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__6855\ : Odrv12
    port map (
            O => \N__34658\,
            I => \pid_side.un1_reset_i_a5_0_2\
        );

    \I__6854\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__34646\,
            I => \pid_side.un1_reset_i_a5_0_3\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34637\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34634\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34628\
        );

    \I__6847\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34628\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34625\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__34634\,
            I => \N__34622\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34619\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34628\,
            I => \pid_front.N_569\
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__34625\,
            I => \pid_front.N_569\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__34622\,
            I => \pid_front.N_569\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34619\,
            I => \pid_front.N_569\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34604\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34609\,
            I => \N__34604\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34604\,
            I => \pid_front.pid_preregZ0Z_14\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34598\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34598\,
            I => \N__34595\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__34595\,
            I => \N__34590\
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__34594\,
            I => \N__34587\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34583\
        );

    \I__6831\ : Span4Mux_h
    port map (
            O => \N__34590\,
            I => \N__34580\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34587\,
            I => \N__34575\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34586\,
            I => \N__34575\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34583\,
            I => \pid_side.pid_preregZ0Z_8\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__34580\,
            I => \pid_side.pid_preregZ0Z_8\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34575\,
            I => \pid_side.pid_preregZ0Z_8\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34562\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__34562\,
            I => \N__34556\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34551\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34551\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34548\
        );

    \I__6819\ : Span4Mux_h
    port map (
            O => \N__34556\,
            I => \N__34543\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34543\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34548\,
            I => \pid_side.pid_preregZ0Z_9\
        );

    \I__6816\ : Odrv4
    port map (
            O => \N__34543\,
            I => \pid_side.pid_preregZ0Z_9\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34526\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34526\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34526\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34526\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__34526\,
            I => \N__34521\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34525\,
            I => \N__34518\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34524\,
            I => \N__34511\
        );

    \I__6808\ : Span4Mux_h
    port map (
            O => \N__34521\,
            I => \N__34506\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34506\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34503\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34497\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34497\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34494\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__34511\,
            I => \N__34489\
        );

    \I__6801\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34489\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__34503\,
            I => \N__34486\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34483\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34497\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34494\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__34489\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__34486\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34483\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34469\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__34469\,
            I => \N__34463\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34456\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34456\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34456\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__34463\,
            I => \N__34453\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34456\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__34453\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6783\ : Odrv4
    port map (
            O => \N__34442\,
            I => \uart_drone.CO0\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34436\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__34433\,
            I => \N__34427\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34424\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34421\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34418\
        );

    \I__6776\ : Sp12to4
    port map (
            O => \N__34427\,
            I => \N__34413\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34424\,
            I => \N__34413\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__34421\,
            I => \pid_side.pid_preregZ0Z_11\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34418\,
            I => \pid_side.pid_preregZ0Z_11\
        );

    \I__6772\ : Odrv12
    port map (
            O => \N__34413\,
            I => \pid_side.pid_preregZ0Z_11\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34403\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34397\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34394\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34391\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34400\,
            I => \N__34388\
        );

    \I__6766\ : Span4Mux_v
    port map (
            O => \N__34397\,
            I => \N__34383\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34394\,
            I => \N__34383\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34391\,
            I => \pid_side.pid_preregZ0Z_7\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34388\,
            I => \pid_side.pid_preregZ0Z_7\
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__34383\,
            I => \pid_side.pid_preregZ0Z_7\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__34370\,
            I => \N__34367\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__34367\,
            I => \pid_side.un1_reset_i_a5_1_5\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34361\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34361\,
            I => \N__34358\
        );

    \I__6755\ : Odrv12
    port map (
            O => \N__34358\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34355\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34346\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__34346\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34343\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34340\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34337\,
            I => \ppm_encoder_1.un1_aileron_cry_13\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34331\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__34331\,
            I => \N__34328\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__34328\,
            I => \N__34323\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34320\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34317\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__34323\,
            I => \N__34314\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34320\,
            I => \N__34311\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34308\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__34314\,
            I => \N__34303\
        );

    \I__6738\ : Span4Mux_v
    port map (
            O => \N__34311\,
            I => \N__34303\
        );

    \I__6737\ : Span12Mux_s1_h
    port map (
            O => \N__34308\,
            I => \N__34300\
        );

    \I__6736\ : Sp12to4
    port map (
            O => \N__34303\,
            I => \N__34297\
        );

    \I__6735\ : Span12Mux_h
    port map (
            O => \N__34300\,
            I => \N__34293\
        );

    \I__6734\ : Span12Mux_h
    port map (
            O => \N__34297\,
            I => \N__34290\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34287\
        );

    \I__6732\ : Odrv12
    port map (
            O => \N__34293\,
            I => drone_altitude_0
        );

    \I__6731\ : Odrv12
    port map (
            O => \N__34290\,
            I => drone_altitude_0
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__34287\,
            I => drone_altitude_0
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__34280\,
            I => \N__34277\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34270\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34267\
        );

    \I__6725\ : Span12Mux_v
    port map (
            O => \N__34270\,
            I => \N__34264\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__34267\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__6723\ : Odrv12
    port map (
            O => \N__34264\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34256\,
            I => \N__34253\
        );

    \I__6720\ : Span4Mux_v
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__34250\,
            I => \N__34244\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34237\
        );

    \I__6717\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34237\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34237\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__34244\,
            I => \pid_side.pid_preregZ0Z_10\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__34237\,
            I => \pid_side.pid_preregZ0Z_10\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__34232\,
            I => \N__34228\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34225\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34228\,
            I => \N__34221\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__34225\,
            I => \N__34218\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34215\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34221\,
            I => side_order_11
        );

    \I__6707\ : Odrv12
    port map (
            O => \N__34218\,
            I => side_order_11
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__34215\,
            I => side_order_11
        );

    \I__6705\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34205\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34201\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__34204\,
            I => \N__34197\
        );

    \I__6702\ : Span4Mux_h
    port map (
            O => \N__34201\,
            I => \N__34194\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__34200\,
            I => \N__34190\
        );

    \I__6700\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34187\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__34194\,
            I => \N__34184\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34181\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34178\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__34187\,
            I => \pid_side.pid_preregZ0Z_6\
        );

    \I__6695\ : Odrv4
    port map (
            O => \N__34184\,
            I => \pid_side.pid_preregZ0Z_6\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34181\,
            I => \pid_side.pid_preregZ0Z_6\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__34178\,
            I => \pid_side.pid_preregZ0Z_6\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34169\,
            I => \ppm_encoder_1.un1_aileron_cry_1\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34166\,
            I => \ppm_encoder_1.un1_aileron_cry_2\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34163\,
            I => \ppm_encoder_1.un1_aileron_cry_3\
        );

    \I__6689\ : InMux
    port map (
            O => \N__34160\,
            I => \ppm_encoder_1.un1_aileron_cry_4\
        );

    \I__6688\ : InMux
    port map (
            O => \N__34157\,
            I => \ppm_encoder_1.un1_aileron_cry_5\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34154\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34151\,
            I => \bfn_14_15_0_\
        );

    \I__6685\ : InMux
    port map (
            O => \N__34148\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34145\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__6683\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34137\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34134\
        );

    \I__6681\ : InMux
    port map (
            O => \N__34140\,
            I => \N__34131\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34128\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34134\,
            I => \N__34125\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__34131\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__6677\ : Odrv12
    port map (
            O => \N__34128\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__6676\ : Odrv4
    port map (
            O => \N__34125\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__34118\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34112\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34112\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__34109\,
            I => \N__34104\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34099\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34099\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34096\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34093\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__34096\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__34093\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__34088\,
            I => \ppm_encoder_1.N_298_cascade_\
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \N__34080\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34084\,
            I => \N__34075\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34075\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34080\,
            I => \N__34072\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__34075\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__34072\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34062\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34057\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34057\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34062\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__34057\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__6653\ : InMux
    port map (
            O => \N__34052\,
            I => \ppm_encoder_1.un1_aileron_cry_0\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34046\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34042\
        );

    \I__6650\ : CascadeMux
    port map (
            O => \N__34045\,
            I => \N__34039\
        );

    \I__6649\ : Span4Mux_v
    port map (
            O => \N__34042\,
            I => \N__34036\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34033\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__34036\,
            I => \N__34030\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__34033\,
            I => \N__34027\
        );

    \I__6645\ : Odrv4
    port map (
            O => \N__34030\,
            I => scaler_4_data_10
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__34027\,
            I => scaler_4_data_10
        );

    \I__6643\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34019\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__34019\,
            I => \N__34016\
        );

    \I__6641\ : Span4Mux_v
    port map (
            O => \N__34016\,
            I => \N__34013\
        );

    \I__6640\ : Odrv4
    port map (
            O => \N__34013\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__6639\ : CascadeMux
    port map (
            O => \N__34010\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34004\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__34004\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33996\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33991\
        );

    \I__6634\ : InMux
    port map (
            O => \N__33999\,
            I => \N__33991\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__33996\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33991\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__33986\,
            I => \ppm_encoder_1.N_297_cascade_\
        );

    \I__6630\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33974\
        );

    \I__6629\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33974\
        );

    \I__6628\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33974\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__33974\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__6626\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33962\
        );

    \I__6625\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33962\
        );

    \I__6624\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33962\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__33962\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__6621\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33952\
        );

    \I__6620\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33949\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33952\,
            I => \N__33946\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33949\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__33946\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33941\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__6615\ : InMux
    port map (
            O => \N__33938\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__33935\,
            I => \N__33932\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33926\
        );

    \I__6612\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33926\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__33926\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__6610\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33919\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33916\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__33919\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__33916\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__6606\ : CascadeMux
    port map (
            O => \N__33911\,
            I => \N__33907\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33902\
        );

    \I__6604\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33902\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__33902\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33895\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33892\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33895\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__33892\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33884\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33880\
        );

    \I__6596\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__6595\ : Odrv4
    port map (
            O => \N__33880\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__33877\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__6593\ : InMux
    port map (
            O => \N__33872\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33869\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33866\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__6590\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33860\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__33860\,
            I => \N__33856\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33853\
        );

    \I__6587\ : Odrv4
    port map (
            O => \N__33856\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__33853\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33848\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33845\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33842\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__33839\,
            I => \N__33836\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33836\,
            I => \N__33833\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33833\,
            I => \N__33829\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33826\
        );

    \I__6578\ : Odrv12
    port map (
            O => \N__33829\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33826\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__6576\ : InMux
    port map (
            O => \N__33821\,
            I => \bfn_14_9_0_\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33818\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33815\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33812\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33805\
        );

    \I__6571\ : InMux
    port map (
            O => \N__33808\,
            I => \N__33802\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__33805\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__33802\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33797\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33794\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33791\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33784\
        );

    \I__6564\ : InMux
    port map (
            O => \N__33787\,
            I => \N__33781\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33784\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33781\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__6561\ : InMux
    port map (
            O => \N__33776\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__6560\ : InMux
    port map (
            O => \N__33773\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33770\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33767\,
            I => \bfn_14_8_0_\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33761\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__33761\,
            I => \N__33757\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33754\
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__33757\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__33754\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33749\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__33746\,
            I => \pid_front.un1_reset_i_a5_1_5_cascade_\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__33743\,
            I => \N__33740\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33737\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__33737\,
            I => \N__33734\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__33734\,
            I => \pid_front.un1_reset_i_a5_1_8\
        );

    \I__6546\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33727\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33724\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__33727\,
            I => \N__33718\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33724\,
            I => \N__33718\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33714\
        );

    \I__6541\ : Span4Mux_v
    port map (
            O => \N__33718\,
            I => \N__33711\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33708\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33714\,
            I => \pid_front.pid_preregZ0Z_10\
        );

    \I__6538\ : Odrv4
    port map (
            O => \N__33711\,
            I => \pid_front.pid_preregZ0Z_10\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__33708\,
            I => \pid_front.pid_preregZ0Z_10\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33701\,
            I => \N__33698\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__33698\,
            I => \dron_frame_decoder_1.drone_H_disp_front_8\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__33695\,
            I => \reset_module_System.reset6_15_cascade_\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33689\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33689\,
            I => \reset_module_System.count_1_1\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__33686\,
            I => \N__33682\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__33685\,
            I => \N__33675\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33666\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33666\
        );

    \I__6527\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33666\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33666\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33653\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33650\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33647\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33665\,
            I => \N__33642\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33642\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33639\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33628\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33628\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33628\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33628\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33628\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33625\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33622\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33617\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33617\
        );

    \I__6510\ : Sp12to4
    port map (
            O => \N__33647\,
            I => \N__33602\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__33642\,
            I => \N__33602\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33602\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33602\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__33625\,
            I => \N__33602\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__33622\,
            I => \N__33602\
        );

    \I__6504\ : Sp12to4
    port map (
            O => \N__33617\,
            I => \N__33602\
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__33602\,
            I => \pid_front.stateZ0Z_1\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__33599\,
            I => \N__33594\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__33598\,
            I => \N__33590\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33575\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33575\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33575\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33575\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33575\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33575\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33569\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33564\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33564\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33561\
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__33569\,
            I => \pid_front.N_287\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33564\,
            I => \pid_front.N_287\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33561\,
            I => \pid_front.N_287\
        );

    \I__6487\ : CascadeMux
    port map (
            O => \N__33554\,
            I => \N__33550\
        );

    \I__6486\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33545\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33545\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__33545\,
            I => \pid_front.N_533\
        );

    \I__6483\ : CEMux
    port map (
            O => \N__33542\,
            I => \N__33539\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__33536\,
            I => \pid_front.state_0_1\
        );

    \I__6480\ : SRMux
    port map (
            O => \N__33533\,
            I => \N__33530\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__33527\,
            I => \N__33523\
        );

    \I__6477\ : SRMux
    port map (
            O => \N__33526\,
            I => \N__33520\
        );

    \I__6476\ : Span4Mux_h
    port map (
            O => \N__33523\,
            I => \N__33514\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__33520\,
            I => \N__33514\
        );

    \I__6474\ : SRMux
    port map (
            O => \N__33519\,
            I => \N__33511\
        );

    \I__6473\ : Span4Mux_v
    port map (
            O => \N__33514\,
            I => \N__33507\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33511\,
            I => \N__33504\
        );

    \I__6471\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33501\
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__33507\,
            I => \pid_front.pid_prereg_RNI2A6A6Z0Z_2\
        );

    \I__6469\ : Odrv12
    port map (
            O => \N__33504\,
            I => \pid_front.pid_prereg_RNI2A6A6Z0Z_2\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33501\,
            I => \pid_front.pid_prereg_RNI2A6A6Z0Z_2\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__33491\,
            I => \pid_front.un1_reset_i_a5_1_6\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33482\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__33482\,
            I => \pid_front.N_315\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33476\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__33476\,
            I => \drone_H_disp_front_1\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__33473\,
            I => \pid_side.state_ns_0_cascade_\
        );

    \I__6459\ : CEMux
    port map (
            O => \N__33470\,
            I => \N__33466\
        );

    \I__6458\ : CEMux
    port map (
            O => \N__33469\,
            I => \N__33463\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33459\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33456\
        );

    \I__6455\ : CEMux
    port map (
            O => \N__33462\,
            I => \N__33453\
        );

    \I__6454\ : Span4Mux_h
    port map (
            O => \N__33459\,
            I => \N__33450\
        );

    \I__6453\ : Span4Mux_v
    port map (
            O => \N__33456\,
            I => \N__33447\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33444\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__33450\,
            I => \N__33439\
        );

    \I__6450\ : Span4Mux_h
    port map (
            O => \N__33447\,
            I => \N__33439\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__33444\,
            I => \N__33436\
        );

    \I__6448\ : Span4Mux_h
    port map (
            O => \N__33439\,
            I => \N__33433\
        );

    \I__6447\ : Span4Mux_v
    port map (
            O => \N__33436\,
            I => \N__33430\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__33433\,
            I => \dron_frame_decoder_1.N_763_0\
        );

    \I__6445\ : Odrv4
    port map (
            O => \N__33430\,
            I => \dron_frame_decoder_1.N_763_0\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33425\,
            I => \N__33422\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33422\,
            I => \N__33419\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__33419\,
            I => \pid_front.un1_reset_i_a5_0_5\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__33416\,
            I => \pid_front.un1_reset_i_1_cascade_\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33409\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33406\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33409\,
            I => \pid_front.N_532\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33406\,
            I => \pid_front.N_532\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33398\,
            I => \pid_front.un1_reset_i_a2_3\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33390\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33394\,
            I => \N__33387\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__33393\,
            I => \N__33383\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33390\,
            I => \N__33378\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33387\,
            I => \N__33378\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33374\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33371\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__33378\,
            I => \N__33368\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__33377\,
            I => \N__33365\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33374\,
            I => \N__33360\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33371\,
            I => \N__33360\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__33368\,
            I => \N__33357\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33354\
        );

    \I__6421\ : Odrv12
    port map (
            O => \N__33360\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__33357\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__33354\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33343\
        );

    \I__6417\ : CascadeMux
    port map (
            O => \N__33346\,
            I => \N__33340\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33337\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33333\
        );

    \I__6414\ : Span12Mux_h
    port map (
            O => \N__33337\,
            I => \N__33330\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33327\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33333\,
            I => \pid_alt.N_557\
        );

    \I__6411\ : Odrv12
    port map (
            O => \N__33330\,
            I => \pid_alt.N_557\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__33327\,
            I => \pid_alt.N_557\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33315\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33308\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33308\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33315\,
            I => \N__33305\
        );

    \I__6405\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33302\
        );

    \I__6404\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33299\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__33308\,
            I => \N__33296\
        );

    \I__6402\ : Span12Mux_h
    port map (
            O => \N__33305\,
            I => \N__33293\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33286\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__33299\,
            I => \N__33286\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__33296\,
            I => \N__33286\
        );

    \I__6398\ : Odrv12
    port map (
            O => \N__33293\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__33286\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33275\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__6392\ : Span4Mux_h
    port map (
            O => \N__33269\,
            I => \N__33266\
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__33266\,
            I => \pid_alt.error_i_acummZ0Z_13\
        );

    \I__6390\ : CEMux
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33260\,
            I => \N__33257\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__33257\,
            I => \N__33252\
        );

    \I__6387\ : CEMux
    port map (
            O => \N__33256\,
            I => \N__33249\
        );

    \I__6386\ : CEMux
    port map (
            O => \N__33255\,
            I => \N__33246\
        );

    \I__6385\ : Span4Mux_h
    port map (
            O => \N__33252\,
            I => \N__33241\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__33249\,
            I => \N__33241\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33238\
        );

    \I__6382\ : Span4Mux_h
    port map (
            O => \N__33241\,
            I => \N__33235\
        );

    \I__6381\ : Span4Mux_v
    port map (
            O => \N__33238\,
            I => \N__33232\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33235\,
            I => \pid_alt.N_72_i_0\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__33232\,
            I => \pid_alt.N_72_i_0\
        );

    \I__6378\ : SRMux
    port map (
            O => \N__33227\,
            I => \N__33222\
        );

    \I__6377\ : SRMux
    port map (
            O => \N__33226\,
            I => \N__33219\
        );

    \I__6376\ : SRMux
    port map (
            O => \N__33225\,
            I => \N__33216\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33222\,
            I => \N__33213\
        );

    \I__6374\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33210\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33216\,
            I => \N__33207\
        );

    \I__6372\ : Span4Mux_h
    port map (
            O => \N__33213\,
            I => \N__33204\
        );

    \I__6371\ : Span4Mux_h
    port map (
            O => \N__33210\,
            I => \N__33201\
        );

    \I__6370\ : Span4Mux_v
    port map (
            O => \N__33207\,
            I => \N__33198\
        );

    \I__6369\ : Span4Mux_v
    port map (
            O => \N__33204\,
            I => \N__33191\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__33201\,
            I => \N__33191\
        );

    \I__6367\ : Span4Mux_s3_h
    port map (
            O => \N__33198\,
            I => \N__33188\
        );

    \I__6366\ : SRMux
    port map (
            O => \N__33197\,
            I => \N__33185\
        );

    \I__6365\ : SRMux
    port map (
            O => \N__33196\,
            I => \N__33182\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__33191\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__33188\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__33185\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__33182\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\
        );

    \I__6360\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33168\
        );

    \I__6359\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33165\
        );

    \I__6358\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33162\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__33168\,
            I => \N__33159\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33154\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33150\
        );

    \I__6354\ : Span4Mux_v
    port map (
            O => \N__33159\,
            I => \N__33147\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33144\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33157\,
            I => \N__33141\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__33154\,
            I => \N__33138\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33135\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__33150\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6348\ : Odrv4
    port map (
            O => \N__33147\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__33144\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__33141\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__33138\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__33135\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__6343\ : SRMux
    port map (
            O => \N__33122\,
            I => \N__33119\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__33119\,
            I => \N__33116\
        );

    \I__6341\ : Span4Mux_v
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__33113\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33107\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33107\,
            I => \ppm_encoder_1.N_291\
        );

    \I__6337\ : InMux
    port map (
            O => \N__33104\,
            I => \N__33101\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__33101\,
            I => \N__33097\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33092\
        );

    \I__6334\ : Span4Mux_h
    port map (
            O => \N__33097\,
            I => \N__33088\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33085\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33082\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33092\,
            I => \N__33078\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__33091\,
            I => \N__33072\
        );

    \I__6329\ : Sp12to4
    port map (
            O => \N__33088\,
            I => \N__33065\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__33085\,
            I => \N__33065\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33065\
        );

    \I__6326\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33062\
        );

    \I__6325\ : Span4Mux_h
    port map (
            O => \N__33078\,
            I => \N__33059\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33054\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33054\
        );

    \I__6322\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33049\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33072\,
            I => \N__33049\
        );

    \I__6320\ : Span12Mux_v
    port map (
            O => \N__33065\,
            I => \N__33046\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__33062\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__33059\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__33054\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__33049\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__6315\ : Odrv12
    port map (
            O => \N__33046\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__33035\,
            I => \N__33032\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33029\,
            I => \N__33024\
        );

    \I__6311\ : InMux
    port map (
            O => \N__33028\,
            I => \N__33019\
        );

    \I__6310\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33016\
        );

    \I__6309\ : Span4Mux_h
    port map (
            O => \N__33024\,
            I => \N__33013\
        );

    \I__6308\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33010\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33007\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__32999\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33016\,
            I => \N__32999\
        );

    \I__6304\ : Span4Mux_v
    port map (
            O => \N__33013\,
            I => \N__32996\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__33010\,
            I => \N__32991\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__33007\,
            I => \N__32991\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32988\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32983\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32983\
        );

    \I__6298\ : Span12Mux_v
    port map (
            O => \N__32999\,
            I => \N__32980\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__32996\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__32991\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__32988\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__32983\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__6293\ : Odrv12
    port map (
            O => \N__32980\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__6292\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32962\
        );

    \I__6291\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32962\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32959\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32955\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32952\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32949\
        );

    \I__6286\ : Span12Mux_h
    port map (
            O => \N__32955\,
            I => \N__32946\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__32952\,
            I => \N__32943\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__32949\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6283\ : Odrv12
    port map (
            O => \N__32946\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6282\ : Odrv12
    port map (
            O => \N__32943\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__6281\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32933\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__32933\,
            I => \N__32929\
        );

    \I__6279\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32926\
        );

    \I__6278\ : Span12Mux_s11_v
    port map (
            O => \N__32929\,
            I => \N__32923\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__32926\,
            I => \N__32920\
        );

    \I__6276\ : Odrv12
    port map (
            O => \N__32923\,
            I => \uart_drone.N_144_1\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__32920\,
            I => \uart_drone.N_144_1\
        );

    \I__6274\ : CascadeMux
    port map (
            O => \N__32915\,
            I => \uart_drone.N_145_cascade_\
        );

    \I__6273\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32904\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32899\
        );

    \I__6270\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32899\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__32904\,
            I => \N__32891\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32899\,
            I => \N__32888\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32883\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32883\
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__32896\,
            I => \N__32880\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32877\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32874\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__32891\,
            I => \N__32871\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__32888\,
            I => \N__32868\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32865\
        );

    \I__6259\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32862\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__32877\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__32874\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__32871\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__32868\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6254\ : Odrv4
    port map (
            O => \N__32865\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__32862\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__6252\ : IoInMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__32846\,
            I => \N__32843\
        );

    \I__6250\ : Span4Mux_s0_v
    port map (
            O => \N__32843\,
            I => \N__32838\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32835\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32828\
        );

    \I__6247\ : Span4Mux_v
    port map (
            O => \N__32838\,
            I => \N__32823\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32823\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32820\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32815\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32815\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32812\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32809\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__32823\,
            I => \N__32806\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32803\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32799\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__32812\,
            I => \N__32796\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__32809\,
            I => \N__32793\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__32806\,
            I => \N__32790\
        );

    \I__6234\ : Span4Mux_v
    port map (
            O => \N__32803\,
            I => \N__32787\
        );

    \I__6233\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32784\
        );

    \I__6232\ : Span4Mux_h
    port map (
            O => \N__32799\,
            I => \N__32781\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__32796\,
            I => \N__32776\
        );

    \I__6230\ : Span4Mux_v
    port map (
            O => \N__32793\,
            I => \N__32776\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__32790\,
            I => \debug_CH1_0A_c\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__32787\,
            I => \debug_CH1_0A_c\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__32784\,
            I => \debug_CH1_0A_c\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__32781\,
            I => \debug_CH1_0A_c\
        );

    \I__6225\ : Odrv4
    port map (
            O => \N__32776\,
            I => \debug_CH1_0A_c\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32762\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__32762\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__6222\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__32756\,
            I => \N__32753\
        );

    \I__6220\ : Span4Mux_h
    port map (
            O => \N__32753\,
            I => \N__32749\
        );

    \I__6219\ : InMux
    port map (
            O => \N__32752\,
            I => \N__32746\
        );

    \I__6218\ : Odrv4
    port map (
            O => \N__32749\,
            I => throttle_order_12
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32746\,
            I => throttle_order_12
        );

    \I__6216\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32738\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32738\,
            I => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__32735\,
            I => \N__32730\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32727\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32724\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32721\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__32727\,
            I => \N__32718\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__32724\,
            I => \N__32715\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32721\,
            I => throttle_order_3
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__32718\,
            I => throttle_order_3
        );

    \I__6206\ : Odrv4
    port map (
            O => \N__32715\,
            I => throttle_order_3
        );

    \I__6205\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32705\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32705\,
            I => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32698\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__32701\,
            I => \N__32695\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32692\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32689\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__32692\,
            I => \N__32686\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32683\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__32686\,
            I => throttle_order_5
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__32683\,
            I => throttle_order_5
        );

    \I__6195\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32675\,
            I => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__32672\,
            I => \N__32667\
        );

    \I__6192\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32664\
        );

    \I__6191\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32661\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32658\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32664\,
            I => \N__32653\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32653\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32648\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__32653\,
            I => \N__32648\
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__32648\,
            I => throttle_order_6
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__32645\,
            I => \ppm_encoder_1.N_314_cascade_\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__32642\,
            I => \ppm_encoder_1.N_288_cascade_\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32635\
        );

    \I__6181\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32632\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32627\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32627\
        );

    \I__6178\ : Odrv12
    port map (
            O => \N__32627\,
            I => scaler_4_data_11
        );

    \I__6177\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32621\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__32621\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__32618\,
            I => \N__32613\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32610\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32607\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32604\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32601\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__32607\,
            I => \N__32598\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__32604\,
            I => throttle_order_11
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__32601\,
            I => throttle_order_11
        );

    \I__6167\ : Odrv4
    port map (
            O => \N__32598\,
            I => throttle_order_11
        );

    \I__6166\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__32588\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32581\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32578\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32581\,
            I => \N__32575\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32578\,
            I => \N__32572\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__32575\,
            I => \N__32569\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__32572\,
            I => \N__32566\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__32569\,
            I => scaler_4_data_13
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__32566\,
            I => scaler_4_data_13
        );

    \I__6156\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32558\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32555\
        );

    \I__6154\ : Odrv4
    port map (
            O => \N__32555\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32549\,
            I => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__32546\,
            I => \N__32541\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32538\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32544\,
            I => \N__32535\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32532\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__32538\,
            I => \N__32529\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32535\,
            I => \N__32526\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32532\,
            I => throttle_order_2
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__32529\,
            I => throttle_order_2
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__32526\,
            I => throttle_order_2
        );

    \I__6142\ : IoInMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32516\,
            I => \N__32512\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__32515\,
            I => \N__32509\
        );

    \I__6139\ : Span12Mux_s8_v
    port map (
            O => \N__32512\,
            I => \N__32506\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32503\
        );

    \I__6137\ : Odrv12
    port map (
            O => \N__32506\,
            I => ppm_output_c
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__32503\,
            I => ppm_output_c
        );

    \I__6135\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32495\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__32495\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__32492\,
            I => \N__32487\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32484\
        );

    \I__6131\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32481\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32478\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32473\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32481\,
            I => \N__32473\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32468\
        );

    \I__6126\ : Span4Mux_v
    port map (
            O => \N__32473\,
            I => \N__32468\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__32468\,
            I => throttle_order_10
        );

    \I__6124\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32460\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32457\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32454\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__32460\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32457\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32454\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32444\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32444\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32441\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32435\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__6113\ : Odrv4
    port map (
            O => \N__32432\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32429\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32426\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32420\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__32420\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__32417\,
            I => \N__32412\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32409\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__32415\,
            I => \N__32406\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32402\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32399\
        );

    \I__6103\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32394\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32405\,
            I => \N__32394\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32402\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6100\ : Odrv12
    port map (
            O => \N__32399\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32394\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__32387\,
            I => \N__32381\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32378\
        );

    \I__6096\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32375\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32370\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32370\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__32378\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__32375\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__32370\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__32363\,
            I => \N__32358\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32355\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32352\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32349\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32355\,
            I => \uart_drone.N_126_li\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32352\,
            I => \uart_drone.N_126_li\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32349\,
            I => \uart_drone.N_126_li\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32336\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__32341\,
            I => \N__32331\
        );

    \I__6081\ : CascadeMux
    port map (
            O => \N__32340\,
            I => \N__32328\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32325\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32322\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32317\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32317\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32314\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32311\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32325\,
            I => \uart_drone.N_143\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__32322\,
            I => \uart_drone.N_143\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32317\,
            I => \uart_drone.N_143\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__32314\,
            I => \uart_drone.N_143\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__32311\,
            I => \uart_drone.N_143\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32296\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32293\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32288\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32288\
        );

    \I__6065\ : Odrv12
    port map (
            O => \N__32288\,
            I => scaler_4_data_12
        );

    \I__6064\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__32282\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__32276\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__6060\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32270\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32266\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32263\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__32266\,
            I => \N__32258\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__32263\,
            I => \N__32258\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__32258\,
            I => scaler_4_data_8
        );

    \I__6054\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32252\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32246\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__32246\,
            I => \N__32242\
        );

    \I__6050\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32239\
        );

    \I__6049\ : Span4Mux_h
    port map (
            O => \N__32242\,
            I => \N__32234\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32234\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__32234\,
            I => scaler_4_data_7
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__32231\,
            I => \pid_front.un1_reset_i_a5_0_2_cascade_\
        );

    \I__6045\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__32225\,
            I => \pid_front.un1_reset_i_a5_0_3\
        );

    \I__6043\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32218\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32213\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__6040\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32207\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32204\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__32213\,
            I => \N__32201\
        );

    \I__6037\ : Span4Mux_v
    port map (
            O => \N__32210\,
            I => \N__32196\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__32207\,
            I => \N__32196\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__32204\,
            I => \pid_front.pid_preregZ0Z_1\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__32201\,
            I => \pid_front.pid_preregZ0Z_1\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__32196\,
            I => \pid_front.pid_preregZ0Z_1\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__32189\,
            I => \N__32185\
        );

    \I__6031\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32180\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32180\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32176\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__32179\,
            I => \N__32173\
        );

    \I__6027\ : Span4Mux_h
    port map (
            O => \N__32176\,
            I => \N__32169\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32166\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32163\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__32169\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__32166\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__32163\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__6021\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32153\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__32153\,
            I => \uart_pc.state_srsts_i_0_2\
        );

    \I__6019\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32143\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32140\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__32143\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__32140\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__32135\,
            I => \N__32132\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32127\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32122\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32130\,
            I => \N__32122\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__32127\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__32122\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32113\
        );

    \I__6007\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32110\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__32113\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32110\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__6004\ : CascadeMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32099\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__32099\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__32093\,
            I => \N__32089\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__32092\,
            I => \N__32086\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__32089\,
            I => \N__32082\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32077\
        );

    \I__5996\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32077\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__32082\,
            I => \uart_drone.N_152\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32077\,
            I => \uart_drone.N_152\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__32072\,
            I => \pid_front.N_533_cascade_\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32057\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32057\
        );

    \I__5990\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32057\
        );

    \I__5989\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32057\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__32057\,
            I => \pid_front.N_10_1\
        );

    \I__5987\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32051\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__32051\,
            I => \N__32048\
        );

    \I__5985\ : Span4Mux_v
    port map (
            O => \N__32048\,
            I => \N__32043\
        );

    \I__5984\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32038\
        );

    \I__5983\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32038\
        );

    \I__5982\ : Sp12to4
    port map (
            O => \N__32043\,
            I => \N__32033\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__32038\,
            I => \N__32033\
        );

    \I__5980\ : Odrv12
    port map (
            O => \N__32033\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32019\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32029\,
            I => \N__32001\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32028\,
            I => \N__32001\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32001\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32001\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32025\,
            I => \N__32001\
        );

    \I__5973\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32001\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32023\,
            I => \N__31998\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32022\,
            I => \N__31995\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__32019\,
            I => \N__31992\
        );

    \I__5969\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31989\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32017\,
            I => \N__31979\
        );

    \I__5967\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31979\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31979\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31976\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31971\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31971\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__31995\,
            I => \N__31965\
        );

    \I__5961\ : Span4Mux_v
    port map (
            O => \N__31992\,
            I => \N__31962\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31959\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31954\
        );

    \I__5958\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31954\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31951\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31943\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31943\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__31971\,
            I => \N__31940\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31933\
        );

    \I__5952\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31933\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31933\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__31965\,
            I => \N__31926\
        );

    \I__5949\ : Span4Mux_h
    port map (
            O => \N__31962\,
            I => \N__31926\
        );

    \I__5948\ : Span4Mux_h
    port map (
            O => \N__31959\,
            I => \N__31926\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31923\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31920\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__31950\,
            I => \N__31917\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__31949\,
            I => \N__31914\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__31948\,
            I => \N__31911\
        );

    \I__5942\ : Span4Mux_h
    port map (
            O => \N__31943\,
            I => \N__31907\
        );

    \I__5941\ : Span4Mux_h
    port map (
            O => \N__31940\,
            I => \N__31902\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31902\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__31926\,
            I => \N__31899\
        );

    \I__5938\ : Span4Mux_v
    port map (
            O => \N__31923\,
            I => \N__31896\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__31920\,
            I => \N__31893\
        );

    \I__5936\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31883\
        );

    \I__5935\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31883\
        );

    \I__5934\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31883\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31883\
        );

    \I__5932\ : Span4Mux_h
    port map (
            O => \N__31907\,
            I => \N__31880\
        );

    \I__5931\ : Span4Mux_v
    port map (
            O => \N__31902\,
            I => \N__31877\
        );

    \I__5930\ : Span4Mux_h
    port map (
            O => \N__31899\,
            I => \N__31870\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__31896\,
            I => \N__31870\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__31893\,
            I => \N__31870\
        );

    \I__5927\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31867\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__31883\,
            I => \pid_alt.N_72_i\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__31880\,
            I => \pid_alt.N_72_i\
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__31877\,
            I => \pid_alt.N_72_i\
        );

    \I__5923\ : Odrv4
    port map (
            O => \N__31870\,
            I => \pid_alt.N_72_i\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31867\,
            I => \pid_alt.N_72_i\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31856\,
            I => \N__31844\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31844\
        );

    \I__5919\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31844\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31839\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31834\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31834\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31844\,
            I => \N__31830\
        );

    \I__5914\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31825\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31842\,
            I => \N__31825\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31839\,
            I => \N__31820\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31820\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31817\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__31830\,
            I => \pid_alt.N_299\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31825\,
            I => \pid_alt.N_299\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__31820\,
            I => \pid_alt.N_299\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__31817\,
            I => \pid_alt.N_299\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31804\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__31807\,
            I => \N__31800\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31797\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31794\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31791\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__31797\,
            I => \N__31784\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31784\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__31791\,
            I => \N__31784\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__31784\,
            I => \N__31781\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__31781\,
            I => \pid_alt.pid_preregZ0Z_7\
        );

    \I__5895\ : SRMux
    port map (
            O => \N__31778\,
            I => \N__31775\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31775\,
            I => \N__31771\
        );

    \I__5893\ : SRMux
    port map (
            O => \N__31774\,
            I => \N__31765\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__31771\,
            I => \N__31762\
        );

    \I__5891\ : SRMux
    port map (
            O => \N__31770\,
            I => \N__31759\
        );

    \I__5890\ : SRMux
    port map (
            O => \N__31769\,
            I => \N__31756\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31753\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31765\,
            I => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__31762\,
            I => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__31759\,
            I => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31756\,
            I => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__31753\,
            I => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\
        );

    \I__5883\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31739\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31739\,
            I => \N__31736\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__31736\,
            I => \ppm_encoder_1.N_292\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__31733\,
            I => \uart_drone.un1_state_7_0_cascade_\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__31730\,
            I => \uart_drone.N_152_cascade_\
        );

    \I__5878\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31715\
        );

    \I__5877\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31715\
        );

    \I__5876\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31715\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31715\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31715\,
            I => \N__31710\
        );

    \I__5873\ : InMux
    port map (
            O => \N__31714\,
            I => \N__31707\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31704\
        );

    \I__5871\ : Span4Mux_v
    port map (
            O => \N__31710\,
            I => \N__31695\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31695\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31692\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31703\,
            I => \N__31689\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31682\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31682\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31682\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__31695\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__31692\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__31689\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__31682\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__31673\,
            I => \N__31670\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31667\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31667\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__31664\,
            I => \N__31658\
        );

    \I__5856\ : CascadeMux
    port map (
            O => \N__31663\,
            I => \N__31655\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31651\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31642\
        );

    \I__5853\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31642\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31642\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31642\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31637\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31634\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31631\
        );

    \I__5847\ : InMux
    port map (
            O => \N__31640\,
            I => \N__31628\
        );

    \I__5846\ : Span12Mux_v
    port map (
            O => \N__31637\,
            I => \N__31623\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__31634\,
            I => \N__31616\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31631\,
            I => \N__31616\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31628\,
            I => \N__31616\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31611\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31611\
        );

    \I__5840\ : Odrv12
    port map (
            O => \N__31623\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__31616\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31611\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31604\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31601\,
            I => \ppm_encoder_1.un1_throttle_cry_13\
        );

    \I__5835\ : CEMux
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31592\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__31592\,
            I => \N__31589\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__31589\,
            I => \pid_alt.N_72_i_1\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31583\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31583\,
            I => \N__31580\
        );

    \I__5829\ : Span4Mux_v
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__5828\ : Odrv4
    port map (
            O => \N__31577\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31567\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31564\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31560\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31557\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31554\
        );

    \I__5821\ : Span4Mux_h
    port map (
            O => \N__31560\,
            I => \N__31551\
        );

    \I__5820\ : Span4Mux_h
    port map (
            O => \N__31557\,
            I => \N__31546\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31546\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__31551\,
            I => \N__31543\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__31546\,
            I => \N__31540\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__31543\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__5815\ : Odrv4
    port map (
            O => \N__31540\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__5813\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31525\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31522\
        );

    \I__5810\ : Span4Mux_v
    port map (
            O => \N__31525\,
            I => \N__31517\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31522\,
            I => \N__31517\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__31517\,
            I => \N__31513\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31510\
        );

    \I__5806\ : Span4Mux_h
    port map (
            O => \N__31513\,
            I => \N__31507\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31504\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__31507\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__31504\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31496\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31496\,
            I => \N__31492\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31489\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__31492\,
            I => \N__31484\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31489\,
            I => \N__31484\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__31484\,
            I => \N__31480\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31483\,
            I => \N__31477\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__31480\,
            I => \N__31474\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31471\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__31474\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__31471\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31462\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31459\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31462\,
            I => \N__31456\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31459\,
            I => \N__31453\
        );

    \I__5787\ : Span4Mux_v
    port map (
            O => \N__31456\,
            I => \N__31450\
        );

    \I__5786\ : Odrv12
    port map (
            O => \N__31453\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__31450\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31433\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31433\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31433\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31433\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31433\,
            I => \pid_alt.N_472_1\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31430\,
            I => \ppm_encoder_1.un1_throttle_cry_3\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31427\,
            I => \ppm_encoder_1.un1_throttle_cry_4\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31424\,
            I => \ppm_encoder_1.un1_throttle_cry_5\
        );

    \I__5776\ : InMux
    port map (
            O => \N__31421\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31418\,
            I => \bfn_12_13_0_\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__31415\,
            I => \N__31411\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31408\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31404\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__31408\,
            I => \N__31401\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31398\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31404\,
            I => throttle_order_9
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__31401\,
            I => throttle_order_9
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31398\,
            I => throttle_order_9
        );

    \I__5766\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__31385\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31382\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31379\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31376\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31373\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31370\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31367\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31364\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__5756\ : InMux
    port map (
            O => \N__31361\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31355\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__31352\,
            I => scaler_4_data_14
        );

    \I__5752\ : InMux
    port map (
            O => \N__31349\,
            I => \bfn_12_11_0_\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31346\,
            I => \ppm_encoder_1.un1_throttle_cry_0\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31343\,
            I => \ppm_encoder_1.un1_throttle_cry_1\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31340\,
            I => \ppm_encoder_1.un1_throttle_cry_2\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \uart_drone.timer_Count_RNO_0_0_1_cascade_\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31329\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31326\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31323\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__31329\,
            I => \N__31320\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31326\,
            I => \N__31317\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__31323\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__31320\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__31317\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__5739\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31307\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__31307\,
            I => \N__31300\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31297\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31294\
        );

    \I__5735\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31286\
        );

    \I__5734\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31286\
        );

    \I__5733\ : Span4Mux_v
    port map (
            O => \N__31300\,
            I => \N__31279\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__31297\,
            I => \N__31279\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31294\,
            I => \N__31279\
        );

    \I__5730\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31272\
        );

    \I__5729\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31272\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31272\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__31286\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__31279\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31272\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__5724\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31262\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31257\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31254\
        );

    \I__5721\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31251\
        );

    \I__5720\ : Span4Mux_v
    port map (
            O => \N__31257\,
            I => \N__31246\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31246\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__31251\,
            I => \uart_pc.N_126_li\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__31246\,
            I => \uart_pc.N_126_li\
        );

    \I__5716\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31217\
        );

    \I__5715\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31217\
        );

    \I__5714\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31217\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31217\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31217\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31217\
        );

    \I__5710\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31217\
        );

    \I__5709\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31217\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31214\
        );

    \I__5707\ : Odrv4
    port map (
            O => \N__31214\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__5706\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31208\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31205\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__31205\,
            I => \N__31201\
        );

    \I__5703\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31198\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__31201\,
            I => \N__31195\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31198\,
            I => \N__31192\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__31195\,
            I => scaler_4_data_6
        );

    \I__5699\ : Odrv4
    port map (
            O => \N__31192\,
            I => scaler_4_data_6
        );

    \I__5698\ : InMux
    port map (
            O => \N__31187\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__5697\ : InMux
    port map (
            O => \N__31184\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__5696\ : InMux
    port map (
            O => \N__31181\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__31178\,
            I => \N__31174\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31177\,
            I => \N__31171\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31168\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__31171\,
            I => \N__31164\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31160\
        );

    \I__5690\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31157\
        );

    \I__5689\ : Span4Mux_v
    port map (
            O => \N__31164\,
            I => \N__31154\
        );

    \I__5688\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31151\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__31160\,
            I => \N__31148\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31144\
        );

    \I__5685\ : Sp12to4
    port map (
            O => \N__31154\,
            I => \N__31139\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31151\,
            I => \N__31139\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__31148\,
            I => \N__31136\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31133\
        );

    \I__5681\ : Sp12to4
    port map (
            O => \N__31144\,
            I => \N__31128\
        );

    \I__5680\ : Span12Mux_h
    port map (
            O => \N__31139\,
            I => \N__31128\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__31136\,
            I => \N__31125\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31133\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__5677\ : Odrv12
    port map (
            O => \N__31128\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__31125\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__5675\ : IoInMux
    port map (
            O => \N__31118\,
            I => \N__31115\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__31115\,
            I => \pid_alt.state_0_0\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__31112\,
            I => \N__31105\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \N__31102\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__31110\,
            I => \N__31095\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \N__31092\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31085\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31085\
        );

    \I__5667\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31085\
        );

    \I__5666\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31082\
        );

    \I__5665\ : InMux
    port map (
            O => \N__31100\,
            I => \N__31079\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31074\
        );

    \I__5663\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31074\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31069\
        );

    \I__5661\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31069\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31066\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__31082\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__31079\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__31074\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__31069\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__31066\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__5654\ : IoInMux
    port map (
            O => \N__31055\,
            I => \N__31051\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31054\,
            I => \N__31043\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31039\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__31050\,
            I => \N__31036\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__31049\,
            I => \N__31033\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__31048\,
            I => \N__31030\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__31047\,
            I => \N__31027\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__31046\,
            I => \N__31022\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31018\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31015\
        );

    \I__5644\ : Span4Mux_s3_v
    port map (
            O => \N__31039\,
            I => \N__31012\
        );

    \I__5643\ : InMux
    port map (
            O => \N__31036\,
            I => \N__30996\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31033\,
            I => \N__30996\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31030\,
            I => \N__30996\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31027\,
            I => \N__30996\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31026\,
            I => \N__30996\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31025\,
            I => \N__30996\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31022\,
            I => \N__30991\
        );

    \I__5636\ : InMux
    port map (
            O => \N__31021\,
            I => \N__30991\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__31018\,
            I => \N__30986\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31015\,
            I => \N__30986\
        );

    \I__5633\ : Span4Mux_v
    port map (
            O => \N__31012\,
            I => \N__30983\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31011\,
            I => \N__30980\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31010\,
            I => \N__30975\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31009\,
            I => \N__30975\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30970\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30991\,
            I => \N__30970\
        );

    \I__5627\ : Span4Mux_v
    port map (
            O => \N__30986\,
            I => \N__30967\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__30983\,
            I => \debug_CH0_16A_c\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__30980\,
            I => \debug_CH0_16A_c\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30975\,
            I => \debug_CH0_16A_c\
        );

    \I__5623\ : Odrv12
    port map (
            O => \N__30970\,
            I => \debug_CH0_16A_c\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__30967\,
            I => \debug_CH0_16A_c\
        );

    \I__5621\ : CascadeMux
    port map (
            O => \N__30956\,
            I => \uart_drone.state_srsts_0_0_0_cascade_\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__30953\,
            I => \N__30950\
        );

    \I__5619\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30947\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30944\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__30944\,
            I => \N__30940\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30937\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__30940\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__30937\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__30929\,
            I => \N__30926\
        );

    \I__5611\ : Odrv12
    port map (
            O => \N__30926\,
            I => \pid_side.un1_pid_prereg_cry_2_THRU_CO\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30919\
        );

    \I__5609\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__30919\,
            I => \N__30913\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30910\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__30913\,
            I => \N__30906\
        );

    \I__5605\ : Span4Mux_v
    port map (
            O => \N__30910\,
            I => \N__30903\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30900\
        );

    \I__5603\ : Sp12to4
    port map (
            O => \N__30906\,
            I => \N__30895\
        );

    \I__5602\ : Sp12to4
    port map (
            O => \N__30903\,
            I => \N__30895\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__30900\,
            I => \pid_side.error_p_regZ0Z_16\
        );

    \I__5600\ : Odrv12
    port map (
            O => \N__30895\,
            I => \pid_side.error_p_regZ0Z_16\
        );

    \I__5599\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30887\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__30887\,
            I => \N__30884\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__30884\,
            I => \N__30881\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__30881\,
            I => \pid_side.un1_pid_prereg_cry_15_THRU_CO\
        );

    \I__5595\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30875\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30872\
        );

    \I__5593\ : Odrv12
    port map (
            O => \N__30872\,
            I => \pid_side.un1_pid_prereg_cry_4_THRU_CO\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30866\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30862\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30859\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__30862\,
            I => \N__30854\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30859\,
            I => \N__30854\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__30854\,
            I => \N__30850\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30847\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__30850\,
            I => \N__30844\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__30847\,
            I => \pid_side.error_p_regZ0Z_5\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__30844\,
            I => \pid_side.error_p_regZ0Z_5\
        );

    \I__5582\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30836\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__30836\,
            I => \N__30833\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__30833\,
            I => \N__30829\
        );

    \I__5579\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30826\
        );

    \I__5578\ : Sp12to4
    port map (
            O => \N__30829\,
            I => \N__30820\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30820\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30817\
        );

    \I__5575\ : Span12Mux_h
    port map (
            O => \N__30820\,
            I => \N__30814\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30817\,
            I => \pid_side.error_p_regZ0Z_13\
        );

    \I__5573\ : Odrv12
    port map (
            O => \N__30814\,
            I => \pid_side.error_p_regZ0Z_13\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30806\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__30806\,
            I => \N__30803\
        );

    \I__5570\ : Span4Mux_h
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__30800\,
            I => \pid_side.un1_pid_prereg_cry_12_THRU_CO\
        );

    \I__5568\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30793\
        );

    \I__5567\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30790\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__30793\,
            I => \N__30787\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__30790\,
            I => \N__30784\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__30787\,
            I => \N__30781\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__30784\,
            I => \N__30778\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__30781\,
            I => \N__30775\
        );

    \I__5561\ : Span4Mux_h
    port map (
            O => \N__30778\,
            I => \N__30772\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__30775\,
            I => \N__30769\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__30772\,
            I => \N__30766\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__30769\,
            I => \N__30761\
        );

    \I__5557\ : Span4Mux_h
    port map (
            O => \N__30766\,
            I => \N__30761\
        );

    \I__5556\ : Odrv4
    port map (
            O => \N__30761\,
            I => xy_kp_1
        );

    \I__5555\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30754\
        );

    \I__5554\ : InMux
    port map (
            O => \N__30757\,
            I => \N__30751\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__30754\,
            I => \N__30748\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30745\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__30748\,
            I => \N__30742\
        );

    \I__5550\ : Span4Mux_s1_h
    port map (
            O => \N__30745\,
            I => \N__30739\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__30742\,
            I => \N__30736\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__30739\,
            I => \N__30733\
        );

    \I__5547\ : Span4Mux_h
    port map (
            O => \N__30736\,
            I => \N__30730\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__30733\,
            I => \N__30727\
        );

    \I__5545\ : Span4Mux_h
    port map (
            O => \N__30730\,
            I => \N__30722\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__30727\,
            I => \N__30722\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__30722\,
            I => xy_kp_7
        );

    \I__5542\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30716\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__30716\,
            I => \pid_alt.un1_reset_i_a5_1_10_8\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30713\,
            I => \N__30710\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__5538\ : Odrv12
    port map (
            O => \N__30707\,
            I => \pid_alt.un1_reset_i_a5_1_10_9\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__30704\,
            I => \pid_alt.un1_reset_i_a5_0_6_cascade_\
        );

    \I__5536\ : CascadeMux
    port map (
            O => \N__30701\,
            I => \pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_\
        );

    \I__5535\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30695\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__30689\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30682\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30679\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30682\,
            I => \pid_alt.N_530\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__30679\,
            I => \pid_alt.N_530\
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30670\,
            I => \N__30665\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__30662\,
            I => \pid_alt.N_535\
        );

    \I__5522\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30652\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30652\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30649\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__30652\,
            I => \N__30645\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30642\
        );

    \I__5517\ : CascadeMux
    port map (
            O => \N__30648\,
            I => \N__30639\
        );

    \I__5516\ : Span4Mux_v
    port map (
            O => \N__30645\,
            I => \N__30633\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__30642\,
            I => \N__30633\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30630\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30627\
        );

    \I__5512\ : Sp12to4
    port map (
            O => \N__30633\,
            I => \N__30620\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30620\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30620\
        );

    \I__5509\ : Odrv12
    port map (
            O => \N__30620\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__30617\,
            I => \pid_alt.N_535_cascade_\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30611\,
            I => \N__30606\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30610\,
            I => \N__30603\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30600\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30606\,
            I => \N__30597\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30603\,
            I => \N__30594\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30600\,
            I => \N__30591\
        );

    \I__5500\ : Span4Mux_h
    port map (
            O => \N__30597\,
            I => \N__30587\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__30594\,
            I => \N__30584\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__30591\,
            I => \N__30581\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30578\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__30587\,
            I => \N__30575\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__30584\,
            I => \N__30572\
        );

    \I__5494\ : Span4Mux_h
    port map (
            O => \N__30581\,
            I => \N__30567\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30578\,
            I => \N__30567\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30575\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__30572\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__5490\ : Odrv4
    port map (
            O => \N__30567\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__5489\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30557\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30557\,
            I => \N__30554\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__30554\,
            I => \N__30551\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__30551\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30544\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30540\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30537\
        );

    \I__5482\ : CascadeMux
    port map (
            O => \N__30543\,
            I => \N__30533\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30530\
        );

    \I__5480\ : Span4Mux_v
    port map (
            O => \N__30537\,
            I => \N__30527\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30524\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30521\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__30530\,
            I => \N__30518\
        );

    \I__5476\ : Sp12to4
    port map (
            O => \N__30527\,
            I => \N__30511\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30511\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30511\
        );

    \I__5473\ : Odrv4
    port map (
            O => \N__30518\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__5472\ : Odrv12
    port map (
            O => \N__30511\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30500\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30500\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__30500\,
            I => \N__30496\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30493\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__30496\,
            I => \N__30485\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30493\,
            I => \N__30485\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30480\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30480\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30477\
        );

    \I__5462\ : Span4Mux_h
    port map (
            O => \N__30485\,
            I => \N__30474\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__30480\,
            I => \N__30469\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30477\,
            I => \N__30469\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__30474\,
            I => \N__30466\
        );

    \I__5458\ : Odrv12
    port map (
            O => \N__30469\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__30466\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__30461\,
            I => \N__30455\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__30460\,
            I => \N__30452\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30448\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30443\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30443\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30438\
        );

    \I__5450\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30438\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30435\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30432\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30429\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__30435\,
            I => \N__30426\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__30432\,
            I => \N__30423\
        );

    \I__5444\ : Span12Mux_v
    port map (
            O => \N__30429\,
            I => \N__30420\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__30426\,
            I => \N__30415\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__30423\,
            I => \N__30415\
        );

    \I__5441\ : Odrv12
    port map (
            O => \N__30420\,
            I => \pid_alt.pid_preregZ0Z_24\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__30415\,
            I => \pid_alt.pid_preregZ0Z_24\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30403\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30403\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30408\,
            I => \N__30400\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__30403\,
            I => \N__30396\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30400\,
            I => \N__30393\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30390\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__30396\,
            I => \N__30383\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__30393\,
            I => \N__30383\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30390\,
            I => \N__30383\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__30380\,
            I => \pid_alt.N_551\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30374\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5426\ : Odrv12
    port map (
            O => \N__30371\,
            I => \pid_side.un1_pid_prereg_cry_6_THRU_CO\
        );

    \I__5425\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30365\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__30362\,
            I => \N__30358\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30355\
        );

    \I__5421\ : Span4Mux_h
    port map (
            O => \N__30358\,
            I => \N__30349\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30349\
        );

    \I__5419\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30346\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__30349\,
            I => \N__30343\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30346\,
            I => \N__30338\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__30343\,
            I => \N__30338\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__30338\,
            I => \pid_side.error_p_regZ0Z_7\
        );

    \I__5414\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30332\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30329\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__30329\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30323\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30323\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30317\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30317\,
            I => \uart_drone.data_Auxce_0_0_4\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30311\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__30311\,
            I => \pid_alt.un1_reset_i_a5_0_6_3\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30302\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__30299\,
            I => \N__30295\
        );

    \I__5401\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30292\
        );

    \I__5400\ : Span4Mux_v
    port map (
            O => \N__30295\,
            I => \N__30287\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30287\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__30287\,
            I => \N__30284\
        );

    \I__5397\ : Span4Mux_h
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__30281\,
            I => \pid_alt.N_306_5\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__30278\,
            I => \pid_alt.un1_reset_i_a5_0_6_2_cascade_\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30271\
        );

    \I__5393\ : InMux
    port map (
            O => \N__30274\,
            I => \N__30268\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30271\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30268\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__30263\,
            I => \N__30259\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30262\,
            I => \N__30256\
        );

    \I__5388\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30253\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__30256\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30253\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30244\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30241\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30244\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__30241\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30232\
        );

    \I__5380\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30229\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__30232\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30229\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__5377\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30220\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30217\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30220\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__30217\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__30212\,
            I => \N__30208\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30205\
        );

    \I__5371\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30202\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__30205\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30202\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__5368\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30193\
        );

    \I__5367\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30190\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__30193\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30190\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30182\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30177\
        );

    \I__5362\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30172\
        );

    \I__5361\ : InMux
    port map (
            O => \N__30180\,
            I => \N__30172\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__30177\,
            I => \N__30167\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30167\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__30164\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__5356\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__30158\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__30155\,
            I => \uart_pc.N_152_cascade_\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__30152\,
            I => \N__30148\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30145\
        );

    \I__5351\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30141\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__30145\,
            I => \N__30133\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30130\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30141\,
            I => \N__30127\
        );

    \I__5347\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30124\
        );

    \I__5346\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30121\
        );

    \I__5345\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30114\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30114\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30136\,
            I => \N__30114\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__30133\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30130\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__30127\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__30124\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__30121\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__30114\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__30101\,
            I => \uart_pc.CO0_cascade_\
        );

    \I__5335\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30089\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30089\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30089\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30085\
        );

    \I__5331\ : InMux
    port map (
            O => \N__30088\,
            I => \N__30082\
        );

    \I__5330\ : Odrv4
    port map (
            O => \N__30085\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__30082\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__5328\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30071\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30071\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30071\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__5325\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30065\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__30065\,
            I => \N__30062\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__30059\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__30056\,
            I => \N__30053\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30047\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30047\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30047\,
            I => \N__30042\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__30046\,
            I => \N__30039\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__30045\,
            I => \N__30033\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__30042\,
            I => \N__30027\
        );

    \I__5314\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30020\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30020\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30020\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30011\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30011\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30011\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30031\,
            I => \N__30011\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30008\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__30027\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__30020\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__30011\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__30008\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29992\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29992\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__29997\,
            I => \N__29985\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__29992\,
            I => \N__29980\
        );

    \I__5298\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29973\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29973\
        );

    \I__5296\ : InMux
    port map (
            O => \N__29989\,
            I => \N__29973\
        );

    \I__5295\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29966\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29966\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29966\
        );

    \I__5292\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29963\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__29980\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__29973\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__29966\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29963\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__5287\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29948\
        );

    \I__5286\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29943\
        );

    \I__5285\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29943\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__29951\,
            I => \N__29937\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__29948\,
            I => \N__29928\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29928\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29921\
        );

    \I__5280\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29921\
        );

    \I__5279\ : InMux
    port map (
            O => \N__29940\,
            I => \N__29921\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29912\
        );

    \I__5277\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29912\
        );

    \I__5276\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29912\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29912\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29909\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__29928\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__29921\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__29912\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__29909\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__5269\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29897\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \N__29890\
        );

    \I__5266\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29887\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29884\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__29887\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__29884\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29876\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29871\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29866\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29866\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__29871\,
            I => \N__29863\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29860\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__29863\,
            I => \N__29857\
        );

    \I__5255\ : Span4Mux_v
    port map (
            O => \N__29860\,
            I => \N__29854\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__29857\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__29854\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29846\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__29843\,
            I => \uart_drone_sync.aux_3__0__0_0\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__29840\,
            I => \uart_drone.timer_Count_0_sqmuxa_cascade_\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__29837\,
            I => \uart_pc.N_145_cascade_\
        );

    \I__5247\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__29831\,
            I => \uart_pc.N_144_1\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__29828\,
            I => \uart_pc.N_144_1_cascade_\
        );

    \I__5244\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__29822\,
            I => \N__29815\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29812\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29807\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29807\
        );

    \I__5239\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29804\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__29815\,
            I => \uart_pc.N_143\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__29812\,
            I => \uart_pc.N_143\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__29807\,
            I => \uart_pc.N_143\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29804\,
            I => \uart_pc.N_143\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29795\,
            I => \N__29792\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__29792\,
            I => \N__29784\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29781\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29778\
        );

    \I__5230\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29773\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29773\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29770\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__29784\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29781\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__29778\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__29773\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29770\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__5222\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29756\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29753\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__5219\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__29747\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29744\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29741\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__29735\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__29726\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29718\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__29722\,
            I => \N__29714\
        );

    \I__5208\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29711\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29718\,
            I => \N__29708\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29703\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29703\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29711\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__29708\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29703\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__5201\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29693\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29686\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__29692\,
            I => \N__29683\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29680\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__29690\,
            I => \N__29677\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__29689\,
            I => \N__29674\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__29686\,
            I => \N__29671\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29668\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29665\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29660\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29674\,
            I => \N__29660\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__29671\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__29668\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__5188\ : Odrv4
    port map (
            O => \N__29665\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29660\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__29651\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\
        );

    \I__5185\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29644\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29644\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__29641\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29629\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29626\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__29629\,
            I => \N__29623\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29626\,
            I => \N__29620\
        );

    \I__5176\ : Span4Mux_h
    port map (
            O => \N__29623\,
            I => \N__29615\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__29620\,
            I => \N__29615\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__29615\,
            I => \drone_H_disp_side_13\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__29612\,
            I => \N__29608\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29603\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29603\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__29600\,
            I => \N__29597\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__29597\,
            I => \N__29594\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__29594\,
            I => \drone_H_disp_side_14\
        );

    \I__5166\ : CEMux
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29588\,
            I => \N__29584\
        );

    \I__5164\ : CEMux
    port map (
            O => \N__29587\,
            I => \N__29581\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__29584\,
            I => \N__29575\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29575\
        );

    \I__5161\ : CEMux
    port map (
            O => \N__29580\,
            I => \N__29572\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__29569\,
            I => \N__29563\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__29566\,
            I => \N__29560\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__29563\,
            I => \N__29557\
        );

    \I__5155\ : Span4Mux_v
    port map (
            O => \N__29560\,
            I => \N__29554\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__29557\,
            I => \dron_frame_decoder_1.N_739_0\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29554\,
            I => \dron_frame_decoder_1.N_739_0\
        );

    \I__5152\ : CascadeMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29543\,
            I => \N__29539\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29542\,
            I => \N__29535\
        );

    \I__5148\ : Span12Mux_s10_h
    port map (
            O => \N__29539\,
            I => \N__29532\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29529\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__29535\,
            I => \drone_H_disp_side_12\
        );

    \I__5145\ : Odrv12
    port map (
            O => \N__29532\,
            I => \drone_H_disp_side_12\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29529\,
            I => \drone_H_disp_side_12\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29513\
        );

    \I__5140\ : Odrv12
    port map (
            O => \N__29513\,
            I => \drone_H_disp_side_i_12\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29507\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29507\,
            I => \drone_H_disp_front_3\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29500\
        );

    \I__5136\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29497\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29494\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29497\,
            I => \N__29491\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__29494\,
            I => \N__29488\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__5131\ : Sp12to4
    port map (
            O => \N__29488\,
            I => \N__29482\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__29485\,
            I => \N__29479\
        );

    \I__5129\ : Span12Mux_s3_h
    port map (
            O => \N__29482\,
            I => \N__29476\
        );

    \I__5128\ : Sp12to4
    port map (
            O => \N__29479\,
            I => \N__29473\
        );

    \I__5127\ : Span12Mux_h
    port map (
            O => \N__29476\,
            I => \N__29470\
        );

    \I__5126\ : Odrv12
    port map (
            O => \N__29473\,
            I => xy_kp_3
        );

    \I__5125\ : Odrv12
    port map (
            O => \N__29470\,
            I => xy_kp_3
        );

    \I__5124\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__29456\,
            I => \uart_drone_sync.aux_2__0__0_0\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__29453\,
            I => \pid_alt.un1_reset_i_a5_1_10_5_cascade_\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29445\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29440\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29440\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29437\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__29437\,
            I => \N__29431\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__5112\ : Span4Mux_h
    port map (
            O => \N__29431\,
            I => \N__29425\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__29428\,
            I => \N__29422\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__29425\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__5109\ : Odrv4
    port map (
            O => \N__29422\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29414\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__5106\ : Span4Mux_v
    port map (
            O => \N__29411\,
            I => \N__29408\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__29408\,
            I => \pid_side.un1_pid_prereg_cry_9_THRU_CO\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29401\
        );

    \I__5103\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29398\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__29401\,
            I => \N__29395\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__29398\,
            I => \N__29392\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__29395\,
            I => \N__29388\
        );

    \I__5099\ : Span12Mux_h
    port map (
            O => \N__29392\,
            I => \N__29385\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29382\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__29388\,
            I => \N__29379\
        );

    \I__5096\ : Odrv12
    port map (
            O => \N__29385\,
            I => \pid_side.error_p_regZ0Z_10\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29382\,
            I => \pid_side.error_p_regZ0Z_10\
        );

    \I__5094\ : Odrv4
    port map (
            O => \N__29379\,
            I => \pid_side.error_p_regZ0Z_10\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__29372\,
            I => \pid_side.un1_reset_i_a2_3_cascade_\
        );

    \I__5092\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29365\
        );

    \I__5091\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29365\,
            I => \pid_side.pid_preregZ0Z_18\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__29362\,
            I => \pid_side.pid_preregZ0Z_18\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29353\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29350\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__29353\,
            I => \pid_side.pid_preregZ0Z_17\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__29350\,
            I => \pid_side.pid_preregZ0Z_17\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__29345\,
            I => \N__29341\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29338\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29335\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__29338\,
            I => \pid_side.pid_preregZ0Z_19\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29335\,
            I => \pid_side.pid_preregZ0Z_19\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__29330\,
            I => \N__29327\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29323\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29320\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__29323\,
            I => \pid_side.pid_preregZ0Z_20\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__29320\,
            I => \pid_side.pid_preregZ0Z_20\
        );

    \I__5074\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29311\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29308\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29311\,
            I => \N__29305\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29308\,
            I => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\
        );

    \I__5070\ : Odrv12
    port map (
            O => \N__29305\,
            I => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29294\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29294\,
            I => \drone_H_disp_side_11\
        );

    \I__5066\ : CEMux
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__5064\ : Span4Mux_v
    port map (
            O => \N__29285\,
            I => \N__29281\
        );

    \I__5063\ : CEMux
    port map (
            O => \N__29284\,
            I => \N__29278\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__29281\,
            I => \N__29275\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__29275\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__5059\ : Odrv12
    port map (
            O => \N__29272\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__5058\ : SRMux
    port map (
            O => \N__29267\,
            I => \N__29263\
        );

    \I__5057\ : SRMux
    port map (
            O => \N__29266\,
            I => \N__29260\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29257\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29260\,
            I => \N__29254\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__29257\,
            I => \N__29251\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__29254\,
            I => \N__29248\
        );

    \I__5052\ : Odrv4
    port map (
            O => \N__29251\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__29248\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__29243\,
            I => \N__29240\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29235\
        );

    \I__5048\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29232\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29229\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__29235\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__29232\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__29229\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__29222\,
            I => \N__29217\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29214\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29207\
        );

    \I__5040\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29200\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29197\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29192\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29187\
        );

    \I__5036\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29187\
        );

    \I__5035\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29184\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29181\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29178\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29171\
        );

    \I__5031\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29171\
        );

    \I__5030\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29171\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29166\
        );

    \I__5028\ : Span4Mux_v
    port map (
            O => \N__29197\,
            I => \N__29166\
        );

    \I__5027\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29161\
        );

    \I__5026\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29161\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__29192\,
            I => uart_drone_data_rdy
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__29187\,
            I => uart_drone_data_rdy
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__29184\,
            I => uart_drone_data_rdy
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__29181\,
            I => uart_drone_data_rdy
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__29178\,
            I => uart_drone_data_rdy
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29171\,
            I => uart_drone_data_rdy
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__29166\,
            I => uart_drone_data_rdy
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29161\,
            I => uart_drone_data_rdy
        );

    \I__5017\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29136\
        );

    \I__5015\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29133\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29130\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__29136\,
            I => \N__29127\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29124\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__29130\,
            I => \N__29121\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__29127\,
            I => \N__29116\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__29124\,
            I => \N__29116\
        );

    \I__5008\ : Span12Mux_h
    port map (
            O => \N__29121\,
            I => \N__29113\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__29116\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__5006\ : Odrv12
    port map (
            O => \N__29113\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__29108\,
            I => \pid_alt.un1_reset_i_a2_3_cascade_\
        );

    \I__5004\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29102\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29102\,
            I => \N__29099\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__29099\,
            I => \N__29094\
        );

    \I__5001\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29089\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29089\
        );

    \I__4999\ : Sp12to4
    port map (
            O => \N__29094\,
            I => \N__29084\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29084\
        );

    \I__4997\ : Odrv12
    port map (
            O => \N__29084\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__4996\ : CascadeMux
    port map (
            O => \N__29081\,
            I => \N__29078\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29078\,
            I => \N__29075\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29071\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29062\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__29065\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29062\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__4988\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29054\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N__29051\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__29051\,
            I => \N__29048\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__29048\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__4984\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29042\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__29033\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__29030\,
            I => \N__29025\
        );

    \I__4978\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29022\
        );

    \I__4977\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29017\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29017\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__29022\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__29017\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__29012\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__4972\ : InMux
    port map (
            O => \N__29009\,
            I => \N__29004\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__29008\,
            I => \N__29001\
        );

    \I__4970\ : InMux
    port map (
            O => \N__29007\,
            I => \N__28997\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__28994\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28989\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28989\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__28997\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__28994\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28989\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28978\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28975\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28969\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__28975\,
            I => \N__28969\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__28974\,
            I => \N__28965\
        );

    \I__4958\ : Span4Mux_v
    port map (
            O => \N__28969\,
            I => \N__28962\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__4956\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28956\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__28962\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28959\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__28956\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__4952\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28945\
        );

    \I__4951\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28942\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28939\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28934\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__28939\,
            I => \N__28931\
        );

    \I__4947\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28928\
        );

    \I__4946\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28925\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__28934\,
            I => \frame_decoder_CH4data_0\
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__28931\,
            I => \frame_decoder_CH4data_0\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__28928\,
            I => \frame_decoder_CH4data_0\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__28925\,
            I => \frame_decoder_CH4data_0\
        );

    \I__4941\ : CEMux
    port map (
            O => \N__28916\,
            I => \N__28913\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28908\
        );

    \I__4939\ : CEMux
    port map (
            O => \N__28912\,
            I => \N__28905\
        );

    \I__4938\ : CEMux
    port map (
            O => \N__28911\,
            I => \N__28902\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__28908\,
            I => \N__28897\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28897\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__28902\,
            I => \N__28894\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__28897\,
            I => \N__28891\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__28894\,
            I => \N__28888\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__28891\,
            I => \N__28885\
        );

    \I__4931\ : Span4Mux_v
    port map (
            O => \N__28888\,
            I => \N__28882\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__28885\,
            I => \N__28879\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__28882\,
            I => \scaler_4.debug_CH3_20A_c_0\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__28879\,
            I => \scaler_4.debug_CH3_20A_c_0\
        );

    \I__4927\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28870\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__28873\,
            I => \N__28867\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__4924\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28861\
        );

    \I__4923\ : Odrv12
    port map (
            O => \N__28864\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__28861\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28849\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__28852\,
            I => \N__28846\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__28849\,
            I => \N__28843\
        );

    \I__4917\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28840\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__28843\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__28840\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__4914\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28832\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28832\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__4912\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28825\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__28828\,
            I => \N__28822\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28819\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28816\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__28819\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28816\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__4906\ : CEMux
    port map (
            O => \N__28811\,
            I => \N__28808\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__28808\,
            I => \pid_alt.state_1_0_0\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__28805\,
            I => \uart_pc.state_srsts_0_0_0_cascade_\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__28802\,
            I => \uart_pc.N_143_cascade_\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__28796\,
            I => \N__28793\
        );

    \I__4900\ : Span4Mux_h
    port map (
            O => \N__28793\,
            I => \N__28788\
        );

    \I__4899\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28783\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28783\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__28788\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28783\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__28778\,
            I => \uart_pc.data_rdyc_1_cascade_\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28770\
        );

    \I__4893\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28766\
        );

    \I__4892\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28763\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__28770\,
            I => \N__28760\
        );

    \I__4890\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28757\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28753\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__28763\,
            I => \N__28750\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__28760\,
            I => \N__28745\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28745\
        );

    \I__4885\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28742\
        );

    \I__4884\ : Span4Mux_v
    port map (
            O => \N__28753\,
            I => \N__28736\
        );

    \I__4883\ : Span4Mux_v
    port map (
            O => \N__28750\,
            I => \N__28736\
        );

    \I__4882\ : Span4Mux_h
    port map (
            O => \N__28745\,
            I => \N__28731\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28742\,
            I => \N__28731\
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__28741\,
            I => \N__28727\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__28736\,
            I => \N__28724\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__28731\,
            I => \N__28721\
        );

    \I__4877\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28716\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28716\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__28724\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__28721\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__28716\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28705\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28702\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28699\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28696\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__28699\,
            I => \N__28692\
        );

    \I__4867\ : Span12Mux_h
    port map (
            O => \N__28696\,
            I => \N__28689\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28686\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__28692\,
            I => \N__28683\
        );

    \I__4864\ : Odrv12
    port map (
            O => \N__28689\,
            I => \pid_side.error_p_regZ0Z_12\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__28686\,
            I => \pid_side.error_p_regZ0Z_12\
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__28683\,
            I => \pid_side.error_p_regZ0Z_12\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__28673\,
            I => \pid_side.un1_pid_prereg_cry_11_THRU_CO\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28667\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28667\,
            I => \pid_side.un1_pid_prereg_cry_17_THRU_CO\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__4856\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28658\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28654\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28651\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__28654\,
            I => \N__28646\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28646\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__28646\,
            I => \N__28642\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28639\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__28642\,
            I => \N__28636\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28639\,
            I => \pid_side.error_p_regZ0Z_18\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__28636\,
            I => \pid_side.error_p_regZ0Z_18\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28628\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__4844\ : Span12Mux_v
    port map (
            O => \N__28625\,
            I => \N__28621\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28618\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__28621\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28618\,
            I => \pid_alt.error_d_reg_prevZ0Z_15\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28609\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__28612\,
            I => \N__28606\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__28609\,
            I => \N__28603\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28600\
        );

    \I__4836\ : Span4Mux_v
    port map (
            O => \N__28603\,
            I => \N__28597\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__28600\,
            I => \N__28594\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__28597\,
            I => \N__28591\
        );

    \I__4833\ : Span12Mux_v
    port map (
            O => \N__28594\,
            I => \N__28588\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__28591\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__4831\ : Odrv12
    port map (
            O => \N__28588\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__28577\,
            I => \N__28573\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28569\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__28573\,
            I => \N__28566\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28563\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__28569\,
            I => \N__28558\
        );

    \I__4823\ : Span4Mux_v
    port map (
            O => \N__28566\,
            I => \N__28558\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28555\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__28558\,
            I => \N__28552\
        );

    \I__4820\ : Span4Mux_v
    port map (
            O => \N__28555\,
            I => \N__28549\
        );

    \I__4819\ : Span4Mux_h
    port map (
            O => \N__28552\,
            I => \N__28546\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__28549\,
            I => \N__28543\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__28546\,
            I => \pid_alt.error_d_regZ0Z_15\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__28543\,
            I => \pid_alt.error_d_regZ0Z_15\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28532\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28532\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4811\ : Span4Mux_h
    port map (
            O => \N__28526\,
            I => \N__28523\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__28523\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28520\,
            I => \N__28517\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__28508\,
            I => \pid_side.error_axb_8_l_ofxZ0\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28496\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28496\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28496\,
            I => side_command_7
        );

    \I__4800\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28490\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28490\,
            I => \N__28487\
        );

    \I__4798\ : Span4Mux_h
    port map (
            O => \N__28487\,
            I => \N__28484\
        );

    \I__4797\ : Span4Mux_h
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__28481\,
            I => \pid_side.error_axbZ0Z_7\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__28475\,
            I => \drone_H_disp_front_2\
        );

    \I__4793\ : InMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28469\,
            I => \drone_H_disp_side_1\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28463\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28463\,
            I => \N__28460\
        );

    \I__4789\ : Odrv12
    port map (
            O => \N__28460\,
            I => \pid_side.error_axbZ0Z_1\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28454\,
            I => \pid_side.un1_pid_prereg_cry_7_THRU_CO\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28447\
        );

    \I__4785\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28444\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28439\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28444\,
            I => \N__28439\
        );

    \I__4782\ : Span4Mux_v
    port map (
            O => \N__28439\,
            I => \N__28435\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28432\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__28435\,
            I => \N__28429\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28432\,
            I => \pid_side.error_p_regZ0Z_8\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__28429\,
            I => \pid_side.error_p_regZ0Z_8\
        );

    \I__4777\ : InMux
    port map (
            O => \N__28424\,
            I => \N__28421\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__28421\,
            I => \N__28417\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28414\
        );

    \I__4774\ : Span4Mux_v
    port map (
            O => \N__28417\,
            I => \N__28409\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28414\,
            I => \N__28409\
        );

    \I__4772\ : Span4Mux_h
    port map (
            O => \N__28409\,
            I => \N__28405\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__4770\ : Span4Mux_h
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__28402\,
            I => \pid_side.error_p_regZ0Z_11\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__28399\,
            I => \pid_side.error_p_regZ0Z_11\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28391\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28391\,
            I => \pid_side.un1_pid_prereg_cry_10_THRU_CO\
        );

    \I__4765\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28385\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28385\,
            I => \pid_side.un1_pid_prereg_cry_3_THRU_CO\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28378\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28375\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28372\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28369\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__28372\,
            I => \N__28363\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__28369\,
            I => \N__28363\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28360\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28360\,
            I => \pid_side.error_p_regZ0Z_4\
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__28357\,
            I => \pid_side.error_p_regZ0Z_4\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28349\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28349\,
            I => \N__28345\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28342\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__28345\,
            I => \N__28337\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28342\,
            I => \N__28337\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__28337\,
            I => \N__28333\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28330\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__28333\,
            I => \N__28327\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28330\,
            I => \pid_side.error_p_regZ0Z_6\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__28327\,
            I => \pid_side.error_p_regZ0Z_6\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__28319\,
            I => \pid_side.un1_pid_prereg_cry_5_THRU_CO\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28313\,
            I => \pid_side.un1_pid_prereg_cry_18_THRU_CO\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__28310\,
            I => \N__28307\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28303\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28300\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28303\,
            I => \N__28297\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__28300\,
            I => \N__28294\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__28297\,
            I => \N__28290\
        );

    \I__4733\ : Span4Mux_v
    port map (
            O => \N__28294\,
            I => \N__28287\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28284\
        );

    \I__4731\ : Sp12to4
    port map (
            O => \N__28290\,
            I => \N__28279\
        );

    \I__4730\ : Sp12to4
    port map (
            O => \N__28287\,
            I => \N__28279\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__28284\,
            I => \pid_side.error_p_regZ0Z_19\
        );

    \I__4728\ : Odrv12
    port map (
            O => \N__28279\,
            I => \pid_side.error_p_regZ0Z_19\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__28271\,
            I => \N__28268\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__28268\,
            I => \N__28264\
        );

    \I__4724\ : InMux
    port map (
            O => \N__28267\,
            I => \N__28261\
        );

    \I__4723\ : Sp12to4
    port map (
            O => \N__28264\,
            I => \N__28255\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28255\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28252\
        );

    \I__4720\ : Span12Mux_v
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__28252\,
            I => \pid_side.error_p_regZ0Z_15\
        );

    \I__4718\ : Odrv12
    port map (
            O => \N__28249\,
            I => \pid_side.error_p_regZ0Z_15\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__28241\,
            I => \pid_side.un1_pid_prereg_cry_14_THRU_CO\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28235\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28231\
        );

    \I__4713\ : InMux
    port map (
            O => \N__28234\,
            I => \N__28228\
        );

    \I__4712\ : Span4Mux_h
    port map (
            O => \N__28231\,
            I => \N__28223\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__28228\,
            I => \N__28223\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__4709\ : Span4Mux_h
    port map (
            O => \N__28220\,
            I => \N__28216\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28213\
        );

    \I__4707\ : Span4Mux_s1_h
    port map (
            O => \N__28216\,
            I => \N__28210\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__28213\,
            I => \pid_side.error_p_regZ0Z_14\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__28210\,
            I => \pid_side.error_p_regZ0Z_14\
        );

    \I__4704\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__28202\,
            I => \pid_side.un1_pid_prereg_cry_13_THRU_CO\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28196\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__28196\,
            I => \pid_side.un1_pid_prereg_cry_16_THRU_CO\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28186\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28183\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__28186\,
            I => \N__28180\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__28183\,
            I => \N__28177\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__28180\,
            I => \N__28173\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__28177\,
            I => \N__28170\
        );

    \I__4693\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28167\
        );

    \I__4692\ : Span4Mux_h
    port map (
            O => \N__28173\,
            I => \N__28164\
        );

    \I__4691\ : Span4Mux_h
    port map (
            O => \N__28170\,
            I => \N__28161\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__28167\,
            I => \pid_side.error_p_regZ0Z_17\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__28164\,
            I => \pid_side.error_p_regZ0Z_17\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__28161\,
            I => \pid_side.error_p_regZ0Z_17\
        );

    \I__4687\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__28151\,
            I => \pid_side.un1_pid_prereg_cry_19_THRU_CO\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28143\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28138\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28138\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__28143\,
            I => \N__28132\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28132\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28129\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28129\,
            I => \pid_side.error_p_regZ0Z_20\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__28126\,
            I => \pid_side.error_p_regZ0Z_20\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__28121\,
            I => \N__28115\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28109\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28109\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28102\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28102\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28102\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__28109\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__28102\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__28088\,
            I => \N__28085\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__28085\,
            I => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__28082\,
            I => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__28079\,
            I => \N__28074\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__28078\,
            I => \N__28071\
        );

    \I__4660\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28066\
        );

    \I__4659\ : InMux
    port map (
            O => \N__28074\,
            I => \N__28066\
        );

    \I__4658\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28063\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__28066\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__28063\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28055\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28055\,
            I => \N__28047\
        );

    \I__4653\ : InMux
    port map (
            O => \N__28054\,
            I => \N__28042\
        );

    \I__4652\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28042\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28037\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28037\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28034\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__28047\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28042\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__28037\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28034\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__4644\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28022\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__28019\,
            I => \dron_frame_decoder_1.N_412_4\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__4640\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__28010\,
            I => \dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0\
        );

    \I__4638\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__28004\,
            I => \dron_frame_decoder_1.N_175\
        );

    \I__4636\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27995\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27990\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27990\
        );

    \I__4633\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27987\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__27995\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__27990\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27987\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__27977\,
            I => \N__27973\
        );

    \I__4627\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27970\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__27973\,
            I => \dron_frame_decoder_1.N_431\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__27970\,
            I => \dron_frame_decoder_1.N_431\
        );

    \I__4624\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27960\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27957\
        );

    \I__4622\ : InMux
    port map (
            O => \N__27963\,
            I => \N__27954\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__27960\,
            I => \dron_frame_decoder_1.N_435\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__27957\,
            I => \dron_frame_decoder_1.N_435\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__27954\,
            I => \dron_frame_decoder_1.N_435\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__27947\,
            I => \N__27943\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__27946\,
            I => \N__27939\
        );

    \I__4616\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27936\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27933\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27930\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__27936\,
            I => \N__27925\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27925\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27930\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__27925\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__4609\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27917\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__27917\,
            I => \N__27914\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__27914\,
            I => \N__27911\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__27911\,
            I => \pid_side.un1_pid_prereg_cry_8_THRU_CO\
        );

    \I__4605\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27904\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__27907\,
            I => \N__27901\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27898\
        );

    \I__4602\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27895\
        );

    \I__4601\ : Span4Mux_h
    port map (
            O => \N__27898\,
            I => \N__27889\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__27895\,
            I => \N__27889\
        );

    \I__4599\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27886\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27878\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__27883\,
            I => \N__27878\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__27878\,
            I => \pid_side.error_p_regZ0Z_9\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27863\
        );

    \I__4593\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27863\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27863\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27856\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27856\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27856\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__27863\,
            I => \N__27849\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27856\,
            I => \N__27849\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27855\,
            I => \N__27844\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27844\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__27849\,
            I => \dron_frame_decoder_1.N_428\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__27844\,
            I => \dron_frame_decoder_1.N_428\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27831\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27828\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__27834\,
            I => \N__27825\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27822\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27819\
        );

    \I__4576\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27816\
        );

    \I__4575\ : Span4Mux_v
    port map (
            O => \N__27822\,
            I => \N__27813\
        );

    \I__4574\ : Odrv12
    port map (
            O => \N__27819\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27816\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__4572\ : Odrv4
    port map (
            O => \N__27813\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__4571\ : CascadeMux
    port map (
            O => \N__27806\,
            I => \dron_frame_decoder_1.N_412_4_cascade_\
        );

    \I__4570\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27798\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27795\
        );

    \I__4568\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27792\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__27798\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__27795\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__27792\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__27785\,
            I => \N__27781\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27777\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27774\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27771\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__27777\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__27774\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__27771\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27758\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__27758\,
            I => \dron_frame_decoder_1.WDT10lt14_0\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__27755\,
            I => \dron_frame_decoder_1.N_177_cascade_\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27746\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27743\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27740\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27737\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__27746\,
            I => \N__27734\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27743\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27740\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__27737\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__27734\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27722\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__27722\,
            I => \dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27710\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27710\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27710\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27707\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27695\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27695\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27695\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27692\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27686\,
            I => \N__27680\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27680\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__27680\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27677\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__27674\,
            I => \N__27671\
        );

    \I__4526\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27665\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27665\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27665\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27662\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27650\
        );

    \I__4520\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27650\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27650\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27647\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__4517\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27640\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__27640\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27637\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__27632\,
            I => \N__27629\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27626\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27623\,
            I => \bfn_9_11_0_\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27620\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__27617\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27594\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27591\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27588\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27585\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27582\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27579\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__27608\,
            I => \N__27574\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27569\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27569\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27564\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27551\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27551\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27551\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27551\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27551\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27551\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27546\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27546\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27541\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27591\,
            I => \N__27541\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27538\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__27585\,
            I => \N__27530\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__27582\,
            I => \N__27530\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27579\,
            I => \N__27527\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27578\,
            I => \N__27524\
        );

    \I__4482\ : InMux
    port map (
            O => \N__27577\,
            I => \N__27519\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27519\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27516\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27511\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27511\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27508\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27551\,
            I => \N__27505\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27498\
        );

    \I__4474\ : Span4Mux_h
    port map (
            O => \N__27541\,
            I => \N__27498\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__27538\,
            I => \N__27498\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27495\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27492\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27488\
        );

    \I__4469\ : Span12Mux_v
    port map (
            O => \N__27530\,
            I => \N__27485\
        );

    \I__4468\ : Span4Mux_h
    port map (
            O => \N__27527\,
            I => \N__27478\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27524\,
            I => \N__27478\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__27519\,
            I => \N__27478\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__27516\,
            I => \N__27471\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27471\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__27508\,
            I => \N__27471\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__27505\,
            I => \N__27468\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__27498\,
            I => \N__27461\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27461\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__27492\,
            I => \N__27461\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27458\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27488\,
            I => uart_pc_data_rdy
        );

    \I__4456\ : Odrv12
    port map (
            O => \N__27485\,
            I => uart_pc_data_rdy
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__27478\,
            I => uart_pc_data_rdy
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27471\,
            I => uart_pc_data_rdy
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__27468\,
            I => uart_pc_data_rdy
        );

    \I__4452\ : Odrv4
    port map (
            O => \N__27461\,
            I => uart_pc_data_rdy
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__27458\,
            I => uart_pc_data_rdy
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__27443\,
            I => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27435\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27430\
        );

    \I__4447\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27430\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27425\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27425\
        );

    \I__4444\ : Odrv12
    port map (
            O => \N__27425\,
            I => \Commands_frame_decoder.N_422\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27416\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27413\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27420\,
            I => \N__27410\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27407\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27403\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__27413\,
            I => \N__27400\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27397\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27394\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27391\
        );

    \I__4434\ : Span12Mux_v
    port map (
            O => \N__27403\,
            I => \N__27386\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__27400\,
            I => \N__27383\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__27397\,
            I => \N__27376\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__27394\,
            I => \N__27376\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27376\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27371\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27371\
        );

    \I__4427\ : Odrv12
    port map (
            O => \N__27386\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__27383\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__27376\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27371\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__27362\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__27359\,
            I => \N__27355\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27352\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27349\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27352\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27349\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27338\,
            I => \N__27335\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__27335\,
            I => \N__27331\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27328\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__27331\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27328\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27317\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__27317\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27314\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__27311\,
            I => \N__27308\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__4404\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27302\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__27302\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27299\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__27293\,
            I => uart_input_pc_c
        );

    \I__4399\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27287\,
            I => \uart_pc_sync.aux_0__0_Z0Z_0\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__27281\,
            I => \uart_pc_sync.aux_1__0_Z0Z_0\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27275\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27275\,
            I => \uart_pc_sync.aux_2__0_Z0Z_0\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__27269\,
            I => \uart_pc_sync.aux_3__0_Z0Z_0\
        );

    \I__4391\ : InMux
    port map (
            O => \N__27266\,
            I => \N__27262\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27265\,
            I => \N__27259\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27262\,
            I => \N__27256\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__27259\,
            I => \N__27251\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__27256\,
            I => \N__27248\
        );

    \I__4386\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27245\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27242\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__27251\,
            I => \N__27239\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__27248\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27245\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27242\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__27239\,
            I => \Commands_frame_decoder.stateZ0Z_14\
        );

    \I__4379\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27226\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__27229\,
            I => \N__27223\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__27226\,
            I => \N__27220\
        );

    \I__4376\ : InMux
    port map (
            O => \N__27223\,
            I => \N__27216\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__27220\,
            I => \N__27213\
        );

    \I__4374\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27210\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__27216\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__27213\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__27210\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__4370\ : IoInMux
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__27200\,
            I => \N__27197\
        );

    \I__4368\ : Span4Mux_s1_v
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__27194\,
            I => \N__27190\
        );

    \I__4366\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27187\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__27190\,
            I => \N__27183\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27187\,
            I => \N__27180\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__27186\,
            I => \N__27177\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__27183\,
            I => \N__27171\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__27180\,
            I => \N__27171\
        );

    \I__4360\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27168\
        );

    \I__4359\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27165\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__27171\,
            I => \debug_CH3_20A_c\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27168\,
            I => \debug_CH3_20A_c\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__27165\,
            I => \debug_CH3_20A_c\
        );

    \I__4355\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27155\,
            I => \N__27151\
        );

    \I__4353\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27148\
        );

    \I__4352\ : Span12Mux_s8_h
    port map (
            O => \N__27151\,
            I => \N__27145\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27142\
        );

    \I__4350\ : Odrv12
    port map (
            O => \N__27145\,
            I => \drone_H_disp_side_0\
        );

    \I__4349\ : Odrv12
    port map (
            O => \N__27142\,
            I => \drone_H_disp_side_0\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__27134\,
            I => \drone_H_disp_side_2\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27128\,
            I => \drone_H_disp_side_3\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__27122\,
            I => \dron_frame_decoder_1.drone_H_disp_side_4\
        );

    \I__4342\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27116\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__27116\,
            I => \dron_frame_decoder_1.drone_H_disp_side_5\
        );

    \I__4340\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__27107\,
            I => \dron_frame_decoder_1.drone_H_disp_side_6\
        );

    \I__4337\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27101\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__27101\,
            I => \dron_frame_decoder_1.drone_H_disp_side_7\
        );

    \I__4335\ : CEMux
    port map (
            O => \N__27098\,
            I => \N__27095\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__27095\,
            I => \N__27092\
        );

    \I__4333\ : Odrv12
    port map (
            O => \N__27092\,
            I => \dron_frame_decoder_1.N_747_0\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27086\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27086\,
            I => \N__27083\
        );

    \I__4330\ : Span4Mux_s1_h
    port map (
            O => \N__27083\,
            I => \N__27080\
        );

    \I__4329\ : Sp12to4
    port map (
            O => \N__27080\,
            I => \N__27077\
        );

    \I__4328\ : Span12Mux_v
    port map (
            O => \N__27077\,
            I => \N__27074\
        );

    \I__4327\ : Odrv12
    port map (
            O => \N__27074\,
            I => alt_ki_7
        );

    \I__4326\ : InMux
    port map (
            O => \N__27071\,
            I => \pid_side.un1_pid_prereg_cry_13\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27068\,
            I => \pid_side.un1_pid_prereg_cry_14\
        );

    \I__4324\ : InMux
    port map (
            O => \N__27065\,
            I => \pid_side.un1_pid_prereg_cry_15\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27062\,
            I => \bfn_8_19_0_\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27059\,
            I => \pid_side.un1_pid_prereg_cry_17\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27056\,
            I => \pid_side.un1_pid_prereg_cry_18\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27053\,
            I => \pid_side.un1_pid_prereg_cry_19\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27050\,
            I => \pid_side.un1_pid_prereg_cry_20\
        );

    \I__4318\ : CEMux
    port map (
            O => \N__27047\,
            I => \N__27044\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__27038\,
            I => \N__27034\
        );

    \I__4314\ : CEMux
    port map (
            O => \N__27037\,
            I => \N__27031\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__27034\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__27031\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27026\,
            I => \pid_side.un1_pid_prereg_cry_4\
        );

    \I__4310\ : InMux
    port map (
            O => \N__27023\,
            I => \pid_side.un1_pid_prereg_cry_5\
        );

    \I__4309\ : InMux
    port map (
            O => \N__27020\,
            I => \pid_side.un1_pid_prereg_cry_6\
        );

    \I__4308\ : InMux
    port map (
            O => \N__27017\,
            I => \pid_side.un1_pid_prereg_cry_7\
        );

    \I__4307\ : InMux
    port map (
            O => \N__27014\,
            I => \bfn_8_18_0_\
        );

    \I__4306\ : InMux
    port map (
            O => \N__27011\,
            I => \pid_side.un1_pid_prereg_cry_9\
        );

    \I__4305\ : InMux
    port map (
            O => \N__27008\,
            I => \pid_side.un1_pid_prereg_cry_10\
        );

    \I__4304\ : InMux
    port map (
            O => \N__27005\,
            I => \pid_side.un1_pid_prereg_cry_11\
        );

    \I__4303\ : InMux
    port map (
            O => \N__27002\,
            I => \pid_side.un1_pid_prereg_cry_12\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__26999\,
            I => \N__26995\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__26998\,
            I => \N__26992\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26987\
        );

    \I__4299\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26980\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26980\
        );

    \I__4297\ : InMux
    port map (
            O => \N__26990\,
            I => \N__26980\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__26987\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__26980\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__26975\,
            I => \N__26971\
        );

    \I__4293\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26966\
        );

    \I__4292\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26966\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__26966\,
            I => \Commands_frame_decoder.stateZ0Z_8\
        );

    \I__4290\ : CEMux
    port map (
            O => \N__26963\,
            I => \N__26960\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__26957\,
            I => \N__26953\
        );

    \I__4287\ : CEMux
    port map (
            O => \N__26956\,
            I => \N__26950\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__26953\,
            I => \N__26947\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26944\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__26947\,
            I => \N__26939\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__26944\,
            I => \N__26939\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__26939\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__4281\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26930\
        );

    \I__4280\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26930\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__26930\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__26924\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__26921\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26904\
        );

    \I__4274\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26904\
        );

    \I__4273\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26904\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26904\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26898\
        );

    \I__4270\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26895\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26890\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26887\
        );

    \I__4267\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26884\
        );

    \I__4266\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26881\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26898\,
            I => \N__26876\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26873\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26868\
        );

    \I__4262\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26868\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__26890\,
            I => \N__26865\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__26887\,
            I => \N__26860\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__26884\,
            I => \N__26860\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26881\,
            I => \N__26857\
        );

    \I__4257\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26852\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26852\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__26876\,
            I => \N__26844\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__26873\,
            I => \N__26844\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26844\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__26865\,
            I => \N__26835\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__26860\,
            I => \N__26835\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__26857\,
            I => \N__26835\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26835\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26832\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__26844\,
            I => \Commands_frame_decoder.N_415\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__26835\,
            I => \Commands_frame_decoder.N_415\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__26832\,
            I => \Commands_frame_decoder.N_415\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__26819\,
            I => \N__26815\
        );

    \I__4241\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26812\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__26815\,
            I => \N__26808\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__26812\,
            I => \N__26805\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26802\
        );

    \I__4237\ : Span4Mux_v
    port map (
            O => \N__26808\,
            I => \N__26799\
        );

    \I__4236\ : Span12Mux_s8_h
    port map (
            O => \N__26805\,
            I => \N__26796\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26802\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__26799\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4233\ : Odrv12
    port map (
            O => \N__26796\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26789\,
            I => \pid_side.un1_pid_prereg_cry_1\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26786\,
            I => \pid_side.un1_pid_prereg_cry_2\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26783\,
            I => \pid_side.un1_pid_prereg_cry_3\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__26771\,
            I => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__26768\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26759\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26759\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__26759\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0\
        );

    \I__4221\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26752\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26749\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__26752\,
            I => \N__26746\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26742\
        );

    \I__4217\ : Span12Mux_s5_h
    port map (
            O => \N__26746\,
            I => \N__26739\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26736\
        );

    \I__4215\ : Span4Mux_s3_h
    port map (
            O => \N__26742\,
            I => \N__26733\
        );

    \I__4214\ : Span12Mux_h
    port map (
            O => \N__26739\,
            I => \N__26730\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26725\
        );

    \I__4212\ : Span4Mux_h
    port map (
            O => \N__26733\,
            I => \N__26725\
        );

    \I__4211\ : Odrv12
    port map (
            O => \N__26730\,
            I => xy_kp_4
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__26725\,
            I => xy_kp_4
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__26720\,
            I => \N__26716\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__26719\,
            I => \N__26713\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26709\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26706\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26703\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26699\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26706\,
            I => \N__26694\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__26703\,
            I => \N__26694\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26702\,
            I => \N__26691\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__26699\,
            I => \N__26688\
        );

    \I__4199\ : Span12Mux_s10_v
    port map (
            O => \N__26694\,
            I => \N__26685\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26691\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__26688\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4196\ : Odrv12
    port map (
            O => \N__26685\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26673\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26668\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26668\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26673\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26668\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26663\,
            I => \dron_frame_decoder_1.un1_WDT_cry_11\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__26660\,
            I => \N__26656\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26656\,
            I => \N__26650\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__26653\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26650\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26645\,
            I => \dron_frame_decoder_1.un1_WDT_cry_12\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26642\,
            I => \dron_frame_decoder_1.un1_WDT_cry_13\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26639\,
            I => \dron_frame_decoder_1.un1_WDT_cry_14\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__26636\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\
        );

    \I__4180\ : SRMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26630\,
            I => \N__26627\
        );

    \I__4178\ : Span4Mux_h
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__26624\,
            I => \N__26620\
        );

    \I__4176\ : SRMux
    port map (
            O => \N__26623\,
            I => \N__26617\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__26620\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__26617\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26609\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26609\,
            I => \dron_frame_decoder_1.WDTZ0Z_3\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26606\,
            I => \dron_frame_decoder_1.un1_WDT_cry_2\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__26603\,
            I => \N__26599\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26593\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26596\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__26593\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26588\,
            I => \dron_frame_decoder_1.un1_WDT_cry_3\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26581\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26578\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26581\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26578\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26573\,
            I => \dron_frame_decoder_1.un1_WDT_cry_4\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26566\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26563\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26566\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26563\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26558\,
            I => \dron_frame_decoder_1.un1_WDT_cry_5\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26551\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26548\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__26551\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26548\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26543\,
            I => \dron_frame_decoder_1.un1_WDT_cry_6\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26536\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26533\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26536\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26533\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26528\,
            I => \bfn_8_12_0_\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26521\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26521\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__26518\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26513\,
            I => \dron_frame_decoder_1.un1_WDT_cry_8\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26506\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26503\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26506\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__26503\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26498\,
            I => \dron_frame_decoder_1.un1_WDT_cry_9\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26490\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26485\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26485\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26490\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26485\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26480\,
            I => \dron_frame_decoder_1.un1_WDT_cry_10\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26474\,
            I => \N__26471\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__26471\,
            I => \scaler_4.N_1684_i_l_ofxZ0\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26468\,
            I => \bfn_8_10_0_\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26465\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__4123\ : SRMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26459\,
            I => \N__26455\
        );

    \I__4121\ : SRMux
    port map (
            O => \N__26458\,
            I => \N__26452\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26446\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__26449\,
            I => \N__26441\
        );

    \I__4117\ : Span4Mux_h
    port map (
            O => \N__26446\,
            I => \N__26441\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__26441\,
            I => \Commands_frame_decoder.un1_state57_iZ0\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__26438\,
            I => \N__26434\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26431\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26428\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26431\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26428\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__26420\,
            I => \dron_frame_decoder_1.WDTZ0Z_0\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26414\,
            I => \dron_frame_decoder_1.WDTZ0Z_1\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26411\,
            I => \dron_frame_decoder_1.un1_WDT_cry_0\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26405\,
            I => \dron_frame_decoder_1.WDTZ0Z_2\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26402\,
            I => \dron_frame_decoder_1.un1_WDT_cry_1\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26396\,
            I => \frame_decoder_CH4data_1\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26387\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26384\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26378\,
            I => \frame_decoder_CH4data_2\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__26369\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26366\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__26360\,
            I => \frame_decoder_CH4data_3\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__26351\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26348\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26342\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26342\,
            I => \frame_decoder_CH4data_4\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__4081\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__26333\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26330\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__26318\,
            I => \frame_decoder_CH4data_5\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__4073\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26309\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__4071\ : InMux
    port map (
            O => \N__26306\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__4070\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26300\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26300\,
            I => \frame_decoder_CH4data_6\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__4064\ : Span4Mux_h
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__26282\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__4062\ : InMux
    port map (
            O => \N__26279\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__4061\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__4059\ : Span12Mux_s9_v
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__4058\ : Odrv12
    port map (
            O => \N__26267\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26264\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26257\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26254\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__26257\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26254\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26249\,
            I => \Commands_frame_decoder.un1_WDT_cry_6\
        );

    \I__4051\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26242\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26239\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__26242\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26239\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26234\,
            I => \bfn_8_8_0_\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__26231\,
            I => \N__26227\
        );

    \I__4045\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26224\
        );

    \I__4044\ : InMux
    port map (
            O => \N__26227\,
            I => \N__26221\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26224\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__26221\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26216\,
            I => \Commands_frame_decoder.un1_WDT_cry_8\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26209\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26206\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__26209\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26206\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__4036\ : InMux
    port map (
            O => \N__26201\,
            I => \Commands_frame_decoder.un1_WDT_cry_9\
        );

    \I__4035\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26193\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26188\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26188\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26193\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26188\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26183\,
            I => \Commands_frame_decoder.un1_WDT_cry_10\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26175\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26170\
        );

    \I__4027\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26170\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26175\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__26170\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26165\,
            I => \Commands_frame_decoder.un1_WDT_cry_11\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__26162\,
            I => \N__26158\
        );

    \I__4022\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26155\
        );

    \I__4021\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26152\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__26155\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__26152\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__4018\ : InMux
    port map (
            O => \N__26147\,
            I => \Commands_frame_decoder.un1_WDT_cry_12\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26131\
        );

    \I__4015\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26131\
        );

    \I__4014\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26131\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__26138\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__26131\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26126\,
            I => \Commands_frame_decoder.un1_WDT_cry_13\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26123\,
            I => \Commands_frame_decoder.un1_WDT_cry_14\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__26120\,
            I => \N__26117\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26109\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26116\,
            I => \N__26109\
        );

    \I__4006\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26106\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26103\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26109\,
            I => \N__26100\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26106\,
            I => \N__26097\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__26103\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__26100\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__26097\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__26087\,
            I => \Commands_frame_decoder.count_1_sqmuxa\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__26084\,
            I => \N__26080\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26083\,
            I => \N__26077\
        );

    \I__3995\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26074\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26077\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__26074\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26066\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__26066\,
            I => \Commands_frame_decoder.WDTZ0Z_0\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__26060\,
            I => \Commands_frame_decoder.WDTZ0Z_1\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26057\,
            I => \Commands_frame_decoder.un1_WDT_cry_0\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26051\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__26051\,
            I => \Commands_frame_decoder.WDTZ0Z_2\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26048\,
            I => \Commands_frame_decoder.un1_WDT_cry_1\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26042\,
            I => \Commands_frame_decoder.WDTZ0Z_3\
        );

    \I__3982\ : InMux
    port map (
            O => \N__26039\,
            I => \Commands_frame_decoder.un1_WDT_cry_2\
        );

    \I__3981\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26032\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26029\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26032\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__26029\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26024\,
            I => \Commands_frame_decoder.un1_WDT_cry_3\
        );

    \I__3976\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26017\
        );

    \I__3975\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26014\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__26017\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__26014\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26009\,
            I => \Commands_frame_decoder.un1_WDT_cry_4\
        );

    \I__3971\ : InMux
    port map (
            O => \N__26006\,
            I => \N__26002\
        );

    \I__3970\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25999\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__26002\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__25999\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25994\,
            I => \Commands_frame_decoder.un1_WDT_cry_5\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__25985\,
            I => \pid_side.error_axbZ0Z_2\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__25976\,
            I => \pid_side.error_axbZ0Z_3\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25970\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__3958\ : Span4Mux_s3_h
    port map (
            O => \N__25967\,
            I => \N__25963\
        );

    \I__3957\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25960\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__25963\,
            I => \N__25957\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25960\,
            I => alt_kp_4
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__25957\,
            I => alt_kp_4
        );

    \I__3953\ : CEMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25944\
        );

    \I__3951\ : CEMux
    port map (
            O => \N__25948\,
            I => \N__25941\
        );

    \I__3950\ : CEMux
    port map (
            O => \N__25947\,
            I => \N__25938\
        );

    \I__3949\ : Span4Mux_s3_h
    port map (
            O => \N__25944\,
            I => \N__25933\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25941\,
            I => \N__25933\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__25938\,
            I => \N__25930\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__25933\,
            I => \N__25925\
        );

    \I__3945\ : Span4Mux_h
    port map (
            O => \N__25930\,
            I => \N__25925\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__25925\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25916\
        );

    \I__3941\ : Span12Mux_s8_v
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__3940\ : Odrv12
    port map (
            O => \N__25913\,
            I => \pid_alt.state_RNIFCSD1Z0Z_0\
        );

    \I__3939\ : IoInMux
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__3937\ : Span4Mux_s1_v
    port map (
            O => \N__25904\,
            I => \N__25901\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__25901\,
            I => \pid_alt.N_850_0\
        );

    \I__3935\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__25895\,
            I => uart_input_drone_c
        );

    \I__3933\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25889\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__25889\,
            I => \uart_drone_sync.aux_0__0__0_0\
        );

    \I__3931\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25883\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25883\,
            I => \uart_drone_sync.aux_1__0__0_0\
        );

    \I__3929\ : CEMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__3926\ : Span4Mux_h
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__25868\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__25859\,
            I => \N__25856\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__25856\,
            I => \pid_alt.pid_preregZ0Z_14\
        );

    \I__3920\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25850\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__25847\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__25835\,
            I => \pid_alt.pid_preregZ0Z_16\
        );

    \I__3913\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__25826\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_5\
        );

    \I__3910\ : CEMux
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__25820\,
            I => \N__25816\
        );

    \I__3908\ : CEMux
    port map (
            O => \N__25819\,
            I => \N__25813\
        );

    \I__3907\ : Span4Mux_s3_h
    port map (
            O => \N__25816\,
            I => \N__25810\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__25813\,
            I => \N__25807\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__25810\,
            I => \N__25804\
        );

    \I__3904\ : Span4Mux_v
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__25804\,
            I => \dron_frame_decoder_1.N_755_0\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__25801\,
            I => \dron_frame_decoder_1.N_755_0\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25793\,
            I => \N__25790\
        );

    \I__3899\ : Odrv12
    port map (
            O => \N__25790\,
            I => \dron_frame_decoder_1.drone_altitude_7\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25783\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25780\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25783\,
            I => \N__25777\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25780\,
            I => \N__25774\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__25774\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__25771\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__25757\,
            I => \drone_H_disp_side_i_4\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__25745\,
            I => \drone_H_disp_side_i_7\
        );

    \I__3883\ : CascadeMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__3882\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25733\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__25733\,
            I => \drone_H_disp_side_i_5\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25727\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__25724\,
            I => \pid_alt.m7_e_4\
        );

    \I__3876\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25718\,
            I => \N__25715\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__25715\,
            I => \N__25710\
        );

    \I__3873\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25705\
        );

    \I__3872\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25705\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25710\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__25705\,
            I => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__25694\,
            I => \pid_alt.error_i_acumm_preregZ0Z_19\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__25691\,
            I => \pid_alt.un1_reset_i_a5_1_10_7_cascade_\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25680\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25675\
        );

    \I__3862\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25675\
        );

    \I__3861\ : Odrv12
    port map (
            O => \N__25680\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__25675\,
            I => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25667\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__25667\,
            I => \pid_alt.error_i_acumm_preregZ0Z_18\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25661\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25661\,
            I => \N__25656\
        );

    \I__3855\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25651\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25651\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__25656\,
            I => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__25651\,
            I => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25643\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25643\,
            I => \pid_alt.error_i_acumm_preregZ0Z_17\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25637\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25632\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25627\
        );

    \I__3846\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25627\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__25632\,
            I => \N__25622\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__25627\,
            I => \N__25622\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__25619\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25613\,
            I => \N__25610\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__25607\,
            I => \N__25604\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__25604\,
            I => \pid_alt.error_i_acumm_preregZ0Z_20\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25598\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25598\,
            I => \N__25593\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25588\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25588\
        );

    \I__3832\ : Odrv12
    port map (
            O => \N__25593\,
            I => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25588\,
            I => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25580\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25580\,
            I => \pid_alt.error_i_acumm_preregZ0Z_16\
        );

    \I__3828\ : CEMux
    port map (
            O => \N__25577\,
            I => \N__25505\
        );

    \I__3827\ : CEMux
    port map (
            O => \N__25576\,
            I => \N__25505\
        );

    \I__3826\ : CEMux
    port map (
            O => \N__25575\,
            I => \N__25505\
        );

    \I__3825\ : CEMux
    port map (
            O => \N__25574\,
            I => \N__25505\
        );

    \I__3824\ : CEMux
    port map (
            O => \N__25573\,
            I => \N__25505\
        );

    \I__3823\ : CEMux
    port map (
            O => \N__25572\,
            I => \N__25505\
        );

    \I__3822\ : CEMux
    port map (
            O => \N__25571\,
            I => \N__25505\
        );

    \I__3821\ : CEMux
    port map (
            O => \N__25570\,
            I => \N__25505\
        );

    \I__3820\ : CEMux
    port map (
            O => \N__25569\,
            I => \N__25505\
        );

    \I__3819\ : CEMux
    port map (
            O => \N__25568\,
            I => \N__25505\
        );

    \I__3818\ : CEMux
    port map (
            O => \N__25567\,
            I => \N__25505\
        );

    \I__3817\ : CEMux
    port map (
            O => \N__25566\,
            I => \N__25505\
        );

    \I__3816\ : CEMux
    port map (
            O => \N__25565\,
            I => \N__25505\
        );

    \I__3815\ : CEMux
    port map (
            O => \N__25564\,
            I => \N__25505\
        );

    \I__3814\ : CEMux
    port map (
            O => \N__25563\,
            I => \N__25505\
        );

    \I__3813\ : CEMux
    port map (
            O => \N__25562\,
            I => \N__25505\
        );

    \I__3812\ : CEMux
    port map (
            O => \N__25561\,
            I => \N__25505\
        );

    \I__3811\ : CEMux
    port map (
            O => \N__25560\,
            I => \N__25505\
        );

    \I__3810\ : CEMux
    port map (
            O => \N__25559\,
            I => \N__25505\
        );

    \I__3809\ : CEMux
    port map (
            O => \N__25558\,
            I => \N__25505\
        );

    \I__3808\ : CEMux
    port map (
            O => \N__25557\,
            I => \N__25505\
        );

    \I__3807\ : CEMux
    port map (
            O => \N__25556\,
            I => \N__25505\
        );

    \I__3806\ : CEMux
    port map (
            O => \N__25555\,
            I => \N__25505\
        );

    \I__3805\ : CEMux
    port map (
            O => \N__25554\,
            I => \N__25505\
        );

    \I__3804\ : GlobalMux
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__3803\ : gio2CtrlBuf
    port map (
            O => \N__25502\,
            I => \pid_alt.state_0_g_0\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25487\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25498\,
            I => \N__25487\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25487\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25487\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25483\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25480\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__25483\,
            I => \N__25477\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25474\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__25477\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__25474\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25463\,
            I => \dron_frame_decoder_1.WDT10lto13_1\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__25460\,
            I => \dron_frame_decoder_1.WDT10lt14_0_cascade_\
        );

    \I__3788\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25454\,
            I => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\
        );

    \I__3786\ : InMux
    port map (
            O => \N__25451\,
            I => \N__25447\
        );

    \I__3785\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25444\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25441\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__25444\,
            I => \N__25438\
        );

    \I__3782\ : Odrv12
    port map (
            O => \N__25441\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__25438\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25430\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25430\,
            I => \N__25426\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__25426\,
            I => \N__25420\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25417\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__25420\,
            I => \N__25414\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__25417\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__25414\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__25409\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25402\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25399\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25402\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25399\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25390\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25387\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25382\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25387\,
            I => \N__25382\
        );

    \I__3763\ : Odrv12
    port map (
            O => \N__25382\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__25373\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25364\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25364\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__25364\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__3756\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25355\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25355\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25355\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__25346\,
            I => \Commands_frame_decoder.N_377_0\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__25343\,
            I => \Commands_frame_decoder.N_377_0_cascade_\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__25337\,
            I => \N__25333\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25330\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__25333\,
            I => \Commands_frame_decoder.N_384\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25330\,
            I => \Commands_frame_decoder.N_384\
        );

    \I__3744\ : CEMux
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3742\ : Span4Mux_v
    port map (
            O => \N__25319\,
            I => \N__25315\
        );

    \I__3741\ : CEMux
    port map (
            O => \N__25318\,
            I => \N__25312\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__25315\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25312\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__25307\,
            I => \N__25303\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__25306\,
            I => \N__25300\
        );

    \I__3736\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25297\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25294\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__25297\,
            I => \N__25291\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25294\,
            I => \Commands_frame_decoder.stateZ0Z_12\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__25291\,
            I => \Commands_frame_decoder.stateZ0Z_12\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25280\
        );

    \I__3730\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25280\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__25280\,
            I => \Commands_frame_decoder.stateZ0Z_13\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25274\,
            I => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \Commands_frame_decoder.WDT8lto13_1_cascade_\
        );

    \I__3725\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__25265\,
            I => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25258\
        );

    \I__3722\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25255\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25258\,
            I => \N__25252\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25248\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__25252\,
            I => \N__25245\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25242\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__25248\,
            I => \N__25239\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__25245\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__25242\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__25239\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__25232\,
            I => \Commands_frame_decoder.WDT8lt14_0_cascade_\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__25226\,
            I => \drone_H_disp_side_i_6\
        );

    \I__3710\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__25217\,
            I => side_command_0
        );

    \I__3707\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25211\,
            I => side_command_1
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25202\,
            I => side_command_2
        );

    \I__3702\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__25196\,
            I => side_command_3
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25187\,
            I => side_command_4
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25178\,
            I => side_command_5
        );

    \I__3694\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25172\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__25172\,
            I => side_command_6
        );

    \I__3692\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25163\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__25163\,
            I => \drone_H_disp_side_15\
        );

    \I__3689\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__25154\,
            I => \dron_frame_decoder_1.drone_altitude_5\
        );

    \I__3686\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25148\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__25145\,
            I => \dron_frame_decoder_1.drone_altitude_6\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25138\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25135\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__25138\,
            I => \N__25132\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__3679\ : Span12Mux_s10_v
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__3678\ : Span4Mux_s3_h
    port map (
            O => \N__25129\,
            I => \N__25123\
        );

    \I__3677\ : Span12Mux_h
    port map (
            O => \N__25126\,
            I => \N__25120\
        );

    \I__3676\ : Span4Mux_v
    port map (
            O => \N__25123\,
            I => \N__25117\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__25120\,
            I => xy_kp_0
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__25117\,
            I => xy_kp_0
        );

    \I__3673\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__3671\ : Span4Mux_s1_h
    port map (
            O => \N__25106\,
            I => \N__25102\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25099\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__25102\,
            I => \N__25096\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25093\
        );

    \I__3667\ : Sp12to4
    port map (
            O => \N__25096\,
            I => \N__25090\
        );

    \I__3666\ : Span4Mux_s2_h
    port map (
            O => \N__25093\,
            I => \N__25087\
        );

    \I__3665\ : Span12Mux_h
    port map (
            O => \N__25090\,
            I => \N__25084\
        );

    \I__3664\ : Span4Mux_h
    port map (
            O => \N__25087\,
            I => \N__25081\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__25084\,
            I => xy_kp_2
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__25081\,
            I => xy_kp_2
        );

    \I__3661\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3659\ : Span4Mux_s3_h
    port map (
            O => \N__25070\,
            I => \N__25066\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25063\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__25063\,
            I => \N__25057\
        );

    \I__3655\ : Span4Mux_v
    port map (
            O => \N__25060\,
            I => \N__25054\
        );

    \I__3654\ : Span4Mux_s2_h
    port map (
            O => \N__25057\,
            I => \N__25051\
        );

    \I__3653\ : Sp12to4
    port map (
            O => \N__25054\,
            I => \N__25048\
        );

    \I__3652\ : Span4Mux_v
    port map (
            O => \N__25051\,
            I => \N__25045\
        );

    \I__3651\ : Odrv12
    port map (
            O => \N__25048\,
            I => xy_kp_6
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__25045\,
            I => xy_kp_6
        );

    \I__3649\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25037\,
            I => \dron_frame_decoder_1.drone_altitude_4\
        );

    \I__3647\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__25025\,
            I => drone_altitude_i_4
        );

    \I__3643\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25019\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__25016\,
            I => \N__25012\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__3639\ : Span4Mux_v
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__3638\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__25006\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25003\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__3635\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24995\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__24989\,
            I => \N__24985\
        );

    \I__3631\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24982\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__24985\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__24982\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__3628\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__24974\,
            I => \N__24970\
        );

    \I__3626\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24967\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__24970\,
            I => \N__24964\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24967\,
            I => \N__24961\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__24964\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__3622\ : Odrv12
    port map (
            O => \N__24961\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__3621\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__24953\,
            I => \drone_H_disp_side_i_13\
        );

    \I__3619\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24946\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \N__24943\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24940\
        );

    \I__3616\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24937\
        );

    \I__3615\ : Span4Mux_v
    port map (
            O => \N__24940\,
            I => \N__24932\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__24937\,
            I => \N__24932\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__24932\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__24929\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\
        );

    \I__3611\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24923\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__24923\,
            I => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\
        );

    \I__3609\ : InMux
    port map (
            O => \N__24920\,
            I => \N__24914\
        );

    \I__3608\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24914\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__24914\,
            I => \N__24911\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__24911\,
            I => \N__24907\
        );

    \I__3605\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__24907\,
            I => \N__24899\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24899\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__24896\,
            I => \N__24893\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__24893\,
            I => \pid_alt.error_d_regZ0Z_19\
        );

    \I__3599\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24887\,
            I => \N__24883\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24880\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__24883\,
            I => \N__24877\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24880\,
            I => \pid_alt.error_d_reg_prevZ0Z_19\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__24877\,
            I => \pid_alt.error_d_reg_prevZ0Z_19\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24866\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24866\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__24866\,
            I => \pid_alt.error_d_reg_prevZ0Z_20\
        );

    \I__3590\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24857\
        );

    \I__3589\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24857\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__3587\ : Span4Mux_h
    port map (
            O => \N__24854\,
            I => \N__24851\
        );

    \I__3586\ : Span4Mux_v
    port map (
            O => \N__24851\,
            I => \N__24848\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__24848\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3584\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24840\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24835\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24835\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__24840\,
            I => \N__24830\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__24835\,
            I => \N__24830\
        );

    \I__3579\ : Span12Mux_v
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__3578\ : Odrv12
    port map (
            O => \N__24827\,
            I => \pid_alt.error_d_regZ0Z_20\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24821\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24821\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \pid_alt.un1_pid_prereg_236_1_cascade_\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__24806\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\
        );

    \I__3570\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24793\
        );

    \I__3569\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24793\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24793\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__24800\,
            I => \N__24790\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__24793\,
            I => \N__24787\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24782\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__24787\,
            I => \N__24779\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24774\
        );

    \I__3562\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24774\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24782\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__24779\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__24774\,
            I => \pid_alt.un1_pid_prereg_236_1\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__3557\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24755\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24755\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24762\,
            I => \N__24755\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24751\
        );

    \I__3553\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24747\
        );

    \I__3552\ : Span4Mux_h
    port map (
            O => \N__24751\,
            I => \N__24744\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24741\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__24747\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__24744\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24741\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__24734\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24717\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24717\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24717\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24717\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24714\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24711\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24717\,
            I => \N__24708\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24703\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24703\
        );

    \I__3537\ : Span4Mux_s3_h
    port map (
            O => \N__24708\,
            I => \N__24698\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__24703\,
            I => \N__24698\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__24698\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24692\,
            I => \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24686\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24686\,
            I => drone_altitude_1
        );

    \I__3530\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__24680\,
            I => drone_altitude_2
        );

    \I__3528\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24674\,
            I => drone_altitude_3
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__24671\,
            I => \N__24667\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__24670\,
            I => \N__24664\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24661\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24658\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__24661\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24658\,
            I => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\
        );

    \I__3520\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24644\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24644\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24644\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__3516\ : Span4Mux_h
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__3515\ : Span4Mux_v
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__24632\,
            I => \pid_alt.error_d_regZ0Z_7\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24620\
        );

    \I__3510\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24620\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24620\,
            I => \pid_alt.error_d_reg_prevZ0Z_7\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24611\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24611\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3504\ : Span4Mux_v
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__24602\,
            I => \pid_alt.error_p_regZ0Z_7\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24596\,
            I => \N__24593\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24593\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24584\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24584\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3496\ : Span4Mux_h
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__24578\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24571\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24568\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24560\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24560\
        );

    \I__3489\ : Span4Mux_v
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__24557\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__24554\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24545\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24545\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24541\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24538\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__24541\,
            I => \N__24535\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24538\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__24535\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24527\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24521\,
            I => \pid_alt.pid_preregZ0Z_20\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__24515\,
            I => \pid_alt.pid_preregZ0Z_19\
        );

    \I__3473\ : CascadeMux
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24506\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24500\,
            I => \pid_alt.pid_preregZ0Z_17\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24494\,
            I => \pid_alt.pid_preregZ0Z_21\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__24488\,
            I => \pid_alt.pid_preregZ0Z_15\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24479\,
            I => \pid_alt.pid_preregZ0Z_23\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24473\,
            I => \pid_alt.pid_preregZ0Z_18\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24467\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24463\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24460\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__24463\,
            I => \N__24457\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24454\
        );

    \I__3454\ : Span4Mux_h
    port map (
            O => \N__24457\,
            I => \N__24449\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__24454\,
            I => \N__24449\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__24449\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__24443\,
            I => \pid_alt.error_i_acumm_preregZ0Z_15\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24437\,
            I => \pid_alt.error_i_acumm_preregZ0Z_14\
        );

    \I__3447\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__24431\,
            I => \N__24428\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__24425\,
            I => \pid_alt.un1_reset_1_i_a5_0_9\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24419\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3441\ : Span4Mux_h
    port map (
            O => \N__24416\,
            I => \N__24413\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__24413\,
            I => \pid_alt.un1_reset_1_i_a5_0_8\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__24410\,
            I => \pid_alt.N_557_cascade_\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__24404\,
            I => \pid_alt.un1_reset_1_i_a5_0_10\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__24401\,
            I => \pid_alt.N_304_cascade_\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__24398\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__24392\,
            I => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\
        );

    \I__3432\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24386\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__24383\,
            I => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24374\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24370\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24367\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__24370\,
            I => \N__24364\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24367\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__24364\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24355\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__24358\,
            I => \N__24352\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24349\
        );

    \I__3419\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24346\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__24349\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__24346\,
            I => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24334\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24331\
        );

    \I__3413\ : Span4Mux_v
    port map (
            O => \N__24334\,
            I => \N__24328\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24331\,
            I => \N__24325\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__24328\,
            I => \N__24322\
        );

    \I__3410\ : Odrv12
    port map (
            O => \N__24325\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__3409\ : Odrv4
    port map (
            O => \N__24322\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24314\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__24311\,
            I => \N__24307\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24304\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__24307\,
            I => \N__24301\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__24304\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__24301\,
            I => \pid_alt.error_d_reg_prevZ0Z_8\
        );

    \I__3401\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__24293\,
            I => \N__24288\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24283\
        );

    \I__3398\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24283\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__24288\,
            I => \N__24280\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__3395\ : Span4Mux_v
    port map (
            O => \N__24280\,
            I => \N__24274\
        );

    \I__3394\ : Span12Mux_v
    port map (
            O => \N__24277\,
            I => \N__24271\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__24274\,
            I => \N__24268\
        );

    \I__3392\ : Odrv12
    port map (
            O => \N__24271\,
            I => \pid_alt.error_d_regZ0Z_8\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24268\,
            I => \pid_alt.error_d_regZ0Z_8\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24257\
        );

    \I__3389\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24257\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24257\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24251\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3385\ : Span4Mux_v
    port map (
            O => \N__24248\,
            I => \N__24243\
        );

    \I__3384\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24240\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__24246\,
            I => \N__24237\
        );

    \I__3382\ : Span4Mux_v
    port map (
            O => \N__24243\,
            I => \N__24232\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24232\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24229\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__24232\,
            I => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24229\,
            I => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\
        );

    \I__3377\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24221\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24216\
        );

    \I__3375\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24211\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24211\
        );

    \I__3373\ : Span4Mux_h
    port map (
            O => \N__24216\,
            I => \N__24208\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__24211\,
            I => \N__24205\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__24208\,
            I => \pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__24205\,
            I => \pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12\
        );

    \I__3369\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24196\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \N__24193\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24190\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24187\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__24190\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__24187\,
            I => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\
        );

    \I__3363\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__24179\,
            I => \N__24174\
        );

    \I__3361\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24171\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24177\,
            I => \N__24168\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__24174\,
            I => \N__24163\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24171\,
            I => \N__24163\
        );

    \I__3357\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24160\
        );

    \I__3356\ : Odrv4
    port map (
            O => \N__24163\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24160\,
            I => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24152\,
            I => \N__24147\
        );

    \I__3352\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24142\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24142\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__24147\,
            I => \N__24139\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__24142\,
            I => \N__24136\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__24139\,
            I => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__24136\,
            I => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24124\
        );

    \I__3344\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24121\
        );

    \I__3343\ : Span4Mux_h
    port map (
            O => \N__24124\,
            I => \N__24117\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24114\
        );

    \I__3341\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24111\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__24117\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__24114\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24111\,
            I => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\
        );

    \I__3337\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__24101\,
            I => \N__24096\
        );

    \I__3335\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24093\
        );

    \I__3334\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24090\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__24096\,
            I => \N__24087\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__24093\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__24090\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__24087\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__3329\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24077\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__24074\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24064\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24061\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__24064\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24061\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__3321\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24052\
        );

    \I__3320\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24049\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__24052\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__24049\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__24044\,
            I => \N__24040\
        );

    \I__3316\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24037\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24034\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__24037\,
            I => \N__24031\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__24034\,
            I => \N__24027\
        );

    \I__3312\ : Span12Mux_s11_v
    port map (
            O => \N__24031\,
            I => \N__24024\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24021\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__24027\,
            I => \N__24018\
        );

    \I__3309\ : Odrv12
    port map (
            O => \N__24024\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24021\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__24018\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__24004\
        );

    \I__3304\ : InMux
    port map (
            O => \N__24007\,
            I => \N__24001\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__24004\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__24001\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__23996\,
            I => \pid_alt.un1_reset_1_i_a5_0_7_cascade_\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__3299\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__3298\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23984\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__23984\,
            I => \pid_alt.error_d_reg_prevZ0Z_12\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23974\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__23977\,
            I => \N__23971\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23974\,
            I => \N__23968\
        );

    \I__3292\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23965\
        );

    \I__3291\ : Span4Mux_v
    port map (
            O => \N__23968\,
            I => \N__23962\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23959\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__23962\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__3288\ : Odrv12
    port map (
            O => \N__23959\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__23945\,
            I => \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\
        );

    \I__3283\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23939\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__3281\ : Span4Mux_v
    port map (
            O => \N__23936\,
            I => \N__23932\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23935\,
            I => \N__23929\
        );

    \I__3279\ : Span4Mux_h
    port map (
            O => \N__23932\,
            I => \N__23924\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23924\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__23918\,
            I => \pid_alt.error_p_regZ0Z_10\
        );

    \I__3274\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23911\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23908\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__23911\,
            I => \N__23905\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__23908\,
            I => \N__23902\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__23905\,
            I => \N__23899\
        );

    \I__3269\ : Span4Mux_v
    port map (
            O => \N__23902\,
            I => \N__23896\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__23899\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__23896\,
            I => \pid_alt.error_d_reg_prevZ0Z_10\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23886\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23883\
        );

    \I__3264\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23880\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__23886\,
            I => \N__23877\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23883\,
            I => \N__23874\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23880\,
            I => \N__23867\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__23877\,
            I => \N__23867\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__23874\,
            I => \N__23867\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__23864\,
            I => \pid_alt.error_d_regZ0Z_10\
        );

    \I__3256\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23858\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__23858\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__23855\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__23852\,
            I => \N__23849\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__23846\,
            I => \N__23842\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__23842\,
            I => \N__23836\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__23839\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__23836\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23825\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23825\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__23825\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23813\
        );

    \I__3242\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23813\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23813\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__23804\,
            I => \pid_alt.error_d_regZ0Z_11\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23792\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23792\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23792\,
            I => \pid_alt.error_d_reg_prevZ0Z_11\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23783\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23783\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__3229\ : Span12Mux_v
    port map (
            O => \N__23780\,
            I => \N__23777\
        );

    \I__3228\ : Odrv12
    port map (
            O => \N__23777\,
            I => \pid_alt.error_p_regZ0Z_11\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23768\
        );

    \I__3226\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23768\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__23768\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23756\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23756\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23756\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__23750\,
            I => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23741\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__23741\,
            I => \N__23737\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__23740\,
            I => \N__23733\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__23737\,
            I => \N__23730\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23725\
        );

    \I__3212\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23725\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__23730\,
            I => \N__23720\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23725\,
            I => \N__23720\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__23720\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__3208\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__23714\,
            I => \N__23710\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23706\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__23710\,
            I => \N__23701\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23698\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23706\,
            I => \N__23695\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23690\
        );

    \I__3201\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23690\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__23701\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23698\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__23695\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__23690\,
            I => \pid_alt.error_d_regZ0Z_0\
        );

    \I__3196\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23675\
        );

    \I__3194\ : Span4Mux_v
    port map (
            O => \N__23675\,
            I => \N__23672\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__23672\,
            I => \pid_alt.error_d_reg_prevZ0Z_0\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__23660\,
            I => \Commands_frame_decoder.state_ns_i_a2_0_2_0\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23652\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23647\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23644\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23652\,
            I => \N__23641\
        );

    \I__3184\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23638\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23635\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23647\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__23644\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__23641\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23638\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23635\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__23615\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_3_2\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23608\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23605\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23608\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23605\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__23600\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23594\,
            I => \N__23589\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23584\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23584\
        );

    \I__3164\ : Span4Mux_h
    port map (
            O => \N__23589\,
            I => \N__23579\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23579\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__23573\,
            I => \pid_alt.error_d_regZ0Z_12\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23570\,
            I => \N__23567\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__23564\,
            I => \Commands_frame_decoder.N_418\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23555\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23555\,
            I => \Commands_frame_decoder.N_382_2\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__23552\,
            I => \Commands_frame_decoder.N_383_cascade_\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23549\,
            I => \Commands_frame_decoder.state_ns_i_0_0_cascade_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23542\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23539\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23542\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23539\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23530\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23526\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23523\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23520\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23526\,
            I => \N__23515\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__23523\,
            I => \N__23515\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23520\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__23515\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23506\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23503\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23506\,
            I => \N__23498\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23498\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__23498\,
            I => \frame_decoder_CH4data_7\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__3132\ : Span4Mux_v
    port map (
            O => \N__23489\,
            I => \N__23486\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__23483\,
            I => \pid_side.error_8\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23480\,
            I => \bfn_4_22_0_\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__23471\,
            I => \drone_H_disp_side_i_9\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__3122\ : Span4Mux_h
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__23456\,
            I => \pid_side.error_9\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23453\,
            I => \pid_side.error_cry_4\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__23441\,
            I => \drone_H_disp_side_i_10\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__3112\ : Span4Mux_v
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__23426\,
            I => \pid_side.error_10\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23423\,
            I => \pid_side.error_cry_5\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23417\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__3107\ : Span4Mux_h
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__23411\,
            I => \N__23408\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23408\,
            I => \pid_side.error_11\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23405\,
            I => \pid_side.error_cry_6\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3100\ : Span4Mux_v
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__23390\,
            I => \pid_side.error_12\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23387\,
            I => \pid_side.error_cry_7\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__3094\ : Span4Mux_v
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__23372\,
            I => \pid_side.error_13\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23369\,
            I => \pid_side.error_cry_8\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__3088\ : Span4Mux_v
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__23354\,
            I => \pid_side.error_14\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23351\,
            I => \pid_side.error_cry_9\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23348\,
            I => \pid_side.error_cry_10\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__3082\ : Span12Mux_s4_h
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3081\ : Odrv12
    port map (
            O => \N__23336\,
            I => \pid_side.error_15\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__23324\,
            I => alt_kp_0
        );

    \I__3076\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23318\,
            I => \pid_side.error_axb_0\
        );

    \I__3074\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3072\ : Span4Mux_s2_h
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__3071\ : Span4Mux_v
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__23303\,
            I => \pid_side.error_1\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23300\,
            I => \pid_side.error_cry_0\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__23291\,
            I => \N__23288\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__23288\,
            I => \pid_side.error_2\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23285\,
            I => \pid_side.error_cry_1\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__3061\ : Span4Mux_s1_h
    port map (
            O => \N__23276\,
            I => \N__23273\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__23270\,
            I => \pid_side.error_3\
        );

    \I__3058\ : InMux
    port map (
            O => \N__23267\,
            I => \pid_side.error_cry_2\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__3055\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__3054\ : Odrv4
    port map (
            O => \N__23255\,
            I => \pid_side.error_4\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23252\,
            I => \pid_side.error_cry_3\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__23240\,
            I => \pid_side.error_5\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23237\,
            I => \pid_side.error_cry_0_0\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23228\
        );

    \I__3045\ : Span4Mux_s1_h
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__3044\ : Span4Mux_v
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__23222\,
            I => \pid_side.error_6\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23219\,
            I => \pid_side.error_cry_1_0\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__3039\ : Span4Mux_s1_h
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__23204\,
            I => \pid_side.error_7\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23201\,
            I => \pid_side.error_cry_2_0\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__23192\,
            I => \drone_H_disp_side_i_8\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__3031\ : InMux
    port map (
            O => \N__23186\,
            I => \N__23182\
        );

    \I__3030\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23179\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23173\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__23176\,
            I => \N__23170\
        );

    \I__3026\ : Span4Mux_v
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__23170\,
            I => \pid_alt.error_d_reg_prev_i_0\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__23167\,
            I => \pid_alt.error_d_reg_prev_i_0\
        );

    \I__3023\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23159\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__23159\,
            I => \dron_frame_decoder_1.drone_H_disp_side_8\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23153\,
            I => \dron_frame_decoder_1.drone_H_disp_side_9\
        );

    \I__3019\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23147\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__23147\,
            I => \dron_frame_decoder_1.drone_H_disp_side_10\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__23141\,
            I => \pid_alt.error_axbZ0Z_1\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23135\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__23132\,
            I => drone_altitude_12
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \N__23126\
        );

    \I__3011\ : InMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__23123\,
            I => \pid_alt.error_axbZ0Z_12\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23117\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__23114\,
            I => \N__23111\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__23111\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23108\,
            I => \pid_alt.un1_pid_prereg_0_cry_21\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__23105\,
            I => \N__23101\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23098\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23095\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23092\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23089\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__23092\,
            I => \N__23086\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__23086\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__23083\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__23078\,
            I => \N__23075\
        );

    \I__2994\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__23069\,
            I => \N__23066\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__23066\,
            I => \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\
        );

    \I__2990\ : InMux
    port map (
            O => \N__23063\,
            I => \bfn_4_18_0_\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23060\,
            I => \pid_alt.un1_pid_prereg_0_cry_23\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23054\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23054\,
            I => \pid_alt.error_axbZ0Z_13\
        );

    \I__2986\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23048\,
            I => drone_altitude_13
        );

    \I__2984\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__23042\,
            I => \pid_alt.error_axbZ0Z_14\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23036\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__23036\,
            I => drone_altitude_14
        );

    \I__2980\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__23030\,
            I => \pid_alt.error_axbZ0Z_2\
        );

    \I__2978\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23024\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__23024\,
            I => \pid_alt.error_axbZ0Z_3\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23017\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23014\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23011\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23014\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__2972\ : Odrv12
    port map (
            O => \N__23011\,
            I => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__23006\,
            I => \N__23003\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__22997\,
            I => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22994\,
            I => \pid_alt.un1_pid_prereg_0_cry_13\
        );

    \I__2966\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__22985\,
            I => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__22982\,
            I => \N__22978\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__22981\,
            I => \N__22975\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22972\
        );

    \I__2960\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22969\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__22972\,
            I => \N__22966\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22963\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__22966\,
            I => \N__22958\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__22963\,
            I => \N__22958\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__22958\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\
        );

    \I__2954\ : InMux
    port map (
            O => \N__22955\,
            I => \bfn_4_17_0_\
        );

    \I__2953\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__22949\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__22946\,
            I => \N__22942\
        );

    \I__2950\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22939\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22936\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__22939\,
            I => \N__22931\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22936\,
            I => \N__22931\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2945\ : Odrv4
    port map (
            O => \N__22928\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22925\,
            I => \pid_alt.un1_pid_prereg_0_cry_15\
        );

    \I__2943\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22919\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__22919\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__22916\,
            I => \N__22912\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__22915\,
            I => \N__22909\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22906\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22903\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__22906\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__22903\,
            I => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\
        );

    \I__2935\ : InMux
    port map (
            O => \N__22898\,
            I => \pid_alt.un1_pid_prereg_0_cry_16\
        );

    \I__2934\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__22889\,
            I => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__22886\,
            I => \N__22882\
        );

    \I__2930\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22876\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__22879\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__22876\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22871\,
            I => \pid_alt.un1_pid_prereg_0_cry_17\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22862\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__22862\,
            I => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__22859\,
            I => \N__22855\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__22858\,
            I => \N__22852\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22849\
        );

    \I__2919\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22846\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22849\,
            I => \N__22843\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22846\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2916\ : Odrv12
    port map (
            O => \N__22843\,
            I => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22838\,
            I => \pid_alt.un1_pid_prereg_0_cry_18\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22835\,
            I => \pid_alt.un1_pid_prereg_0_cry_19\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22832\,
            I => \pid_alt.un1_pid_prereg_0_cry_20\
        );

    \I__2912\ : InMux
    port map (
            O => \N__22829\,
            I => \pid_alt.un1_pid_prereg_0_cry_4\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__2909\ : Span4Mux_h
    port map (
            O => \N__22820\,
            I => \N__22817\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__22817\,
            I => \pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__22814\,
            I => \N__22810\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__22813\,
            I => \N__22807\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22804\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22801\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__22804\,
            I => \N__22798\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22795\
        );

    \I__2901\ : Span4Mux_h
    port map (
            O => \N__22798\,
            I => \N__22792\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__22792\,
            I => \pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__22789\,
            I => \pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4\
        );

    \I__2897\ : InMux
    port map (
            O => \N__22784\,
            I => \pid_alt.un1_pid_prereg_0_cry_5\
        );

    \I__2896\ : InMux
    port map (
            O => \N__22781\,
            I => \bfn_4_16_0_\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22778\,
            I => \pid_alt.un1_pid_prereg_0_cry_7\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__22769\,
            I => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\
        );

    \I__2891\ : InMux
    port map (
            O => \N__22766\,
            I => \pid_alt.un1_pid_prereg_0_cry_8\
        );

    \I__2890\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__22760\,
            I => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22750\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22747\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22744\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22747\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__22744\,
            I => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22739\,
            I => \pid_alt.un1_pid_prereg_0_cry_9\
        );

    \I__2881\ : InMux
    port map (
            O => \N__22736\,
            I => \pid_alt.un1_pid_prereg_0_cry_10\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2878\ : Odrv12
    port map (
            O => \N__22727\,
            I => \pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11\
        );

    \I__2877\ : InMux
    port map (
            O => \N__22724\,
            I => \pid_alt.un1_pid_prereg_0_cry_11\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__22715\,
            I => \pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22709\,
            I => \N__22705\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__22708\,
            I => \N__22702\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22699\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22702\,
            I => \N__22696\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__22699\,
            I => \N__22693\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22696\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11\
        );

    \I__2866\ : Odrv4
    port map (
            O => \N__22693\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11\
        );

    \I__2865\ : InMux
    port map (
            O => \N__22688\,
            I => \pid_alt.un1_pid_prereg_0_cry_12\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__22685\,
            I => \pid_alt.N_294_cascade_\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22677\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22667\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22680\,
            I => \N__22667\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22667\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22676\,
            I => \N__22667\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__22667\,
            I => \pid_alt.N_294\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22655\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22655\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22652\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__22652\,
            I => \N__22644\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22635\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22635\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22635\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22635\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__22647\,
            I => \N__22632\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__22644\,
            I => \N__22625\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22622\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22611\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22611\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22611\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22611\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22611\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__22625\,
            I => \pid_alt.N_295\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__22622\,
            I => \pid_alt.N_295\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22611\,
            I => \pid_alt.N_295\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22600\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22597\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22591\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22591\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22588\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__22591\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22588\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__22580\,
            I => \pid_alt.error_i_acummZ0Z_4\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2825\ : Span4Mux_s2_h
    port map (
            O => \N__22568\,
            I => \N__22564\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22561\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__22564\,
            I => \pid_alt.un1_pid_prereg_0\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22561\,
            I => \pid_alt.un1_pid_prereg_0\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__22544\,
            I => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22541\,
            I => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__22529\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22526\,
            I => \pid_alt.un1_pid_prereg_0_cry_0\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22517\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__22514\,
            I => \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22511\,
            I => \pid_alt.un1_pid_prereg_0_cry_1\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__2803\ : Span4Mux_h
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__22499\,
            I => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22496\,
            I => \pid_alt.un1_pid_prereg_0_cry_2\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22486\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22483\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22478\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22478\
        );

    \I__2795\ : Span4Mux_h
    port map (
            O => \N__22478\,
            I => \N__22475\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__22475\,
            I => \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2792\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__22463\,
            I => \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22460\,
            I => \pid_alt.un1_pid_prereg_0_cry_3\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__22451\,
            I => \pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__22448\,
            I => \N__22444\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22441\
        );

    \I__2783\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22438\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22433\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22433\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__22433\,
            I => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__22430\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22418\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22418\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22418\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2774\ : Span4Mux_h
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__22409\,
            I => \pid_alt.error_d_regZ0Z_14\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22397\
        );

    \I__2769\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22397\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22397\,
            I => \pid_alt.error_d_reg_prevZ0Z_14\
        );

    \I__2767\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22388\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22388\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__22382\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22376\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22376\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22367\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__22364\,
            I => \pid_alt.N_295_cascade_\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22358\,
            I => \pid_alt.error_i_acummZ0Z_1\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22352\,
            I => \pid_alt.error_i_acummZ0Z_2\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__22346\,
            I => \pid_alt.error_i_acummZ0Z_3\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22334\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22334\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__22334\,
            I => \pid_alt.m39_i_a2_3\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22327\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22322\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22322\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__22319\,
            I => \pid_alt.m39_i_a2_4\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22309\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22309\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22306\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22309\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__22306\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__2736\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22297\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22294\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__22297\,
            I => \N__22291\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__2732\ : Span12Mux_v
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__2731\ : Span12Mux_v
    port map (
            O => \N__22288\,
            I => \N__22282\
        );

    \I__2730\ : Odrv12
    port map (
            O => \N__22285\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__22282\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__2728\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22270\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22267\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__22270\,
            I => \N__22264\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22267\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__22264\,
            I => \pid_alt.error_d_reg_prevZ0Z_13\
        );

    \I__2722\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22254\
        );

    \I__2721\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22251\
        );

    \I__2720\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22248\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22243\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__22251\,
            I => \N__22243\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__22248\,
            I => \N__22240\
        );

    \I__2716\ : Span4Mux_v
    port map (
            O => \N__22243\,
            I => \N__22235\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__22240\,
            I => \N__22235\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__22232\,
            I => \pid_alt.error_d_regZ0Z_13\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22223\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22223\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__22223\,
            I => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22214\
        );

    \I__2708\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22214\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__22202\,
            I => \pid_alt.error_p_regZ0Z_12\
        );

    \I__2702\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__22196\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__22193\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\
        );

    \I__2699\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2697\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__22181\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__22178\,
            I => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\
        );

    \I__2694\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22172\,
            I => \N__22168\
        );

    \I__2692\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22165\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__22168\,
            I => \N__22162\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__22165\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__22162\,
            I => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22151\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22151\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__2684\ : Span4Mux_v
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__22139\,
            I => \pid_alt.error_p_regZ0Z_14\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__22136\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__2679\ : InMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__22127\,
            I => \Commands_frame_decoder.state_ns_0_a3_3_1\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__22121\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__22118\,
            I => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\
        );

    \I__2674\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22108\
        );

    \I__2673\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22108\
        );

    \I__2672\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22105\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22108\,
            I => \N__22102\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__22105\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__22102\,
            I => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\
        );

    \I__2668\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__22091\,
            I => \N__22086\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22083\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22080\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__22086\,
            I => \N__22077\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__22083\,
            I => \N__22074\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22071\
        );

    \I__2660\ : Sp12to4
    port map (
            O => \N__22077\,
            I => \N__22068\
        );

    \I__2659\ : Span4Mux_s3_h
    port map (
            O => \N__22074\,
            I => \N__22065\
        );

    \I__2658\ : Span4Mux_s3_h
    port map (
            O => \N__22071\,
            I => \N__22062\
        );

    \I__2657\ : Span12Mux_s3_h
    port map (
            O => \N__22068\,
            I => \N__22057\
        );

    \I__2656\ : Sp12to4
    port map (
            O => \N__22065\,
            I => \N__22057\
        );

    \I__2655\ : Span4Mux_v
    port map (
            O => \N__22062\,
            I => \N__22054\
        );

    \I__2654\ : Odrv12
    port map (
            O => \N__22057\,
            I => \pid_alt.error_14\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__22054\,
            I => \pid_alt.error_14\
        );

    \I__2652\ : InMux
    port map (
            O => \N__22049\,
            I => \pid_alt.error_cry_13\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__22043\,
            I => drone_altitude_15
        );

    \I__2649\ : InMux
    port map (
            O => \N__22040\,
            I => \pid_alt.error_cry_14\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22034\,
            I => \N__22029\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22026\
        );

    \I__2645\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22023\
        );

    \I__2644\ : Span12Mux_s7_v
    port map (
            O => \N__22029\,
            I => \N__22018\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__22026\,
            I => \N__22018\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22015\
        );

    \I__2641\ : Span12Mux_v
    port map (
            O => \N__22018\,
            I => \N__22010\
        );

    \I__2640\ : Span12Mux_s10_v
    port map (
            O => \N__22015\,
            I => \N__22010\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__22010\,
            I => \pid_alt.error_15\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__22004\,
            I => \dron_frame_decoder_1.drone_altitude_11\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__21998\,
            I => drone_altitude_i_11
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__21995\,
            I => \N__21991\
        );

    \I__2633\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21988\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21985\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21982\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__21985\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__2629\ : Odrv12
    port map (
            O => \N__21982\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__21971\,
            I => \N__21967\
        );

    \I__2625\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__21967\,
            I => \N__21961\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__21964\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__21961\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__2621\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2619\ : Span4Mux_s3_h
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__21947\,
            I => alt_kp_1
        );

    \I__2617\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__2615\ : Span4Mux_s3_h
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__21935\,
            I => alt_kp_7
        );

    \I__2613\ : CEMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21924\
        );

    \I__2611\ : CEMux
    port map (
            O => \N__21928\,
            I => \N__21921\
        );

    \I__2610\ : CEMux
    port map (
            O => \N__21927\,
            I => \N__21918\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__21924\,
            I => \N__21915\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__21921\,
            I => \N__21912\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__21918\,
            I => \N__21909\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__21915\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__21912\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__21909\,
            I => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__21902\,
            I => \N__21898\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__21901\,
            I => \N__21895\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21892\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21889\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21892\,
            I => alt_command_2
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__21889\,
            I => alt_command_2
        );

    \I__2597\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21880\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21877\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21874\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21877\,
            I => \N__21870\
        );

    \I__2593\ : Span4Mux_s3_h
    port map (
            O => \N__21874\,
            I => \N__21867\
        );

    \I__2592\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21864\
        );

    \I__2591\ : Span4Mux_s3_h
    port map (
            O => \N__21870\,
            I => \N__21861\
        );

    \I__2590\ : Span4Mux_v
    port map (
            O => \N__21867\,
            I => \N__21858\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__21864\,
            I => \N__21855\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__21861\,
            I => \N__21852\
        );

    \I__2587\ : Sp12to4
    port map (
            O => \N__21858\,
            I => \N__21847\
        );

    \I__2586\ : Span12Mux_s3_h
    port map (
            O => \N__21855\,
            I => \N__21847\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__21852\,
            I => \pid_alt.error_6\
        );

    \I__2584\ : Odrv12
    port map (
            O => \N__21847\,
            I => \pid_alt.error_6\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21842\,
            I => \pid_alt.error_cry_5\
        );

    \I__2582\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__21836\,
            I => drone_altitude_i_7
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__21833\,
            I => \N__21829\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__21832\,
            I => \N__21826\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21823\
        );

    \I__2577\ : InMux
    port map (
            O => \N__21826\,
            I => \N__21820\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21823\,
            I => alt_command_3
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__21820\,
            I => alt_command_3
        );

    \I__2574\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21807\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21804\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21801\
        );

    \I__2570\ : Span12Mux_s6_v
    port map (
            O => \N__21807\,
            I => \N__21796\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21796\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21801\,
            I => \N__21793\
        );

    \I__2567\ : Span12Mux_v
    port map (
            O => \N__21796\,
            I => \N__21788\
        );

    \I__2566\ : Span12Mux_s11_v
    port map (
            O => \N__21793\,
            I => \N__21788\
        );

    \I__2565\ : Odrv12
    port map (
            O => \N__21788\,
            I => \pid_alt.error_7\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21785\,
            I => \pid_alt.error_cry_6\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__21779\,
            I => drone_altitude_i_8
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__21770\,
            I => alt_command_4
        );

    \I__2558\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21760\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21756\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__21760\,
            I => \N__21753\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21750\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__21756\,
            I => \N__21747\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__21753\,
            I => \N__21744\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__21750\,
            I => \N__21741\
        );

    \I__2550\ : Span4Mux_s3_h
    port map (
            O => \N__21747\,
            I => \N__21738\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__21744\,
            I => \N__21735\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__21741\,
            I => \N__21732\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__21738\,
            I => \N__21729\
        );

    \I__2546\ : Span4Mux_h
    port map (
            O => \N__21735\,
            I => \N__21724\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__21732\,
            I => \N__21724\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__21729\,
            I => \pid_alt.error_8\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__21724\,
            I => \pid_alt.error_8\
        );

    \I__2542\ : InMux
    port map (
            O => \N__21719\,
            I => \bfn_3_20_0_\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__21713\,
            I => drone_altitude_i_9
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__2538\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__21704\,
            I => alt_command_5
        );

    \I__2536\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21693\
        );

    \I__2534\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21690\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21687\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__21693\,
            I => \N__21684\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21690\,
            I => \N__21681\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21678\
        );

    \I__2529\ : Sp12to4
    port map (
            O => \N__21684\,
            I => \N__21675\
        );

    \I__2528\ : Span4Mux_s3_h
    port map (
            O => \N__21681\,
            I => \N__21672\
        );

    \I__2527\ : Span4Mux_s3_h
    port map (
            O => \N__21678\,
            I => \N__21669\
        );

    \I__2526\ : Span12Mux_s3_h
    port map (
            O => \N__21675\,
            I => \N__21666\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__21672\,
            I => \N__21663\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__21669\,
            I => \N__21660\
        );

    \I__2523\ : Odrv12
    port map (
            O => \N__21666\,
            I => \pid_alt.error_9\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__21663\,
            I => \pid_alt.error_9\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__21660\,
            I => \pid_alt.error_9\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21653\,
            I => \pid_alt.error_cry_8\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21647\,
            I => drone_altitude_i_10
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21638\,
            I => alt_command_6
        );

    \I__2514\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21627\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21624\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21621\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__21627\,
            I => \N__21618\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21615\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21612\
        );

    \I__2507\ : Sp12to4
    port map (
            O => \N__21618\,
            I => \N__21609\
        );

    \I__2506\ : Span4Mux_s3_h
    port map (
            O => \N__21615\,
            I => \N__21606\
        );

    \I__2505\ : Span4Mux_s3_h
    port map (
            O => \N__21612\,
            I => \N__21603\
        );

    \I__2504\ : Span12Mux_s3_h
    port map (
            O => \N__21609\,
            I => \N__21600\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__21606\,
            I => \N__21597\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__21603\,
            I => \N__21594\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__21600\,
            I => \pid_alt.error_10\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__21597\,
            I => \pid_alt.error_10\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__21594\,
            I => \pid_alt.error_10\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21587\,
            I => \pid_alt.error_cry_9\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21578\,
            I => alt_command_7
        );

    \I__2494\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21570\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21567\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21564\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__21570\,
            I => \N__21561\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21567\,
            I => \N__21558\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21564\,
            I => \N__21555\
        );

    \I__2488\ : Span12Mux_s3_h
    port map (
            O => \N__21561\,
            I => \N__21552\
        );

    \I__2487\ : Span4Mux_s3_h
    port map (
            O => \N__21558\,
            I => \N__21549\
        );

    \I__2486\ : Span4Mux_s3_h
    port map (
            O => \N__21555\,
            I => \N__21546\
        );

    \I__2485\ : Span12Mux_v
    port map (
            O => \N__21552\,
            I => \N__21543\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__21549\,
            I => \N__21540\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__21546\,
            I => \N__21537\
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__21543\,
            I => \pid_alt.error_11\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__21540\,
            I => \pid_alt.error_11\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__21537\,
            I => \pid_alt.error_11\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21530\,
            I => \pid_alt.error_cry_10\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__21521\,
            I => \N__21516\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21513\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21510\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__21516\,
            I => \N__21507\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21504\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21510\,
            I => \N__21501\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__21507\,
            I => \N__21498\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__21504\,
            I => \N__21495\
        );

    \I__2468\ : Span12Mux_s3_h
    port map (
            O => \N__21501\,
            I => \N__21492\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__21498\,
            I => \N__21487\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__21495\,
            I => \N__21487\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__21492\,
            I => \pid_alt.error_12\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__21487\,
            I => \pid_alt.error_12\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21482\,
            I => \pid_alt.error_cry_11\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21476\,
            I => \N__21472\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__2459\ : Span4Mux_s2_h
    port map (
            O => \N__21472\,
            I => \N__21465\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21469\,
            I => \N__21462\
        );

    \I__2457\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21459\
        );

    \I__2456\ : Sp12to4
    port map (
            O => \N__21465\,
            I => \N__21456\
        );

    \I__2455\ : Span4Mux_s3_h
    port map (
            O => \N__21462\,
            I => \N__21453\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21450\
        );

    \I__2453\ : Span12Mux_v
    port map (
            O => \N__21456\,
            I => \N__21447\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__21453\,
            I => \N__21444\
        );

    \I__2451\ : Span12Mux_s3_h
    port map (
            O => \N__21450\,
            I => \N__21441\
        );

    \I__2450\ : Odrv12
    port map (
            O => \N__21447\,
            I => \pid_alt.error_13\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__21444\,
            I => \pid_alt.error_13\
        );

    \I__2448\ : Odrv12
    port map (
            O => \N__21441\,
            I => \pid_alt.error_13\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21434\,
            I => \pid_alt.error_cry_12\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21422\
        );

    \I__2445\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21422\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21422\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21422\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21416\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__21416\,
            I => \N__21413\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__21413\,
            I => \N__21409\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21412\,
            I => \N__21406\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__21409\,
            I => \N__21403\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21406\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1_0\
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__21403\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1_0\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21393\
        );

    \I__2434\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21390\
        );

    \I__2433\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21387\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21393\,
            I => \N__21384\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21381\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__21387\,
            I => \N__21378\
        );

    \I__2429\ : Span4Mux_s3_h
    port map (
            O => \N__21384\,
            I => \N__21375\
        );

    \I__2428\ : Span4Mux_v
    port map (
            O => \N__21381\,
            I => \N__21372\
        );

    \I__2427\ : Span4Mux_s3_h
    port map (
            O => \N__21378\,
            I => \N__21369\
        );

    \I__2426\ : Sp12to4
    port map (
            O => \N__21375\,
            I => \N__21366\
        );

    \I__2425\ : Span4Mux_h
    port map (
            O => \N__21372\,
            I => \N__21363\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__21369\,
            I => \N__21360\
        );

    \I__2423\ : Odrv12
    port map (
            O => \N__21366\,
            I => \pid_alt.error_1\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__21363\,
            I => \pid_alt.error_1\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__21360\,
            I => \pid_alt.error_1\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21353\,
            I => \pid_alt.error_cry_0\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21347\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__21344\,
            I => \N__21339\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21336\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21333\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__21339\,
            I => \N__21328\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21336\,
            I => \N__21328\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21333\,
            I => \N__21325\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__21328\,
            I => \N__21322\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__21325\,
            I => \N__21319\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__21322\,
            I => \N__21314\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__21319\,
            I => \N__21314\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__21314\,
            I => \pid_alt.error_2\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21311\,
            I => \pid_alt.error_cry_1\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21300\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21297\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21303\,
            I => \N__21294\
        );

    \I__2401\ : Span4Mux_s3_h
    port map (
            O => \N__21300\,
            I => \N__21291\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21288\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21285\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__21291\,
            I => \N__21282\
        );

    \I__2397\ : Span4Mux_s3_h
    port map (
            O => \N__21288\,
            I => \N__21279\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__21285\,
            I => \N__21276\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__21282\,
            I => \N__21273\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__21279\,
            I => \N__21270\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__21276\,
            I => \N__21267\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__21273\,
            I => \pid_alt.error_3\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__21270\,
            I => \pid_alt.error_3\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__21267\,
            I => \pid_alt.error_3\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21260\,
            I => \pid_alt.error_cry_2\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__21257\,
            I => \N__21253\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__21256\,
            I => \N__21250\
        );

    \I__2386\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21247\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21244\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__21247\,
            I => alt_command_0
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__21244\,
            I => alt_command_0
        );

    \I__2382\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21236\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__2380\ : Span4Mux_s1_h
    port map (
            O => \N__21233\,
            I => \N__21229\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21226\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__21229\,
            I => \N__21220\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21220\
        );

    \I__2376\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21217\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__21220\,
            I => \N__21214\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__21217\,
            I => \N__21211\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__21214\,
            I => \N__21208\
        );

    \I__2372\ : Span4Mux_s3_h
    port map (
            O => \N__21211\,
            I => \N__21205\
        );

    \I__2371\ : Span4Mux_s1_h
    port map (
            O => \N__21208\,
            I => \N__21202\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__21205\,
            I => \N__21199\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__21202\,
            I => \pid_alt.error_4\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__21199\,
            I => \pid_alt.error_4\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21194\,
            I => \pid_alt.error_cry_3\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21188\,
            I => drone_altitude_i_5
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__21185\,
            I => \N__21181\
        );

    \I__2363\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21178\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21175\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__21178\,
            I => alt_command_1
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21175\,
            I => alt_command_1
        );

    \I__2359\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21166\
        );

    \I__2358\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21162\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21159\
        );

    \I__2356\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21156\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__21162\,
            I => \N__21153\
        );

    \I__2354\ : Span12Mux_s2_h
    port map (
            O => \N__21159\,
            I => \N__21150\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21147\
        );

    \I__2352\ : Span4Mux_s3_h
    port map (
            O => \N__21153\,
            I => \N__21144\
        );

    \I__2351\ : Span12Mux_v
    port map (
            O => \N__21150\,
            I => \N__21141\
        );

    \I__2350\ : Span12Mux_s3_h
    port map (
            O => \N__21147\,
            I => \N__21138\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__21144\,
            I => \N__21135\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__21141\,
            I => \pid_alt.error_5\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__21138\,
            I => \pid_alt.error_5\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__21135\,
            I => \pid_alt.error_5\
        );

    \I__2345\ : InMux
    port map (
            O => \N__21128\,
            I => \pid_alt.error_cry_4\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__21122\,
            I => drone_altitude_i_6
        );

    \I__2342\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21110\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21110\
        );

    \I__2340\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21110\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__2338\ : Span12Mux_s10_h
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__2337\ : Span12Mux_v
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2336\ : Odrv12
    port map (
            O => \N__21101\,
            I => \pid_alt.error_d_regZ0Z_16\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__2334\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21089\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21089\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21089\,
            I => \pid_alt.error_d_reg_prevZ0Z_16\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21080\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21080\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__2328\ : Span4Mux_h
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__21074\,
            I => \N__21071\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__21071\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__21065\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__21062\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__21059\,
            I => \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__21056\,
            I => \Commands_frame_decoder.source_CH1data8_cascade_\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__2318\ : Span4Mux_h
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__21041\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__2315\ : InMux
    port map (
            O => \N__21038\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_18\
        );

    \I__2314\ : InMux
    port map (
            O => \N__21035\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21026\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21026\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__2310\ : Span4Mux_h
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__21017\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21014\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21008\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__21005\,
            I => \N__21001\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20998\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__20998\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__20995\,
            I => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20982\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20979\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20976\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__20982\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__20979\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__20976\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\
        );

    \I__2292\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20965\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20962\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20959\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__20962\,
            I => \N__20954\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__20959\,
            I => \N__20954\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__20951\,
            I => \pid_alt.error_p_regZ0Z_17\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__20945\,
            I => \N__20941\
        );

    \I__2283\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20938\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__20941\,
            I => \N__20935\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__20938\,
            I => \pid_alt.error_d_reg_prevZ0Z_17\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__20935\,
            I => \pid_alt.error_d_reg_prevZ0Z_17\
        );

    \I__2279\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20922\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20917\
        );

    \I__2276\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20917\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__20922\,
            I => \N__20914\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20911\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__20914\,
            I => \N__20908\
        );

    \I__2272\ : Span12Mux_v
    port map (
            O => \N__20911\,
            I => \N__20905\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__20908\,
            I => \N__20902\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__20905\,
            I => \pid_alt.error_d_regZ0Z_17\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__20902\,
            I => \pid_alt.error_d_regZ0Z_17\
        );

    \I__2268\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__20894\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__20891\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20882\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__20882\,
            I => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__2261\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__20867\,
            I => \pid_alt.error_i_regZ0Z_11\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20864\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_10\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__20855\,
            I => \N__20852\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__20846\,
            I => \pid_alt.error_i_regZ0Z_12\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20843\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_11\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__2248\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__20825\,
            I => \pid_alt.error_i_regZ0Z_13\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20822\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_12\
        );

    \I__2242\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__2240\ : Span4Mux_v
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__20807\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20804\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_13\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__20795\,
            I => \N__20792\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__20789\,
            I => \pid_alt.error_i_regZ0Z_15\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20786\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_14\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__20771\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20768\,
            I => \bfn_3_16_0_\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__2222\ : Span4Mux_v
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__20753\,
            I => \pid_alt.error_i_regZ0Z_17\
        );

    \I__2219\ : InMux
    port map (
            O => \N__20750\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_16\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20744\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__2216\ : Span12Mux_v
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__2215\ : Odrv12
    port map (
            O => \N__20738\,
            I => \pid_alt.error_i_regZ0Z_18\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20735\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_17\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__20720\,
            I => \pid_alt.error_i_regZ0Z_3\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20717\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_2\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__20699\,
            I => \pid_alt.error_i_regZ0Z_4\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20691\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20686\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20686\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20691\,
            I => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__20686\,
            I => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20681\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_3\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__2193\ : Span4Mux_v
    port map (
            O => \N__20672\,
            I => \N__20669\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__20669\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20661\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20656\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20656\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20661\,
            I => \pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20656\,
            I => \pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20651\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_4\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20644\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20641\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20638\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__20641\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__20638\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2177\ : Span4Mux_v
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__20621\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20618\,
            I => \N__20612\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20612\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20608\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20605\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__20608\,
            I => \N__20602\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__20605\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__20602\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20597\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20585\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__20582\,
            I => \pid_alt.error_i_regZ0Z_7\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20579\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20572\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20569\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20572\,
            I => \N__20566\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20569\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__20566\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20555\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__20546\,
            I => \pid_alt.error_i_regZ0Z_8\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20543\,
            I => \bfn_3_15_0_\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20536\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20533\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20530\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20533\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__20530\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__20525\,
            I => \N__20522\
        );

    \I__2143\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20519\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__20513\,
            I => \N__20510\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__20510\,
            I => \pid_alt.error_i_regZ0Z_9\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20502\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20497\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20497\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20502\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20497\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20492\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20485\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20482\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__20479\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__20474\,
            I => \N__20471\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__20462\,
            I => \pid_alt.error_i_regZ0Z_10\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20459\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20456\,
            I => \N__20451\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20446\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20446\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20451\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20446\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20436\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__20440\,
            I => \N__20433\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20439\,
            I => \N__20430\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20427\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20422\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20422\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__20427\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__20422\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20406\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20403\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20400\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__20406\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20403\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20400\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20390\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20390\,
            I => \N__20385\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20382\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20379\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__20385\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20382\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20379\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__20363\,
            I => \pid_alt.error_i_regZ0Z_1\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20360\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_0\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__20345\,
            I => \pid_alt.error_i_regZ0Z_2\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20342\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_1\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__20333\,
            I => \pid_alt.O_2_6\
        );

    \I__2079\ : CEMux
    port map (
            O => \N__20330\,
            I => \N__20279\
        );

    \I__2078\ : CEMux
    port map (
            O => \N__20329\,
            I => \N__20279\
        );

    \I__2077\ : CEMux
    port map (
            O => \N__20328\,
            I => \N__20279\
        );

    \I__2076\ : CEMux
    port map (
            O => \N__20327\,
            I => \N__20279\
        );

    \I__2075\ : CEMux
    port map (
            O => \N__20326\,
            I => \N__20279\
        );

    \I__2074\ : CEMux
    port map (
            O => \N__20325\,
            I => \N__20279\
        );

    \I__2073\ : CEMux
    port map (
            O => \N__20324\,
            I => \N__20279\
        );

    \I__2072\ : CEMux
    port map (
            O => \N__20323\,
            I => \N__20279\
        );

    \I__2071\ : CEMux
    port map (
            O => \N__20322\,
            I => \N__20279\
        );

    \I__2070\ : CEMux
    port map (
            O => \N__20321\,
            I => \N__20279\
        );

    \I__2069\ : CEMux
    port map (
            O => \N__20320\,
            I => \N__20279\
        );

    \I__2068\ : CEMux
    port map (
            O => \N__20319\,
            I => \N__20279\
        );

    \I__2067\ : CEMux
    port map (
            O => \N__20318\,
            I => \N__20279\
        );

    \I__2066\ : CEMux
    port map (
            O => \N__20317\,
            I => \N__20279\
        );

    \I__2065\ : CEMux
    port map (
            O => \N__20316\,
            I => \N__20279\
        );

    \I__2064\ : CEMux
    port map (
            O => \N__20315\,
            I => \N__20279\
        );

    \I__2063\ : CEMux
    port map (
            O => \N__20314\,
            I => \N__20279\
        );

    \I__2062\ : GlobalMux
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__2061\ : gio2CtrlBuf
    port map (
            O => \N__20276\,
            I => \pid_alt.N_850_0_g\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__2058\ : Span4Mux_s2_h
    port map (
            O => \N__20267\,
            I => \N__20264\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__20264\,
            I => alt_kp_2
        );

    \I__2056\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20258\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__2053\ : Sp12to4
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__2052\ : Odrv12
    port map (
            O => \N__20249\,
            I => alt_kp_3
        );

    \I__2051\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__2049\ : Span4Mux_s3_h
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__20237\,
            I => alt_kp_5
        );

    \I__2047\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__2045\ : Span4Mux_s2_h
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__20225\,
            I => alt_kp_6
        );

    \I__2043\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__20219\,
            I => \N__20216\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__20213\,
            I => alt_kd_3
        );

    \I__2039\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__2037\ : Span4Mux_s3_h
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__20201\,
            I => alt_kd_0
        );

    \I__2035\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__2033\ : Span4Mux_s3_h
    port map (
            O => \N__20192\,
            I => \N__20189\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__20189\,
            I => alt_kd_4
        );

    \I__2031\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20183\,
            I => \dron_frame_decoder_1.drone_altitude_10\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__20177\,
            I => \dron_frame_decoder_1.drone_altitude_8\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__20171\,
            I => \dron_frame_decoder_1.drone_altitude_9\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20162\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__2022\ : Span4Mux_v
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__20156\,
            I => \pid_alt.error_p_regZ0Z_5\
        );

    \I__2020\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20147\
        );

    \I__2019\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20147\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__20147\,
            I => \pid_alt.error_d_reg_prevZ0Z_5\
        );

    \I__2017\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20135\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20135\
        );

    \I__2015\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20135\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__2013\ : Span12Mux_v
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__20129\,
            I => \pid_alt.error_d_regZ0Z_5\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__2010\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20117\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20117\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__20114\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\
        );

    \I__2006\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20105\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20105\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__20099\,
            I => \pid_alt.error_p_regZ0Z_6\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20090\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20090\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__20090\,
            I => \pid_alt.error_d_reg_prevZ0Z_6\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20078\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20078\
        );

    \I__1996\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20078\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20075\
        );

    \I__1994\ : Span12Mux_v
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__1993\ : Odrv12
    port map (
            O => \N__20072\,
            I => \pid_alt.error_d_regZ0Z_6\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__20060\,
            I => \pid_side.O_0_24\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__20048\,
            I => \pid_side.O_0_13\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20039\
        );

    \I__1983\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20039\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__20039\,
            I => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\
        );

    \I__1981\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20027\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20027\
        );

    \I__1979\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20027\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__20015\,
            I => \pid_alt.error_d_regZ0Z_18\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__20012\,
            I => \N__20009\
        );

    \I__1972\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20003\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20003\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__20003\,
            I => \pid_alt.error_d_reg_prevZ0Z_18\
        );

    \I__1969\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19994\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19994\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__19988\,
            I => \pid_alt.error_p_regZ0Z_18\
        );

    \I__1964\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__19982\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\
        );

    \I__1962\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19973\
        );

    \I__1961\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19973\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__19970\,
            I => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__19967\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\
        );

    \I__1957\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__19961\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19949\
        );

    \I__1953\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19949\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__19949\,
            I => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__19946\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19934\
        );

    \I__1949\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19934\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19941\,
            I => \N__19934\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__1945\ : Span4Mux_v
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__19925\,
            I => \pid_alt.error_d_regZ0Z_9\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19913\
        );

    \I__1941\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19913\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__19913\,
            I => \pid_alt.error_d_reg_prevZ0Z_9\
        );

    \I__1939\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19904\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19904\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__19895\,
            I => \pid_alt.error_p_regZ0Z_9\
        );

    \I__1933\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__19889\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\
        );

    \I__1931\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19880\
        );

    \I__1930\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19880\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__1928\ : Span4Mux_h
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__19874\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__19871\,
            I => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__19865\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__19862\,
            I => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19856\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\
        );

    \I__1920\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19847\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19847\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19847\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19835\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19835\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__19826\,
            I => \pid_alt.error_p_regZ0Z_4\
        );

    \I__1910\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19817\
        );

    \I__1909\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19817\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__19814\,
            I => \pid_alt.error_d_reg_prevZ0Z_4\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19803\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19798\
        );

    \I__1903\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19798\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__19803\,
            I => \N__19793\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19793\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__19793\,
            I => \pid_alt.error_d_regZ0Z_4\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__19790\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__19784\,
            I => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__1894\ : Span4Mux_s2_h
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__19772\,
            I => alt_ki_5
        );

    \I__1892\ : InMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__19760\,
            I => \pid_alt.O_2_5\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__19748\,
            I => \pid_alt.O_2_4\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__1882\ : Span4Mux_s2_h
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__19736\,
            I => alt_kd_5
        );

    \I__1880\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__1878\ : Span4Mux_s2_h
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__19724\,
            I => alt_kd_1
        );

    \I__1876\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__19712\,
            I => \pid_alt.O_1_9\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__19700\,
            I => alt_ki_0
        );

    \I__1868\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19694\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__1866\ : Span4Mux_s2_h
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__19688\,
            I => alt_ki_4
        );

    \I__1864\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19682\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__19676\,
            I => alt_ki_1
        );

    \I__1860\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__19667\,
            I => \N__19664\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__19664\,
            I => alt_ki_2
        );

    \I__1856\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__1854\ : Span4Mux_s2_h
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__19652\,
            I => alt_ki_3
        );

    \I__1852\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__19646\,
            I => \pid_alt.O_3_9\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19640\,
            I => \pid_alt.O_3_10\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__19634\,
            I => \pid_alt.O_3_11\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__19628\,
            I => \pid_alt.O_3_13\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19622\,
            I => \N__19619\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__19616\,
            I => \pid_alt.O_1_8\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__1838\ : Span4Mux_h
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__19604\,
            I => \pid_alt.O_1_11\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__19595\,
            I => alt_kd_6
        );

    \I__1833\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19589\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__19586\,
            I => alt_kd_2
        );

    \I__1830\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19580\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1828\ : Span4Mux_s2_h
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__19574\,
            I => alt_kd_7
        );

    \I__1826\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19568\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__19562\,
            I => \pid_alt.O_3_24\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__19553\,
            I => \pid_alt.O_3_20\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__19547\,
            I => \N__19544\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__19544\,
            I => \pid_alt.O_3_21\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__19535\,
            I => \pid_alt.O_3_22\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19526\,
            I => \pid_alt.O_3_23\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__19517\,
            I => \pid_alt.O_3_15\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__19508\,
            I => \pid_alt.O_3_19\
        );

    \I__1804\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__19502\,
            I => \pid_alt.O_3_14\
        );

    \I__1802\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__19496\,
            I => \pid_alt.O_3_8\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__19490\,
            I => \N__19487\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__19487\,
            I => \pid_alt.O_3_6\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \N__19480\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19476\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19469\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19469\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19466\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19461\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19474\,
            I => \N__19461\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19458\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__19466\,
            I => \N__19453\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19453\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19458\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19453\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__1785\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__19445\,
            I => \pid_alt.O_3_7\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19442\,
            I => \N__19438\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19434\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19431\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19428\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19425\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__19431\,
            I => \N__19420\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N__19420\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__19425\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__19420\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__1774\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__19412\,
            I => \pid_alt.O_3_5\
        );

    \I__1772\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19399\
        );

    \I__1771\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19399\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19394\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19394\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19405\,
            I => \N__19389\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19389\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19382\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__19394\,
            I => \N__19382\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__19389\,
            I => \N__19382\
        );

    \I__1763\ : Odrv12
    port map (
            O => \N__19382\,
            I => \pid_alt.error_p_regZ0Z_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__19373\,
            I => \pid_alt.O_3_12\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__19364\,
            I => \pid_alt.O_3_16\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__19355\,
            I => \pid_alt.O_3_17\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__19346\,
            I => \pid_alt.O_3_18\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19340\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__19337\,
            I => \N__19332\
        );

    \I__1747\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19324\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19324\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19319\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19319\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19314\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19314\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19324\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19319\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__19314\,
            I => \pid_alt.error_d_reg_prevZ0Z_1\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19296\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19296\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19289\
        );

    \I__1735\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19289\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19289\
        );

    \I__1733\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19284\
        );

    \I__1732\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19284\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19277\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__19289\,
            I => \N__19277\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__19284\,
            I => \N__19277\
        );

    \I__1728\ : Odrv12
    port map (
            O => \N__19277\,
            I => \pid_alt.error_d_regZ0Z_1\
        );

    \I__1727\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__19271\,
            I => \pid_alt.N_3_1\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__19265\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19262\,
            I => \N__19254\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19261\,
            I => \N__19249\
        );

    \I__1721\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19249\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19242\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19242\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19242\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19235\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__19249\,
            I => \N__19235\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__19242\,
            I => \N__19235\
        );

    \I__1714\ : Odrv12
    port map (
            O => \N__19235\,
            I => \pid_alt.error_d_regZ0Z_2\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__19229\,
            I => \N__19222\
        );

    \I__1711\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19217\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19217\
        );

    \I__1709\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19212\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19212\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__19222\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__19217\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__19212\,
            I => \pid_alt.error_d_reg_prevZ0Z_2\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__19199\,
            I => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__19190\,
            I => \N__19185\
        );

    \I__1698\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19180\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19180\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__19185\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__19180\,
            I => \pid_alt.error_d_reg_prevZ0Z_3\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19165\
        );

    \I__1693\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19165\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19165\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19162\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19159\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__19162\,
            I => \N__19154\
        );

    \I__1688\ : Span12Mux_v
    port map (
            O => \N__19159\,
            I => \N__19154\
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__19154\,
            I => \pid_alt.error_d_regZ0Z_3\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__19145\,
            I => \pid_alt.g0_4_0\
        );

    \I__1683\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__19139\,
            I => \pid_alt.N_1505_i_0\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__19133\,
            I => \pid_alt.N_3_0\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__1678\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__19124\,
            I => \pid_alt.N_1507_0\
        );

    \I__1676\ : InMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19118\,
            I => \pid_alt.N_5\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__19112\,
            I => \pid_alt.N_1511_0\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__19109\,
            I => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\
        );

    \I__1671\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19102\
        );

    \I__1670\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19097\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19102\,
            I => \N__19094\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19089\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19089\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19097\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__19094\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__19089\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19079\,
            I => \pid_alt.N_1505_i_1\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1660\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__19070\,
            I => \pid_alt.N_1507_1\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__19067\,
            I => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\
        );

    \I__1657\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__1655\ : Span12Mux_s4_h
    port map (
            O => \N__19058\,
            I => \N__19055\
        );

    \I__1654\ : Span12Mux_v
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__1653\ : Odrv12
    port map (
            O => \N__19052\,
            I => \pid_alt.O_1_4\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__1649\ : Span4Mux_s1_h
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__19037\,
            I => \pid_alt.O_3_4\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__1646\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__19028\,
            I => \pid_alt.N_1505_i\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \pid_alt.N_1505_i_cascade_\
        );

    \I__1643\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__19019\,
            I => \pid_alt.un1_pid_prereg_0_axb_2_1\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__19016\,
            I => \pid_alt.N_1513_0_cascade_\
        );

    \I__1640\ : InMux
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19010\,
            I => \pid_side.O_0_11\
        );

    \I__1638\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__19004\,
            I => \pid_side.O_0_6\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__18998\,
            I => \pid_side.O_0_17\
        );

    \I__1634\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__18992\,
            I => \pid_side.O_0_16\
        );

    \I__1632\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__18986\,
            I => \pid_side.O_0_12\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18980\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__18980\,
            I => \pid_side.O_0_20\
        );

    \I__1628\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__18974\,
            I => \pid_side.O_0_21\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__18968\,
            I => \pid_side.O_0_22\
        );

    \I__1624\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18962\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__18962\,
            I => \pid_side.O_0_9\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__18953\,
            I => \pid_side.O_0_19\
        );

    \I__1619\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__18947\,
            I => \pid_side.O_0_14\
        );

    \I__1617\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__18941\,
            I => \pid_side.O_0_8\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__18935\,
            I => \pid_side.O_0_10\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__18926\,
            I => \pid_side.O_0_23\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__18917\,
            I => \pid_side.O_0_15\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__18908\,
            I => \pid_side.O_0_18\
        );

    \I__1604\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__18902\,
            I => \pid_alt.O_2_17\
        );

    \I__1602\ : InMux
    port map (
            O => \N__18899\,
            I => \N__18896\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__1600\ : Span4Mux_v
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__18890\,
            I => \pid_alt.O_1_6\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18884\,
            I => \pid_alt.O_2_12\
        );

    \I__1596\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__18878\,
            I => \pid_alt.O_2_19\
        );

    \I__1594\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__18872\,
            I => \pid_alt.O_2_14\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__18866\,
            I => \pid_alt.O_2_15\
        );

    \I__1590\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__1588\ : Span4Mux_h
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__18851\,
            I => \pid_alt.O_1_5\
        );

    \I__1585\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18845\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__1583\ : Span4Mux_h
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__18839\,
            I => \pid_alt.O_2_22\
        );

    \I__1581\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__18833\,
            I => \pid_alt.O_2_11\
        );

    \I__1579\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__18824\,
            I => \pid_alt.O_2_24\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__18818\,
            I => \pid_alt.O_2_7\
        );

    \I__1574\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__18812\,
            I => \pid_alt.O_2_8\
        );

    \I__1572\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__18803\,
            I => \pid_alt.O_2_23\
        );

    \I__1569\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__18797\,
            I => \pid_alt.O_2_10\
        );

    \I__1567\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18791\,
            I => \pid_alt.O_2_9\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__18782\,
            I => \pid_alt.O_2_16\
        );

    \I__1562\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__18773\,
            I => \pid_alt.O_1_24\
        );

    \I__1559\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__18767\,
            I => \pid_alt.O_1_13\
        );

    \I__1557\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__18761\,
            I => \pid_alt.O_1_14\
        );

    \I__1555\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__18755\,
            I => \pid_alt.O_1_10\
        );

    \I__1553\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__18749\,
            I => \pid_alt.O_1_21\
        );

    \I__1551\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__18740\,
            I => \pid_alt.O_2_13\
        );

    \I__1548\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__18731\,
            I => \pid_alt.O_2_21\
        );

    \I__1545\ : InMux
    port map (
            O => \N__18728\,
            I => \N__18725\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__18722\,
            I => \pid_alt.O_2_18\
        );

    \I__1542\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__18713\,
            I => \pid_alt.O_2_20\
        );

    \I__1539\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__18707\,
            I => \pid_alt.O_1_15\
        );

    \I__1537\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__18698\,
            I => \pid_alt.O_1_16\
        );

    \I__1534\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__18689\,
            I => \pid_alt.O_1_17\
        );

    \I__1531\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__18680\,
            I => \pid_alt.O_1_19\
        );

    \I__1528\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__18671\,
            I => \pid_alt.O_1_20\
        );

    \I__1525\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18665\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__18665\,
            I => \pid_alt.O_1_7\
        );

    \I__1523\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18659\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__18659\,
            I => \pid_alt.O_1_22\
        );

    \I__1521\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__18653\,
            I => \pid_alt.O_1_23\
        );

    \I__1519\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__18647\,
            I => \pid_alt.O_1_18\
        );

    \I__1517\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__18641\,
            I => \pid_alt.O_1_12\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_6\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_14\,
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_22\,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_15_12_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.un1_pid_prereg_cry_8\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.un1_pid_prereg_cry_16\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_18_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_22_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.un1_pid_prereg_cry_8\,
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.un1_pid_prereg_cry_16\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_cry_7\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_4_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_21_0_\
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_side.error_cry_3_0\,
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_front.error_cry_3_0\,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \dron_frame_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Commands_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_8_8_0_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__42143\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_661_g\
        );

    \pid_alt.state_RNICP2N1_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25910\,
            GLOBALBUFFEROUTPUT => \pid_alt.N_850_0_g\
        );

    \reset_module_System.reset_RNITC69_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__48314\,
            GLOBALBUFFEROUTPUT => \N_851_g\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__49034\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pid_alt.state_RNIH1EN_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31118\,
            GLOBALBUFFEROUTPUT => \pid_alt.state_0_g_0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_8_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18644\,
            lcout => \pid_alt.error_d_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_11_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_12_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_13_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18695\,
            lcout => \pid_alt.error_d_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_15_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18686\,
            lcout => \pid_alt.error_d_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_16_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18677\,
            lcout => \pid_alt.error_d_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51542\,
            ce => \N__20330\,
            sr => \N__50717\
        );

    \pid_alt.error_d_reg_esr_3_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_18_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18662\,
            lcout => \pid_alt.error_d_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_19_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18656\,
            lcout => \pid_alt.error_d_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_14_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18650\,
            lcout => \pid_alt.error_d_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_20_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18779\,
            lcout => \pid_alt.error_d_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_9_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18770\,
            lcout => \pid_alt.error_d_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_10_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18764\,
            lcout => \pid_alt.error_d_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_6_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18758\,
            lcout => \pid_alt.error_d_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51540\,
            ce => \N__20328\,
            sr => \N__50715\
        );

    \pid_alt.error_d_reg_esr_17_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18752\,
            lcout => \pid_alt.error_d_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51537\,
            ce => \N__20327\,
            sr => \N__50714\
        );

    \pid_alt.error_i_reg_esr_9_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18746\,
            lcout => \pid_alt.error_i_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51531\,
            ce => \N__20325\,
            sr => \N__50712\
        );

    \pid_alt.error_i_reg_esr_17_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18737\,
            lcout => \pid_alt.error_i_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51531\,
            ce => \N__20325\,
            sr => \N__50712\
        );

    \pid_alt.error_i_reg_esr_14_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18728\,
            lcout => \pid_alt.error_i_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51531\,
            ce => \N__20325\,
            sr => \N__50712\
        );

    \pid_alt.error_i_reg_esr_16_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18719\,
            lcout => \pid_alt.error_i_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51531\,
            ce => \N__20325\,
            sr => \N__50712\
        );

    \pid_alt.error_i_reg_esr_18_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \pid_alt.error_i_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51531\,
            ce => \N__20325\,
            sr => \N__50712\
        );

    \pid_alt.error_i_reg_esr_7_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18836\,
            lcout => \pid_alt.error_i_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_20_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18830\,
            lcout => \pid_alt.error_i_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_3_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18821\,
            lcout => \pid_alt.error_i_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_4_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18815\,
            lcout => \pid_alt.error_i_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_19_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18809\,
            lcout => \pid_alt.error_i_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_6_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18800\,
            lcout => \pid_alt.error_i_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_5_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18794\,
            lcout => \pid_alt.error_i_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_12_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18788\,
            lcout => \pid_alt.error_i_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51527\,
            ce => \N__20324\,
            sr => \N__50711\
        );

    \pid_alt.error_i_reg_esr_13_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18905\,
            lcout => \pid_alt.error_i_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_d_reg_esr_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18899\,
            lcout => \pid_alt.error_d_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_i_reg_esr_8_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18887\,
            lcout => \pid_alt.error_i_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_i_reg_esr_15_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18881\,
            lcout => \pid_alt.error_i_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_i_reg_esr_10_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18875\,
            lcout => \pid_alt.error_i_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_i_reg_esr_11_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18869\,
            lcout => \pid_alt.error_i_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51522\,
            ce => \N__20323\,
            sr => \N__50710\
        );

    \pid_alt.error_d_reg_esr_1_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18863\,
            lcout => \pid_alt.error_d_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51517\,
            ce => \N__20321\,
            sr => \N__50708\
        );

    \pid_alt.error_d_reg_prev_esr_13_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22259\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51511\,
            ce => \N__25564\,
            sr => \N__49537\
        );

    \pid_alt.error_d_reg_prev_esr_4_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19811\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51511\,
            ce => \N__25564\,
            sr => \N__49537\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_3_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19441\,
            in1 => \N__19196\,
            in2 => \_gnd_net_\,
            in3 => \N__19172\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_13_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__22301\,
            in1 => \N__22273\,
            in2 => \_gnd_net_\,
            in3 => \N__22258\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHMZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_5_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50204\,
            in1 => \N__30853\,
            in2 => \_gnd_net_\,
            in3 => \N__18965\,
            lcout => \pid_side.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_15_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18959\,
            in1 => \N__50206\,
            in2 => \_gnd_net_\,
            in3 => \N__28260\,
            lcout => \pid_side.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_10_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50202\,
            in1 => \N__29391\,
            in2 => \_gnd_net_\,
            in3 => \N__18950\,
            lcout => \pid_side.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_4_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28368\,
            in1 => \N__50208\,
            in2 => \_gnd_net_\,
            in3 => \N__18944\,
            lcout => \pid_side.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_6_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18938\,
            in1 => \_gnd_net_\,
            in2 => \N__50226\,
            in3 => \N__28336\,
            lcout => \pid_side.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_19_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28293\,
            in1 => \N__50207\,
            in2 => \_gnd_net_\,
            in3 => \N__18932\,
            lcout => \pid_side.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_11_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50203\,
            in1 => \N__28408\,
            in2 => \_gnd_net_\,
            in3 => \N__18923\,
            lcout => \pid_side.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_14_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28219\,
            in1 => \N__50205\,
            in2 => \_gnd_net_\,
            in3 => \N__18914\,
            lcout => \pid_side.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51494\,
            ce => 'H',
            sr => \N__50705\
        );

    \pid_side.error_p_reg_7_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30354\,
            in1 => \N__50217\,
            in2 => \_gnd_net_\,
            in3 => \N__19013\,
            lcout => \pid_side.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_2_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__19007\,
            in1 => \_gnd_net_\,
            in2 => \N__50227\,
            in3 => \N__34701\,
            lcout => \pid_side.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_13_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30825\,
            in1 => \N__50215\,
            in2 => \_gnd_net_\,
            in3 => \N__19001\,
            lcout => \pid_side.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_12_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50212\,
            in1 => \N__28695\,
            in2 => \_gnd_net_\,
            in3 => \N__18995\,
            lcout => \pid_side.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_8_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28438\,
            in1 => \N__50218\,
            in2 => \_gnd_net_\,
            in3 => \N__18989\,
            lcout => \pid_side.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_16_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50213\,
            in1 => \N__30909\,
            in2 => \_gnd_net_\,
            in3 => \N__18983\,
            lcout => \pid_side.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_17_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28176\,
            in1 => \N__50216\,
            in2 => \_gnd_net_\,
            in3 => \N__18977\,
            lcout => \pid_side.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_side.error_p_reg_18_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50214\,
            in1 => \N__28645\,
            in2 => \_gnd_net_\,
            in3 => \N__18971\,
            lcout => \pid_side.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51485\,
            ce => 'H',
            sr => \N__50704\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_3_2_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19483\,
            in1 => \N__19232\,
            in2 => \_gnd_net_\,
            in3 => \N__19262\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI0J511_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIIGU44_1_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24182\,
            in2 => \N__19067\,
            in3 => \N__19022\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIIGU44Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI3SMI1_0_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__22577\,
            in1 => \N__19101\,
            in2 => \_gnd_net_\,
            in3 => \N__23705\,
            lcout => \pid_alt.error_p_reg_esr_RNI3SMI1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_1_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19336\,
            in1 => \N__19409\,
            in2 => \N__19034\,
            in3 => \N__19307\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL2AQ1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_0_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19064\,
            lcout => \pid_alt.error_d_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51472\,
            ce => \N__20318\,
            sr => \N__50703\
        );

    \pid_alt.error_p_reg_esr_0_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19049\,
            lcout => \pid_alt.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51472\,
            ce => \N__20318\,
            sr => \N__50703\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19100\,
            in2 => \_gnd_net_\,
            in3 => \N__23704\,
            lcout => \pid_alt.N_1505_i\,
            ltout => \pid_alt.N_1505_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL2AQ1_0_1_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010110010"
        )
    port map (
            in0 => \N__19335\,
            in1 => \N__19408\,
            in2 => \N__19025\,
            in3 => \N__19306\,
            lcout => \pid_alt.un1_pid_prereg_0_axb_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5LS3_0_1_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110001"
        )
    port map (
            in0 => \N__19142\,
            in1 => \N__19121\,
            in2 => \N__19130\,
            in3 => \N__19136\,
            lcout => OPEN,
            ltout => \pid_alt.N_1513_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNILE0V5_3_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011010100"
        )
    port map (
            in0 => \N__19151\,
            in1 => \N__19115\,
            in2 => \N__19016\,
            in3 => \N__19442\,
            lcout => \pid_alt.error_p_reg_esr_RNILE0V5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_0_0_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19105\,
            in2 => \_gnd_net_\,
            in3 => \N__23709\,
            lcout => \pid_alt.N_1505_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_1_1_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19406\,
            in1 => \N__19331\,
            in2 => \_gnd_net_\,
            in3 => \N__19303\,
            lcout => \pid_alt.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_1_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__19304\,
            in1 => \_gnd_net_\,
            in2 => \N__19337\,
            in3 => \N__19407\,
            lcout => \pid_alt.N_1507_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_1_2_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19227\,
            in1 => \N__19479\,
            in2 => \_gnd_net_\,
            in3 => \N__19260\,
            lcout => \pid_alt.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111010"
        )
    port map (
            in0 => \N__19261\,
            in1 => \_gnd_net_\,
            in2 => \N__19484\,
            in3 => \N__19228\,
            lcout => \pid_alt.N_1511_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_1_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19305\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51459\,
            ce => \N__25575\,
            sr => \N__49579\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5LS3_1_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110001"
        )
    port map (
            in0 => \N__19082\,
            in1 => \N__19343\,
            in2 => \N__19076\,
            in3 => \N__19274\,
            lcout => OPEN,
            ltout => \pid_alt.error_d_reg_prev_esr_RNII5LS3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNILDG87_2_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__19205\,
            in2 => \N__19109\,
            in3 => \N__19268\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNILDG87Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIOI4P_1_0_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19106\,
            in2 => \_gnd_net_\,
            in3 => \N__23713\,
            lcout => \pid_alt.N_1505_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_0_1_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19405\,
            in1 => \N__19330\,
            in2 => \_gnd_net_\,
            in3 => \N__19302\,
            lcout => \pid_alt.N_1507_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_2_2_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19474\,
            in1 => \N__19225\,
            in2 => \_gnd_net_\,
            in3 => \N__19257\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNITF511_2_1_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19404\,
            in1 => \N__19329\,
            in2 => \_gnd_net_\,
            in3 => \N__19301\,
            lcout => \pid_alt.N_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI0J511_0_2_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19475\,
            in1 => \N__19226\,
            in2 => \_gnd_net_\,
            in3 => \N__19258\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI0J511_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_2_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51442\,
            ce => \N__25576\,
            sr => \N__49587\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_17_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__20968\,
            in1 => \N__20944\,
            in2 => \_gnd_net_\,
            in3 => \N__20925\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IMZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_17_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51428\,
            ce => \N__25577\,
            sr => \N__49596\
        );

    \pid_alt.error_d_reg_prev_esr_RNI3M511_0_3_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19437\,
            in1 => \N__19188\,
            in2 => \_gnd_net_\,
            in3 => \N__19173\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI3M511_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_3_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51428\,
            ce => \N__25577\,
            sr => \N__49596\
        );

    \pid_alt.error_d_reg_prev_esr_RNIE77K_3_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19189\,
            in2 => \_gnd_net_\,
            in3 => \N__19174\,
            lcout => \pid_alt.g0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_8_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24337\,
            in1 => \N__24310\,
            in2 => \_gnd_net_\,
            in3 => \N__24291\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_8_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51428\,
            ce => \N__25577\,
            sr => \N__49596\
        );

    \pid_alt.error_p_reg_esr_2_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19493\,
            lcout => \pid_alt.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51414\,
            ce => \N__20317\,
            sr => \N__50701\
        );

    \pid_alt.error_p_reg_esr_3_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19448\,
            lcout => \pid_alt.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_1_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19415\,
            lcout => \pid_alt.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_8_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \pid_alt.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_12_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19370\,
            lcout => \pid_alt.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_13_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19361\,
            lcout => \pid_alt.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_14_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19352\,
            lcout => \pid_alt.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_20_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19571\,
            lcout => \pid_alt.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51400\,
            ce => \N__20316\,
            sr => \N__50700\
        );

    \pid_alt.error_p_reg_esr_16_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19559\,
            lcout => \pid_alt.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_17_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19550\,
            lcout => \pid_alt.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_18_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19541\,
            lcout => \pid_alt.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_19_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19532\,
            lcout => \pid_alt.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_11_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19523\,
            lcout => \pid_alt.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_15_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_10_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19505\,
            lcout => \pid_alt.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_4_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19499\,
            lcout => \pid_alt.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51385\,
            ce => \N__20315\,
            sr => \N__50699\
        );

    \pid_alt.error_p_reg_esr_5_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19649\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51374\,
            ce => \N__20314\,
            sr => \N__50698\
        );

    \pid_alt.error_p_reg_esr_6_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19643\,
            lcout => \pid_alt.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51374\,
            ce => \N__20314\,
            sr => \N__50698\
        );

    \pid_alt.error_p_reg_esr_7_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19637\,
            lcout => \pid_alt.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51374\,
            ce => \N__20314\,
            sr => \N__50698\
        );

    \pid_alt.error_p_reg_esr_9_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19631\,
            lcout => \pid_alt.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51374\,
            ce => \N__20314\,
            sr => \N__50698\
        );

    \pid_alt.error_d_reg_esr_4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19625\,
            lcout => \pid_alt.error_d_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51541\,
            ce => \N__20329\,
            sr => \N__50716\
        );

    \pid_alt.error_d_reg_esr_7_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19613\,
            lcout => \pid_alt.error_d_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51541\,
            ce => \N__20329\,
            sr => \N__50716\
        );

    \Commands_frame_decoder.source_alt_kd_6_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40110\,
            lcout => alt_kd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51538\,
            ce => \N__21927\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39500\,
            in2 => \_gnd_net_\,
            in3 => \N__50823\,
            lcout => alt_kd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51538\,
            ce => \N__21927\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_7_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40012\,
            in2 => \_gnd_net_\,
            in3 => \N__50825\,
            lcout => alt_kd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51538\,
            ce => \N__21927\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_5_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40273\,
            in2 => \_gnd_net_\,
            in3 => \N__50819\,
            lcout => alt_kd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51535\,
            ce => \N__21932\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39626\,
            in2 => \_gnd_net_\,
            in3 => \N__50818\,
            lcout => alt_kd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51535\,
            ce => \N__21932\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_esr_5_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19721\,
            lcout => \pid_alt.error_d_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51532\,
            ce => \N__20326\,
            sr => \N__50713\
        );

    \Commands_frame_decoder.source_alt_ki_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39749\,
            in2 => \_gnd_net_\,
            in3 => \N__50817\,
            lcout => alt_ki_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51528\,
            ce => \N__38841\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40395\,
            in2 => \_gnd_net_\,
            in3 => \N__50815\,
            lcout => alt_ki_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51523\,
            ce => \N__38832\,
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25393\,
            in2 => \_gnd_net_\,
            in3 => \N__23509\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39625\,
            in2 => \_gnd_net_\,
            in3 => \N__50812\,
            lcout => alt_ki_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51523\,
            ce => \N__38832\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_2_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39488\,
            lcout => alt_ki_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51523\,
            ce => \N__38832\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_3_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39362\,
            in2 => \_gnd_net_\,
            in3 => \N__50814\,
            lcout => alt_ki_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51523\,
            ce => \N__38832\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_5_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40262\,
            lcout => alt_ki_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51523\,
            ce => \N__38832\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_10_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23889\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51518\,
            ce => \N__25557\,
            sr => \N__49518\
        );

    \pid_alt.error_i_reg_esr_1_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19769\,
            lcout => \pid_alt.error_i_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51512\,
            ce => \N__20320\,
            sr => \N__50707\
        );

    \pid_alt.error_i_reg_esr_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19757\,
            lcout => \pid_alt.error_i_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51505\,
            ce => \N__20319\,
            sr => \N__50706\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI8HDV_8_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__20389\,
            in2 => \N__33377\,
            in3 => \N__20410\,
            lcout => \pid_alt.m39_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_8_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24373\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51495\,
            ce => \N__25565\,
            sr => \N__49538\
        );

    \pid_alt.error_i_acumm_prereg_esr_9_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20507\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51495\,
            ce => \N__25565\,
            sr => \N__49538\
        );

    \pid_alt.error_i_acumm_prereg_esr_13_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22113\,
            lcout => \pid_alt.error_i_acumm7lto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51495\,
            ce => \N__25565\,
            sr => \N__49538\
        );

    \pid_alt.error_i_acumm_prereg_esr_21_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51495\,
            ce => \N__25565\,
            sr => \N__49538\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_0_20_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24801\,
            in1 => \N__24762\,
            in2 => \_gnd_net_\,
            in3 => \N__24728\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_1_20_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24730\,
            in1 => \_gnd_net_\,
            in2 => \N__24767\,
            in3 => \N__24803\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12_1Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS0U12_20_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__24802\,
            in1 => \N__24763\,
            in2 => \_gnd_net_\,
            in3 => \N__24729\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS0U12Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI11TA9_3_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19859\,
            in1 => \N__19852\,
            in2 => \N__22493\,
            in3 => \N__20694\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI11TA9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_0_4_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__19840\,
            in1 => \N__19822\,
            in2 => \_gnd_net_\,
            in3 => \N__19806\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI6P511_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICISB3_3_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19853\,
            in2 => \N__19844\,
            in3 => \N__20695\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICISB3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_0_10_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__23935\,
            in1 => \N__23914\,
            in2 => \_gnd_net_\,
            in3 => \N__23890\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHM_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI6P511_4_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19841\,
            in1 => \N__19823\,
            in2 => \_gnd_net_\,
            in3 => \N__19807\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI6P511Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI1FQN6_4_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__22447\,
            in1 => \N__20122\,
            in2 => \N__19790\,
            in3 => \N__20664\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI1FQN6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNILSTB3_4_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__20665\,
            in1 => \_gnd_net_\,
            in2 => \N__20126\,
            in3 => \N__19787\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNILSTB3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_9_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19909\,
            in1 => \N__19918\,
            in2 => \_gnd_net_\,
            in3 => \N__19941\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIL8611Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAR62_9_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21004\,
            in2 => \N__19946\,
            in3 => \N__20986\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAR62Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_9_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19943\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51473\,
            ce => \N__25569\,
            sr => \N__49550\
        );

    \pid_alt.error_d_reg_prev_esr_RNIG75T2_8_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19892\,
            in1 => \N__19886\,
            in2 => \_gnd_net_\,
            in3 => \N__20506\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIG75T2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL8611_0_9_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__19942\,
            in1 => \_gnd_net_\,
            in2 => \N__19922\,
            in3 => \N__19910\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIL8611_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIN49Q5_8_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__24359\,
            in1 => \N__19885\,
            in2 => \N__19871\,
            in3 => \N__20505\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIN49Q5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8IQ14_18_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20044\,
            in1 => \N__19868\,
            in2 => \N__22858\,
            in3 => \N__25713\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8IQ14Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_18_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__19999\,
            in1 => \N__20008\,
            in2 => \_gnd_net_\,
            in3 => \N__20034\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IMZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOTT02_18_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__20045\,
            in1 => \_gnd_net_\,
            in2 => \N__19862\,
            in3 => \N__25714\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOTT02Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_0_19_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24466\,
            in1 => \N__24890\,
            in2 => \_gnd_net_\,
            in3 => \N__24910\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IM_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_18_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51461\,
            ce => \N__25572\,
            sr => \N__49560\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGKS02_17_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__19985\,
            in1 => \N__19979\,
            in2 => \_gnd_net_\,
            in3 => \N__25684\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGKS02Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI53IM_0_18_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__20035\,
            in1 => \_gnd_net_\,
            in2 => \N__20012\,
            in3 => \N__20000\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI53IM_0Z0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOVN14_17_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__22885\,
            in1 => \N__19978\,
            in2 => \N__19967\,
            in3 => \N__25683\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOVN14Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIA5V86_5_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19954\,
            in1 => \N__19964\,
            in2 => \N__22814\,
            in3 => \N__20617\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIA5V86Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_0_6_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20110\,
            in1 => \N__20095\,
            in2 => \_gnd_net_\,
            in3 => \N__20085\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNICV511_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIL81T2_5_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__19955\,
            in1 => \_gnd_net_\,
            in2 => \N__19958\,
            in3 => \N__20618\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIL81T2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_5_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__20153\,
            in2 => \_gnd_net_\,
            in3 => \N__20143\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_5_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51443\,
            ce => \N__25573\,
            sr => \N__49568\
        );

    \pid_alt.error_d_reg_prev_esr_RNI9S511_0_5_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20167\,
            in1 => \N__20152\,
            in2 => \_gnd_net_\,
            in3 => \N__20142\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI9S511_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_6_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20087\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51443\,
            ce => \N__25573\,
            sr => \N__49568\
        );

    \pid_alt.error_d_reg_prev_esr_RNICV511_6_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__20111\,
            in1 => \N__20096\,
            in2 => \_gnd_net_\,
            in3 => \N__20086\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICV511Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_20_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28137\,
            in1 => \_gnd_net_\,
            in2 => \N__50228\,
            in3 => \N__20069\,
            lcout => \pid_side.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51429\,
            ce => 'H',
            sr => \N__50702\
        );

    \pid_side.error_p_reg_9_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27894\,
            in1 => \N__50222\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \pid_side.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51429\,
            ce => 'H',
            sr => \N__50702\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25160\,
            lcout => drone_altitude_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25151\,
            lcout => drone_altitude_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25796\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20180\,
            lcout => drone_altitude_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20174\,
            lcout => drone_altitude_i_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20186\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_i_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_10_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37130\,
            lcout => \dron_frame_decoder_1.drone_altitude_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \dron_frame_decoder_1.source_Altitude_esr_11_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37052\,
            lcout => \dron_frame_decoder_1.drone_altitude_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \dron_frame_decoder_1.source_Altitude_esr_12_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36946\,
            lcout => drone_altitude_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \dron_frame_decoder_1.source_Altitude_esr_15_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36632\,
            lcout => drone_altitude_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \dron_frame_decoder_1.source_Altitude_esr_8_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42611\,
            lcout => \dron_frame_decoder_1.drone_altitude_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \dron_frame_decoder_1.source_Altitude_esr_9_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36808\,
            lcout => \dron_frame_decoder_1.drone_altitude_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51417\,
            ce => \N__25823\,
            sr => \N__49588\
        );

    \Commands_frame_decoder.source_CH1data_esr_4_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40396\,
            lcout => alt_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51402\,
            ce => \N__25880\,
            sr => \N__49597\
        );

    \Commands_frame_decoder.source_CH1data_esr_5_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40250\,
            lcout => alt_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51402\,
            ce => \N__25880\,
            sr => \N__49597\
        );

    \Commands_frame_decoder.source_CH1data_esr_6_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40142\,
            lcout => alt_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51402\,
            ce => \N__25880\,
            sr => \N__49597\
        );

    \Commands_frame_decoder.source_CH1data_esr_7_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40011\,
            lcout => alt_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51402\,
            ce => \N__25880\,
            sr => \N__49597\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50806\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39527\,
            lcout => alt_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51376\,
            ce => \N__25952\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_3_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50807\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39380\,
            lcout => alt_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51376\,
            ce => \N__25952\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40272\,
            in2 => \_gnd_net_\,
            in3 => \N__50805\,
            lcout => alt_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51376\,
            ce => \N__25952\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_5_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50808\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40141\,
            lcout => alt_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51376\,
            ce => \N__25952\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_3_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39334\,
            lcout => alt_kd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51539\,
            ce => \N__21928\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_0_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39769\,
            in2 => \_gnd_net_\,
            in3 => \N__50820\,
            lcout => alt_kd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51539\,
            ce => \N__21928\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kd_4_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40379\,
            in2 => \_gnd_net_\,
            in3 => \N__50822\,
            lcout => alt_kd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51539\,
            ce => \N__21928\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_2_0_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__39742\,
            in1 => \N__23651\,
            in2 => \N__39497\,
            in3 => \N__21419\,
            lcout => \Commands_frame_decoder.N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_2_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20339\,
            lcout => \pid_alt.error_i_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51519\,
            ce => \N__20322\,
            sr => \N__50709\
        );

    \Commands_frame_decoder.source_offset4data_esr_6_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40122\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51513\,
            ce => \N__26963\,
            sr => \N__49515\
        );

    \pid_alt.error_i_acumm_10_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__20441\,
            in1 => \N__20488\,
            in2 => \N__31948\,
            in3 => \N__22648\,
            lcout => \pid_alt.error_i_acummZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51506\,
            ce => 'H',
            sr => \N__33225\
        );

    \pid_alt.error_i_acumm_6_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__20456\,
            in1 => \N__20647\,
            in2 => \N__31949\,
            in3 => \N__22649\,
            lcout => \pid_alt.error_i_acummZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51506\,
            ce => 'H',
            sr => \N__33225\
        );

    \pid_alt.error_i_acumm_8_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__20393\,
            in1 => \N__20575\,
            in2 => \N__31950\,
            in3 => \N__22650\,
            lcout => \pid_alt.error_i_acummZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51506\,
            ce => 'H',
            sr => \N__33225\
        );

    \pid_alt.error_i_acumm_9_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__22651\,
            in1 => \N__31910\,
            in2 => \N__20417\,
            in3 => \N__20539\,
            lcout => \pid_alt.error_i_acummZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51506\,
            ce => 'H',
            sr => \N__33225\
        );

    \pid_alt.pid_prereg_esr_RNIL6HQ_3_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31466\,
            in2 => \_gnd_net_\,
            in3 => \N__31892\,
            lcout => \pid_alt.N_306_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI08CV_10_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20455\,
            in1 => \N__23736\,
            in2 => \N__20440\,
            in3 => \N__24030\,
            lcout => \pid_alt.m39_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20611\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51496\,
            ce => \N__25561\,
            sr => \N__49523\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIGERC1_10_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20454\,
            in1 => \N__22314\,
            in2 => \N__20439\,
            in3 => \N__22596\,
            lcout => \pid_alt.un1_reset_1_i_a5_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20696\,
            lcout => \pid_alt.error_i_acumm7lto4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51496\,
            ce => \N__25561\,
            sr => \N__49523\
        );

    \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20666\,
            lcout => \pid_alt.error_i_acumm7lto5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51496\,
            ce => \N__25561\,
            sr => \N__49523\
        );

    \pid_alt.error_i_acumm_prereg_esr_10_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51496\,
            ce => \N__25561\,
            sr => \N__49523\
        );

    \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24544\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51496\,
            ce => \N__25561\,
            sr => \N__49523\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI6ECV_11_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20409\,
            in1 => \N__20388\,
            in2 => \N__23740\,
            in3 => \N__24104\,
            lcout => \pid_alt.un1_reset_1_i_a5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIB9IP_0_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24988\,
            in2 => \N__25015\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.un1_pid_prereg_0\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIQMD91_1_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22361\,
            in2 => \N__20372\,
            in3 => \N__20360\,
            lcout => \pid_alt.error_i_acumm_esr_RNIQMD91Z0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNITQE91_2_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22355\,
            in2 => \N__20357\,
            in3 => \N__20342\,
            lcout => \pid_alt.error_i_acumm_esr_RNITQE91Z0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI0VF91_3_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22349\,
            in2 => \N__20732\,
            in3 => \N__20717\,
            lcout => \pid_alt.error_i_acumm_esr_RNI0VF91Z0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI33H91_4_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22583\,
            in2 => \N__20714\,
            in3 => \N__20681\,
            lcout => \pid_alt.error_i_acumm_esr_RNI33H91Z0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNI67I91_5_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20678\,
            in2 => \N__22373\,
            in3 => \N__20651\,
            lcout => \pid_alt.error_i_acumm_esr_RNI67I91Z0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20648\,
            in2 => \N__20633\,
            in3 => \N__20597\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_5_c_RNI0DLQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21977\,
            in2 => \N__20594\,
            in3 => \N__20579\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_6_c_RNI3HMQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20576\,
            in2 => \N__20561\,
            in3 => \N__20543\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_7_c_RNI6LNQ\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_8_c_RNI9POQ_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20540\,
            in2 => \N__20525\,
            in3 => \N__20492\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_8_c_RNI9POQ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_9_c_RNIQN3F_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20489\,
            in2 => \N__20474\,
            in3 => \N__20459\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_9_c_RNIQN3F\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI4NMP_11_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21994\,
            in2 => \N__20879\,
            in3 => \N__20864\,
            lcout => \pid_alt.error_i_reg_esr_RNI4NMPZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIG2KM_12_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24080\,
            in2 => \N__20861\,
            in3 => \N__20843\,
            lcout => \pid_alt.error_i_acumm_esr_RNIG2KMZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_RNIJ6LM_13_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33281\,
            in2 => \N__20840\,
            in3 => \N__20822\,
            lcout => \pid_alt.error_i_acumm_esr_RNIJ6LMZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI15KJ_14_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20819\,
            in2 => \_gnd_net_\,
            in3 => \N__20804\,
            lcout => \pid_alt.error_i_reg_esr_RNI15KJZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI38LJ_15_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20801\,
            in2 => \_gnd_net_\,
            in3 => \N__20786\,
            lcout => \pid_alt.error_i_reg_esr_RNI38LJZ0Z_15\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI5BMJ_16_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20783\,
            in2 => \_gnd_net_\,
            in3 => \N__20768\,
            lcout => \pid_alt.error_i_reg_esr_RNI5BMJZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI7ENJ_17_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20765\,
            in2 => \_gnd_net_\,
            in3 => \N__20750\,
            lcout => \pid_alt.error_i_reg_esr_RNI7ENJZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNI9HOJ_18_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20747\,
            in2 => \_gnd_net_\,
            in3 => \N__20735\,
            lcout => \pid_alt.error_i_reg_esr_RNI9HOJZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_RNIBKPJ_19_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21053\,
            in2 => \_gnd_net_\,
            in3 => \N__21038\,
            lcout => \pid_alt.error_i_reg_esr_RNIBKPJZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21031\,
            in2 => \_gnd_net_\,
            in3 => \N__21035\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_19_c_RNI4FRJ\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_20_c_RNISVKK_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21014\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_20_c_RNISVKK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICI045_9_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__21011\,
            in1 => \N__22753\,
            in2 => \N__21005\,
            in3 => \N__20985\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICI045Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI88G14_14_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22175\,
            in1 => \N__22190\,
            in2 => \N__22982\,
            in3 => \N__24120\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI88G14Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8DL14_16_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20897\,
            in1 => \N__25659\,
            in2 => \N__22916\,
            in3 => \N__20887\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8DL14Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI20IM_0_17_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__20969\,
            in1 => \N__20948\,
            in2 => \_gnd_net_\,
            in3 => \N__20930\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI20IM_0Z0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI8BR02_16_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25660\,
            in2 => \N__20891\,
            in3 => \N__20888\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI8BR02Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_16_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__21085\,
            in1 => \N__21094\,
            in2 => \_gnd_net_\,
            in3 => \N__21117\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHMZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_16_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51444\,
            ce => \N__25570\,
            sr => \N__49551\
        );

    \pid_alt.error_d_reg_prev_esr_RNI02Q02_15_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__21068\,
            in1 => \N__25597\,
            in2 => \_gnd_net_\,
            in3 => \N__28538\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI02Q02Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIVSHM_0_16_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__21118\,
            in1 => \_gnd_net_\,
            in2 => \N__21098\,
            in3 => \N__21086\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIVSHM_0Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOQI14_15_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__22945\,
            in1 => \N__25596\,
            in2 => \N__21062\,
            in3 => \N__28537\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOQI14Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto3_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__39498\,
            in1 => \N__39364\,
            in2 => \_gnd_net_\,
            in3 => \N__39633\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto7_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40138\,
            in1 => \N__40400\,
            in2 => \N__21059\,
            in3 => \N__21412\,
            lcout => \Commands_frame_decoder.source_CH1data8\,
            ltout => \Commands_frame_decoder.source_CH1data8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_1_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__25497\,
            in1 => \N__21184\,
            in2 => \N__21056\,
            in3 => \N__39634\,
            lcout => alt_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51430\,
            ce => 'H',
            sr => \N__49561\
        );

    \Commands_frame_decoder.source_CH1data_2_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__21430\,
            in1 => \N__39499\,
            in2 => \N__21902\,
            in3 => \N__25498\,
            lcout => alt_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51430\,
            ce => 'H',
            sr => \N__49561\
        );

    \Commands_frame_decoder.source_CH1data_3_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__25499\,
            in1 => \N__39365\,
            in2 => \N__21833\,
            in3 => \N__21431\,
            lcout => alt_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51430\,
            ce => 'H',
            sr => \N__49561\
        );

    \Commands_frame_decoder.source_CH1data_0_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__21429\,
            in1 => \N__39770\,
            in2 => \N__21257\,
            in3 => \N__25496\,
            lcout => alt_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51430\,
            ce => 'H',
            sr => \N__49561\
        );

    \Commands_frame_decoder.source_CH1data8lto7_1_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39994\,
            in2 => \_gnd_net_\,
            in3 => \N__40257\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \pid_alt.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_RNI1N2F_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23144\,
            in2 => \_gnd_net_\,
            in3 => \N__21353\,
            lcout => \pid_alt.error_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_0\,
            carryout => \pid_alt.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_1_c_RNI3Q3F_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23033\,
            in2 => \_gnd_net_\,
            in3 => \N__21311\,
            lcout => \pid_alt.error_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_1\,
            carryout => \pid_alt.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_2_c_RNI5T4F_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23027\,
            in2 => \_gnd_net_\,
            in3 => \N__21260\,
            lcout => \pid_alt.error_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_2\,
            carryout => \pid_alt.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_3_c_RNIKE1T_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25034\,
            in2 => \N__21256\,
            in3 => \N__21194\,
            lcout => \pid_alt.error_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_3\,
            carryout => \pid_alt.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_4_c_RNINI2T_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21191\,
            in2 => \N__21185\,
            in3 => \N__21128\,
            lcout => \pid_alt.error_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_4\,
            carryout => \pid_alt.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_5_c_RNIQM3T_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21125\,
            in2 => \N__21901\,
            in3 => \N__21842\,
            lcout => \pid_alt.error_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_5\,
            carryout => \pid_alt.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_6_c_RNITQ4T_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21839\,
            in2 => \N__21832\,
            in3 => \N__21785\,
            lcout => \pid_alt.error_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_6\,
            carryout => \pid_alt.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_7_c_RNI9LEM_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21782\,
            in2 => \N__21776\,
            in3 => \N__21719\,
            lcout => \pid_alt.error_8\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \pid_alt.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_8_c_RNICPFM_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21716\,
            in2 => \N__21710\,
            in3 => \N__21653\,
            lcout => \pid_alt.error_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_8\,
            carryout => \pid_alt.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_9_c_RNIMMUJ_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21650\,
            in2 => \N__21644\,
            in3 => \N__21587\,
            lcout => \pid_alt.error_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_9\,
            carryout => \pid_alt.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_10_c_RNI0SDO_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22001\,
            in2 => \N__21584\,
            in3 => \N__21530\,
            lcout => \pid_alt.error_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_10\,
            carryout => \pid_alt.error_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_11_c_RNI5JAH_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23129\,
            in3 => \N__21482\,
            lcout => \pid_alt.error_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_11\,
            carryout => \pid_alt.error_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_12_c_RNI7MBH_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23057\,
            in2 => \_gnd_net_\,
            in3 => \N__21434\,
            lcout => \pid_alt.error_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_12\,
            carryout => \pid_alt.error_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_13_c_RNI9PCH_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23045\,
            in2 => \_gnd_net_\,
            in3 => \N__22049\,
            lcout => \pid_alt.error_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_13\,
            carryout => \pid_alt.error_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_14_c_RNIBSDH_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22046\,
            in2 => \_gnd_net_\,
            in3 => \N__22040\,
            lcout => \pid_alt.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22007\,
            lcout => drone_altitude_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_11_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__23747\,
            in1 => \N__31988\,
            in2 => \N__21995\,
            in3 => \N__22660\,
            lcout => \pid_alt.error_i_acummZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51377\,
            ce => 'H',
            sr => \N__33227\
        );

    \pid_alt.error_i_acumm_7_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__21970\,
            in2 => \N__22664\,
            in3 => \N__24043\,
            lcout => \pid_alt.error_i_acummZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51377\,
            ce => 'H',
            sr => \N__33227\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39652\,
            in2 => \_gnd_net_\,
            in3 => \N__50803\,
            lcout => alt_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51362\,
            ce => \N__25948\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_6_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40010\,
            lcout => alt_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51362\,
            ce => \N__25948\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIRSI31_11_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__23534\,
            in1 => \N__27612\,
            in2 => \_gnd_net_\,
            in3 => \N__49772\,
            lcout => \Commands_frame_decoder.state_RNIRSI31Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_1_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39761\,
            in2 => \_gnd_net_\,
            in3 => \N__40001\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23545\,
            in1 => \N__39483\,
            in2 => \N__22136\,
            in3 => \N__40261\,
            lcout => \Commands_frame_decoder.state_ns_0_a3_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__26901\,
            in2 => \N__22133\,
            in3 => \N__27440\,
            lcout => \Commands_frame_decoder.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51524\,
            ce => 'H',
            sr => \N__49504\
        );

    \Commands_frame_decoder.state_RNI6QPK_14_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27265\,
            in2 => \_gnd_net_\,
            in3 => \N__23650\,
            lcout => \Commands_frame_decoder.N_382_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_ess_7_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39983\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51514\,
            ce => \N__25318\,
            sr => \N__49509\
        );

    \Commands_frame_decoder.source_CH4data_esr_5_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40246\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51514\,
            ce => \N__25318\,
            sr => \N__49509\
        );

    \pid_alt.state_1_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.N_72_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51507\,
            ce => 'H',
            sr => \N__49512\
        );

    \Commands_frame_decoder.state_5_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__23612\,
            in1 => \N__25451\,
            in2 => \_gnd_net_\,
            in3 => \N__26903\,
            lcout => \Commands_frame_decoder.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51507\,
            ce => 'H',
            sr => \N__49512\
        );

    \pid_alt.error_d_reg_prev_esr_RNIFBF74_12_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22228\,
            in1 => \N__22124\,
            in2 => \N__22708\,
            in3 => \N__22114\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIFBF74Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_12_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__22219\,
            in1 => \N__23989\,
            in2 => \_gnd_net_\,
            in3 => \N__23592\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHMZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISAO32_12_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__22229\,
            in1 => \_gnd_net_\,
            in2 => \N__22118\,
            in3 => \N__22115\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISAO32Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIMJHM_0_13_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__22300\,
            in1 => \N__22277\,
            in2 => \_gnd_net_\,
            in3 => \N__22257\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIMJHM_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJ0N32_11_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22199\,
            in1 => \N__23774\,
            in2 => \_gnd_net_\,
            in3 => \N__24220\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJ0N32Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJGHM_0_12_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__23593\,
            in1 => \_gnd_net_\,
            in2 => \N__23993\,
            in3 => \N__22220\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIJGHM_0Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIKFGA4_11_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__23845\,
            in1 => \N__23773\,
            in2 => \N__22193\,
            in3 => \N__24219\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIKFGA4Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_14_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__22426\,
            in1 => \_gnd_net_\,
            in2 => \N__22406\,
            in3 => \N__22157\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIPMHMZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIOOO02_14_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22171\,
            in2 => \N__22178\,
            in3 => \N__24127\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIOOO02Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_0_15_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__28624\,
            in1 => \_gnd_net_\,
            in2 => \N__28612\,
            in3 => \N__28572\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHM_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIPMHM_0_14_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__22156\,
            in1 => \N__22402\,
            in2 => \_gnd_net_\,
            in3 => \N__22425\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIPMHM_0Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNICQF44_13_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22393\,
            in1 => \N__23020\,
            in2 => \N__22430\,
            in3 => \N__24150\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNICQF44Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_14_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22427\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51486\,
            ce => \N__25558\,
            sr => \N__49519\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGFN02_13_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__22394\,
            in1 => \N__22379\,
            in2 => \_gnd_net_\,
            in3 => \N__24151\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGFN02Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_5_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__22316\,
            in1 => \N__22330\,
            in2 => \N__22343\,
            in3 => \N__22628\,
            lcout => \pid_alt.error_i_acummZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI175B_12_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__33336\,
            in1 => \N__33314\,
            in2 => \N__33393\,
            in3 => \N__24099\,
            lcout => \pid_alt.N_295\,
            ltout => \pid_alt.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_1_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22676\,
            in2 => \N__22364\,
            in3 => \N__24056\,
            lcout => \pid_alt.error_i_acummZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.error_i_acumm_esr_2_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__22630\,
            in1 => \_gnd_net_\,
            in2 => \N__22682\,
            in3 => \N__24011\,
            lcout => \pid_alt.error_i_acummZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.error_i_acumm_esr_3_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24071\,
            in1 => \N__22631\,
            in2 => \_gnd_net_\,
            in3 => \N__22680\,
            lcout => \pid_alt.error_i_acummZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIP4VR2_4_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__22603\,
            in1 => \N__22339\,
            in2 => \N__22331\,
            in3 => \N__22315\,
            lcout => \pid_alt.N_294\,
            ltout => \pid_alt.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22629\,
            in2 => \N__22685\,
            in3 => \N__24977\,
            lcout => \pid_alt.error_i_acummZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.error_i_acumm_esr_4_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__22681\,
            in1 => \_gnd_net_\,
            in2 => \N__22647\,
            in3 => \N__22604\,
            lcout => \pid_alt.error_i_acummZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51474\,
            ce => \N__33256\,
            sr => \N__33197\
        );

    \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23185\,
            in2 => \N__23189\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_0_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22567\,
            in2 => \N__22556\,
            in3 => \N__22541\,
            lcout => \pid_alt.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_0\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_1_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22538\,
            in2 => \N__24199\,
            in3 => \N__22526\,
            lcout => \pid_alt.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_0\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_1\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_2_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22523\,
            in2 => \N__24177\,
            in3 => \N__22511\,
            lcout => \pid_alt.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_1\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_2\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_3_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22508\,
            in2 => \N__24246\,
            in3 => \N__22496\,
            lcout => \pid_alt.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_2\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_3\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_4_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22489\,
            in2 => \N__22472\,
            in3 => \N__22460\,
            lcout => \pid_alt.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_3\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_4\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_5_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22457\,
            in2 => \N__22448\,
            in3 => \N__22829\,
            lcout => \pid_alt.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_4\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_5\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_6_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22826\,
            in2 => \N__22813\,
            in3 => \N__22784\,
            lcout => \pid_alt.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_5\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_6\,
            clk => \N__51462\,
            ce => \N__25562\,
            sr => \N__49531\
        );

    \pid_alt.pid_prereg_esr_7_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24530\,
            in2 => \N__24575\,
            in3 => \N__22781\,
            lcout => \pid_alt.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_7\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_8_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24395\,
            in2 => \N__24670\,
            in3 => \N__22778\,
            lcout => \pid_alt.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_7\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_8\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_9_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22775\,
            in2 => \N__24358\,
            in3 => \N__22766\,
            lcout => \pid_alt.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_8\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_9\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_10_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22763\,
            in2 => \N__22757\,
            in3 => \N__22739\,
            lcout => \pid_alt.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_9\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_10\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_11_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23954\,
            in2 => \N__23977\,
            in3 => \N__22736\,
            lcout => \pid_alt.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_10\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_11\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_12_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22733\,
            in2 => \N__23852\,
            in3 => \N__22724\,
            lcout => \pid_alt.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_11\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_12\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_13_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22721\,
            in2 => \N__22712\,
            in3 => \N__22688\,
            lcout => \pid_alt.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_12\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_13\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_14_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23021\,
            in2 => \N__23006\,
            in3 => \N__22994\,
            lcout => \pid_alt.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_13\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_14\,
            clk => \N__51445\,
            ce => \N__25566\,
            sr => \N__49539\
        );

    \pid_alt.pid_prereg_esr_15_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22991\,
            in2 => \N__22981\,
            in3 => \N__22955\,
            lcout => \pid_alt.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_15\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_16_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22952\,
            in2 => \N__22946\,
            in3 => \N__22925\,
            lcout => \pid_alt.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_15\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_16\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_17_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22922\,
            in2 => \N__22915\,
            in3 => \N__22898\,
            lcout => \pid_alt.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_16\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_17\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_18_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22895\,
            in2 => \N__22886\,
            in3 => \N__22871\,
            lcout => \pid_alt.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_17\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_18\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_19_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22868\,
            in2 => \N__22859\,
            in3 => \N__22838\,
            lcout => \pid_alt.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_18\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_19\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_20_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24926\,
            in2 => \N__24949\,
            in3 => \N__22835\,
            lcout => \pid_alt.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_19\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_20\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_21_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24695\,
            in2 => \N__24815\,
            in3 => \N__22832\,
            lcout => \pid_alt.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_20\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_21\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_22_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23120\,
            in2 => \N__23105\,
            in3 => \N__23108\,
            lcout => \pid_alt.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_21\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_22\,
            clk => \N__51431\,
            ce => \N__25567\,
            sr => \N__49546\
        );

    \pid_alt.pid_prereg_esr_23_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23104\,
            in2 => \N__23078\,
            in3 => \N__23063\,
            lcout => \pid_alt.pid_preregZ0Z_23\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_23\,
            clk => \N__51418\,
            ce => \N__25571\,
            sr => \N__49552\
        );

    \pid_alt.pid_prereg_esr_24_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000101111110"
        )
    port map (
            in0 => \N__24754\,
            in1 => \N__24727\,
            in2 => \N__24800\,
            in3 => \N__23060\,
            lcout => \pid_alt.pid_preregZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51418\,
            ce => \N__25571\,
            sr => \N__49552\
        );

    \pid_alt.error_axb_13_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23051\,
            lcout => \pid_alt.error_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_13_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36879\,
            lcout => drone_altitude_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51403\,
            ce => \N__25819\,
            sr => \N__49562\
        );

    \pid_alt.error_axb_14_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23039\,
            lcout => \pid_alt.error_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48435\,
            lcout => drone_altitude_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51403\,
            ce => \N__25819\,
            sr => \N__49562\
        );

    \pid_alt.error_axb_2_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24683\,
            lcout => \pid_alt.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_3_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24677\,
            lcout => \pid_alt.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI2Q08_0_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23681\,
            lcout => \pid_alt.error_d_reg_prev_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIKAP4_8_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23162\,
            lcout => \drone_H_disp_side_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_8_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42606\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51388\,
            ce => \N__29587\,
            sr => \N__49569\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNILBP4_9_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23156\,
            lcout => \drone_H_disp_side_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_9_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36807\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51388\,
            ce => \N__29587\,
            sr => \N__49569\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIT4RD_10_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23150\,
            lcout => \drone_H_disp_side_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_10_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37128\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51388\,
            ce => \N__29587\,
            sr => \N__49569\
        );

    \pid_alt.error_axb_1_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24689\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_12_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \pid_alt.error_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_0_c_inv_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23321\,
            in2 => \_gnd_net_\,
            in3 => \N__27154\,
            lcout => \pid_side.error_axb_0\,
            ltout => OPEN,
            carryin => \bfn_4_21_0_\,
            carryout => \pid_side.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_0_c_RNI43F5_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28466\,
            in2 => \_gnd_net_\,
            in3 => \N__23300\,
            lcout => \pid_side.error_1\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_0\,
            carryout => \pid_side.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_1_c_RNI66G5_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25991\,
            in2 => \_gnd_net_\,
            in3 => \N__23285\,
            lcout => \pid_side.error_2\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_1\,
            carryout => \pid_side.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_2_c_RNI89H5_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25982\,
            in2 => \_gnd_net_\,
            in3 => \N__23267\,
            lcout => \pid_side.error_3\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_2\,
            carryout => \pid_side.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_3_c_RNI1SDJ_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25223\,
            in2 => \N__25766\,
            in3 => \N__23252\,
            lcout => \pid_side.error_4\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_3\,
            carryout => \pid_side.error_cry_0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_0_0_c_RNIF3ET_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25214\,
            in2 => \N__25742\,
            in3 => \N__23237\,
            lcout => \pid_side.error_5\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_0_0\,
            carryout => \pid_side.error_cry_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_1_0_c_RNII9K11_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25229\,
            in2 => \N__25208\,
            in3 => \N__23219\,
            lcout => \pid_side.error_6\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_1_0\,
            carryout => \pid_side.error_cry_2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_2_0_c_RNILFQL_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25199\,
            in2 => \N__25754\,
            in3 => \N__23201\,
            lcout => \pid_side.error_7\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_2_0\,
            carryout => \pid_side.error_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_3_0_c_RNIOL0Q_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23198\,
            in2 => \N__25193\,
            in3 => \N__23480\,
            lcout => \pid_side.error_8\,
            ltout => OPEN,
            carryin => \bfn_4_22_0_\,
            carryout => \pid_side.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_4_c_RNIC8FJ_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23477\,
            in2 => \N__25184\,
            in3 => \N__23453\,
            lcout => \pid_side.error_9\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_4\,
            carryout => \pid_side.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_5_c_RNIM4IS_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25175\,
            in2 => \N__23450\,
            in3 => \N__23423\,
            lcout => \pid_side.error_10\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_5\,
            carryout => \pid_side.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_6_c_RNIQBMT_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28493\,
            in2 => \_gnd_net_\,
            in3 => \N__23405\,
            lcout => \pid_side.error_11\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_6\,
            carryout => \pid_side.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_7_c_RNIPRDP1_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28520\,
            in2 => \N__29549\,
            in3 => \N__23387\,
            lcout => \pid_side.error_12\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_7\,
            carryout => \pid_side.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_8_c_RNIUUKS_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29636\,
            in2 => \N__29522\,
            in3 => \N__23369\,
            lcout => \pid_side.error_13\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_8\,
            carryout => \pid_side.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_9_c_RNI13MS_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24956\,
            in2 => \N__29612\,
            in3 => \N__23351\,
            lcout => \pid_side.error_14\,
            ltout => OPEN,
            carryin => \pid_side.error_cry_9\,
            carryout => \pid_side.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_cry_10_c_RNIBCT11_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__25169\,
            in1 => \N__29611\,
            in2 => \_gnd_net_\,
            in3 => \N__23348\,
            lcout => \pid_side.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_0_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39768\,
            in2 => \_gnd_net_\,
            in3 => \N__50802\,
            lcout => alt_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51352\,
            ce => \N__25947\,
            sr => \_gnd_net_\
        );

    \pid_alt.state_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31147\,
            in1 => \N__32842\,
            in2 => \_gnd_net_\,
            in3 => \N__32022\,
            lcout => \pid_alt.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51529\,
            ce => 'H',
            sr => \N__49498\
        );

    \Commands_frame_decoder.state_12_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23533\,
            in1 => \N__27609\,
            in2 => \N__25306\,
            in3 => \N__26913\,
            lcout => \Commands_frame_decoder.stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51525\,
            ce => 'H',
            sr => \N__49500\
        );

    \Commands_frame_decoder.state_RNO_1_0_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__23560\,
            in1 => \N__27438\,
            in2 => \N__23669\,
            in3 => \N__23570\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_0_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__23546\,
            in1 => \N__23561\,
            in2 => \N__23552\,
            in3 => \N__25352\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__26880\,
            in1 => \N__23656\,
            in2 => \N__23549\,
            in3 => \N__25340\,
            lcout => \Commands_frame_decoder.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51520\,
            ce => 'H',
            sr => \N__49502\
        );

    \Commands_frame_decoder.state_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__27439\,
            in1 => \N__23621\,
            in2 => \N__25429\,
            in3 => \N__26879\,
            lcout => \Commands_frame_decoder.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51520\,
            ce => 'H',
            sr => \N__49502\
        );

    \Commands_frame_decoder.preinit_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25251\,
            in2 => \_gnd_net_\,
            in3 => \N__27607\,
            lcout => \Commands_frame_decoder.preinitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51515\,
            ce => 'H',
            sr => \N__49505\
        );

    \Commands_frame_decoder.state_11_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27606\,
            in1 => \N__23529\,
            in2 => \N__26825\,
            in3 => \N__26902\,
            lcout => \Commands_frame_decoder.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51515\,
            ce => 'H',
            sr => \N__49505\
        );

    \scaler_4.N_1684_i_l_ofx_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25394\,
            in2 => \_gnd_net_\,
            in3 => \N__23510\,
            lcout => \scaler_4.N_1684_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_3_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39697\,
            in1 => \N__39974\,
            in2 => \N__39467\,
            in3 => \N__40238\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_2_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__39975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39698\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_2_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__39439\,
            in1 => \N__23657\,
            in2 => \N__23624\,
            in3 => \N__40239\,
            lcout => \Commands_frame_decoder.state_ns_0_a3_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_2_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28769\,
            in1 => \N__27421\,
            in2 => \N__39474\,
            in3 => \N__28874\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIHL1J_5_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23611\,
            in2 => \_gnd_net_\,
            in3 => \N__27568\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIE28S_5_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23600\,
            in3 => \N__49750\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28775\,
            in1 => \N__27420\,
            in2 => \N__27344\,
            in3 => \N__39706\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIQRI31_10_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__27567\,
            in1 => \N__26818\,
            in2 => \_gnd_net_\,
            in3 => \N__49749\,
            lcout => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_15_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28576\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51487\,
            ce => \N__25554\,
            sr => \N__49513\
        );

    \pid_alt.error_d_reg_prev_esr_12_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23597\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51487\,
            ce => \N__25554\,
            sr => \N__49513\
        );

    \pid_alt.error_d_reg_prev_esr_RNITPKD4_10_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23830\,
            in1 => \N__23861\,
            in2 => \N__23981\,
            in3 => \N__23763\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNITPKD4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIDAHM_10_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__23942\,
            in1 => \N__23915\,
            in2 => \_gnd_net_\,
            in3 => \N__23891\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIDAHMZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI1FP62_10_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__23831\,
            in1 => \_gnd_net_\,
            in2 => \N__23855\,
            in3 => \N__23764\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI1FP62Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGDHM_0_11_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__23788\,
            in1 => \N__23797\,
            in2 => \_gnd_net_\,
            in3 => \N__23820\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGDHM_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_11_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23822\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51475\,
            ce => \N__25555\,
            sr => \N__49516\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGDHM_11_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001010"
        )
    port map (
            in0 => \N__23821\,
            in1 => \_gnd_net_\,
            in2 => \N__23801\,
            in3 => \N__23789\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGDHMZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_11_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23765\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51475\,
            ce => \N__25555\,
            sr => \N__49516\
        );

    \pid_alt.error_d_reg_prev_esr_0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23717\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_3_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24247\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_12_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24224\,
            lcout => \pid_alt.error_i_acumm7lto12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_1_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24200\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_2_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24178\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_14_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24155\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_prereg_esr_15_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24131\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51463\,
            ce => \N__25559\,
            sr => \N__49520\
        );

    \pid_alt.error_i_acumm_esr_12_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__33319\,
            in1 => \N__33395\,
            in2 => \N__33346\,
            in3 => \N__24100\,
            lcout => \pid_alt.error_i_acummZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51446\,
            ce => \N__33255\,
            sr => \N__33196\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIRFAQ1_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24067\,
            in1 => \N__24055\,
            in2 => \N__24044\,
            in3 => \N__24973\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_1_i_a5_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIE78O2_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33318\,
            in1 => \N__24007\,
            in2 => \N__23996\,
            in3 => \N__31968\,
            lcout => \pid_alt.un1_reset_1_i_a5_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIRRP7_14_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__24446\,
            in1 => \N__25730\,
            in2 => \N__25616\,
            in3 => \N__24440\,
            lcout => \pid_alt.N_557\,
            ltout => \pid_alt.N_557_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIVV9C5_10_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24434\,
            in1 => \N__24422\,
            in2 => \N__24410\,
            in3 => \N__24407\,
            lcout => OPEN,
            ltout => \pid_alt.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI8HS46_21_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__31969\,
            in1 => \N__33394\,
            in2 => \N__24401\,
            in3 => \N__49042\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21\,
            ltout => \pid_alt.error_i_acumm_prereg_esr_RNI8HS46Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIT64J6_1_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24398\,
            in3 => \N__31970\,
            lcout => \pid_alt.N_72_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI5G6Q5_7_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24262\,
            in1 => \N__24389\,
            in2 => \N__24671\,
            in3 => \N__24379\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI5G6Q5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_7_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24616\,
            in1 => \N__24625\,
            in2 => \_gnd_net_\,
            in3 => \N__24651\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIF2611Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI7T3T2_7_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__24263\,
            in1 => \_gnd_net_\,
            in2 => \N__24383\,
            in3 => \N__24380\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI7T3T2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNII5611_0_8_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24341\,
            in1 => \N__24317\,
            in2 => \_gnd_net_\,
            in3 => \N__24296\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNII5611_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_7_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51432\,
            ce => \N__25563\,
            sr => \N__49532\
        );

    \pid_alt.error_d_reg_prev_esr_RNIUI2T2_6_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__24590\,
            in1 => \_gnd_net_\,
            in2 => \N__24599\,
            in3 => \N__24551\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIUI2T2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIF2611_0_7_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__24652\,
            in1 => \_gnd_net_\,
            in2 => \N__24629\,
            in3 => \N__24617\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIF2611_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIJR3Q5_6_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__24589\,
            in1 => \N__24574\,
            in2 => \N__24554\,
            in3 => \N__24550\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIJR3Q5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNICSUM_17_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24524\,
            in1 => \N__24518\,
            in2 => \N__24512\,
            in3 => \N__24503\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIBRUM_15_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24497\,
            in1 => \N__24491\,
            in2 => \N__24485\,
            in3 => \N__24476\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_20_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__24862\,
            in1 => \N__24871\,
            in2 => \_gnd_net_\,
            in3 => \N__24843\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIGGKMZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNI86IM_19_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__24919\,
            in1 => \N__24470\,
            in2 => \_gnd_net_\,
            in3 => \N__24886\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNI86IMZ0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIK3024_19_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__24950\,
            in1 => \N__24785\,
            in2 => \N__24929\,
            in3 => \N__25635\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIK3024Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_19_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24920\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51404\,
            ce => \N__25568\,
            sr => \N__49547\
        );

    \pid_alt.error_d_reg_prev_esr_20_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24844\,
            lcout => \pid_alt.error_d_reg_prevZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51404\,
            ce => \N__25568\,
            sr => \N__49547\
        );

    \pid_alt.error_d_reg_prev_esr_RNIGGKM_0_20_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__24872\,
            in1 => \N__24863\,
            in2 => \_gnd_net_\,
            in3 => \N__24845\,
            lcout => \pid_alt.un1_pid_prereg_236_1\,
            ltout => \pid_alt.un1_pid_prereg_236_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIS5212_19_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24824\,
            in2 => \N__24818\,
            in3 => \N__25636\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19\,
            ltout => \pid_alt.error_d_reg_prev_esr_RNIS5212Z0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_d_reg_prev_esr_RNIO6034_20_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24786\,
            in1 => \N__24750\,
            in2 => \N__24734\,
            in3 => \N__24726\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNIO6034Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_1_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36796\,
            lcout => drone_altitude_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \dron_frame_decoder_1.source_Altitude_esr_2_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37118\,
            lcout => drone_altitude_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \dron_frame_decoder_1.source_Altitude_esr_3_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37044\,
            lcout => drone_altitude_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36969\,
            lcout => \dron_frame_decoder_1.drone_altitude_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \dron_frame_decoder_1.source_Altitude_esr_5_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36878\,
            lcout => \dron_frame_decoder_1.drone_altitude_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48434\,
            lcout => \dron_frame_decoder_1.drone_altitude_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51389\,
            ce => \N__33470\,
            sr => \N__49553\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_0_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39755\,
            in2 => \_gnd_net_\,
            in3 => \N__50809\,
            lcout => xy_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51378\,
            ce => \N__39026\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_2_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39525\,
            in2 => \_gnd_net_\,
            in3 => \N__50810\,
            lcout => xy_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51378\,
            ce => \N__39026\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_5_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40093\,
            lcout => xy_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51378\,
            ce => \N__39026\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25040\,
            lcout => drone_altitude_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_0_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25022\,
            in2 => \_gnd_net_\,
            in3 => \N__24998\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51363\,
            ce => \N__25574\,
            sr => \N__49570\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNI08RD_13_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29632\,
            lcout => \drone_H_disp_side_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNII8P4_6_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27113\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_side_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_0_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39759\,
            lcout => side_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_1_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39653\,
            lcout => side_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_2_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39526\,
            lcout => side_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_3_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39366\,
            lcout => side_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_4_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40402\,
            lcout => side_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_5_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40274\,
            lcout => side_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \Commands_frame_decoder.source_CH2data_esr_6_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40121\,
            lcout => side_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51353\,
            ce => \N__27047\,
            sr => \N__49580\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_15_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36627\,
            lcout => \drone_H_disp_side_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51343\,
            ce => \N__29591\,
            sr => \N__49589\
        );

    \Commands_frame_decoder.source_data_valid_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__26090\,
            in1 => \N__25262\,
            in2 => \N__27186\,
            in3 => \N__27614\,
            lcout => \debug_CH3_20A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51521\,
            ce => 'H',
            sr => \N__49499\
        );

    \Commands_frame_decoder.state_13_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__25286\,
            in2 => \N__25307\,
            in3 => \N__26851\,
            lcout => \Commands_frame_decoder.stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51516\,
            ce => 'H',
            sr => \N__49501\
        );

    \Commands_frame_decoder.state_14_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__25285\,
            in1 => \N__27598\,
            in2 => \_gnd_net_\,
            in3 => \N__25336\,
            lcout => \Commands_frame_decoder.stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51516\,
            ce => 'H',
            sr => \N__49501\
        );

    \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__26178\,
            in1 => \N__26196\,
            in2 => \N__26162\,
            in3 => \N__26212\,
            lcout => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNII19A1_4_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26245\,
            in1 => \N__26020\,
            in2 => \N__26231\,
            in3 => \N__26035\,
            lcout => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNID7P31_6_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__26179\,
            in1 => \N__26005\,
            in2 => \_gnd_net_\,
            in3 => \N__26197\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__26260\,
            in1 => \N__25277\,
            in2 => \N__25271\,
            in3 => \N__25268\,
            lcout => \Commands_frame_decoder.WDT8lt14_0\,
            ltout => \Commands_frame_decoder.WDT8lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIF92K5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__26141\,
            in1 => \N__25261\,
            in2 => \N__25232\,
            in3 => \N__26115\,
            lcout => \Commands_frame_decoder.state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__25361\,
            in1 => \N__26143\,
            in2 => \N__27608\,
            in3 => \N__26116\,
            lcout => \Commands_frame_decoder.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__26142\,
            in1 => \N__27577\,
            in2 => \N__26120\,
            in3 => \N__25360\,
            lcout => \Commands_frame_decoder.N_377_0\,
            ltout => \Commands_frame_decoder.N_377_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNIA5DM6_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__27254\,
            in1 => \N__27230\,
            in2 => \N__25343\,
            in3 => \N__27578\,
            lcout => \Commands_frame_decoder.N_384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH4data_esr_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39754\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_CH4data_esr_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39577\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_CH4data_esr_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_CH4data_esr_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39344\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_CH4data_esr_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40359\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_CH4data_esr_6_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40106\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51498\,
            ce => \N__25325\,
            sr => \N__49506\
        );

    \Commands_frame_decoder.source_offset4data_esr_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39753\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_esr_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39594\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_esr_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39466\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39343\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_esr_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40378\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_esr_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40254\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.source_offset4data_ess_7_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39982\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51488\,
            ce => \N__26956\,
            sr => \N__49508\
        );

    \Commands_frame_decoder.state_6_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__25379\,
            in1 => \N__26702\,
            in2 => \_gnd_net_\,
            in3 => \N__26894\,
            lcout => \Commands_frame_decoder.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51476\,
            ce => 'H',
            sr => \N__49510\
        );

    \uart_pc.data_rdy_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40704\,
            in2 => \_gnd_net_\,
            in3 => \N__28799\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51476\,
            ce => 'H',
            sr => \N__49510\
        );

    \Commands_frame_decoder.state_RNIGK1J_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25369\,
            in2 => \_gnd_net_\,
            in3 => \N__27491\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_4_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__25370\,
            in1 => \N__25786\,
            in2 => \_gnd_net_\,
            in3 => \N__26893\,
            lcout => \Commands_frame_decoder.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51476\,
            ce => 'H',
            sr => \N__49510\
        );

    \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__26676\,
            in1 => \N__26493\,
            in2 => \_gnd_net_\,
            in3 => \N__26569\,
            lcout => \dron_frame_decoder_1.WDT10lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26524\,
            in1 => \N__26584\,
            in2 => \N__26603\,
            in3 => \N__26539\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__26554\,
            in1 => \N__25457\,
            in2 => \N__25469\,
            in3 => \N__25466\,
            lcout => \dron_frame_decoder_1.WDT10lt14_0\,
            ltout => \dron_frame_decoder_1.WDT10lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27780\,
            in2 => \N__25460\,
            in3 => \N__27801\,
            lcout => \dron_frame_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__26494\,
            in1 => \N__26509\,
            in2 => \N__26660\,
            in3 => \N__26677\,
            lcout => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNID18S_4_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25450\,
            in2 => \_gnd_net_\,
            in3 => \N__49748\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_6_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28774\,
            in1 => \N__27422\,
            in2 => \N__40562\,
            in3 => \N__39930\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51447\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25405\,
            in2 => \_gnd_net_\,
            in3 => \N__27536\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIEI1J_2_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \_gnd_net_\,
            in3 => \N__27537\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0\,
            ltout => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25406\,
            in2 => \N__25409\,
            in3 => \N__26914\,
            lcout => \Commands_frame_decoder.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51433\,
            ce => 'H',
            sr => \N__49521\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIIDE4_16_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25670\,
            in1 => \N__25646\,
            in2 => \N__25700\,
            in3 => \N__25583\,
            lcout => \pid_alt.m7_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_19_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25721\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51419\,
            ce => \N__25556\,
            sr => \N__49524\
        );

    \pid_alt.pid_prereg_esr_RNI046H1_1_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30590\,
            in1 => \N__31483\,
            in2 => \N__30648\,
            in3 => \N__31516\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_i_a5_1_10_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIJF5N2_10_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30547\,
            in1 => \N__30298\,
            in2 => \N__25691\,
            in3 => \N__29140\,
            lcout => \pid_alt.un1_reset_i_a5_1_10_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_18_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25688\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51405\,
            ce => \N__25560\,
            sr => \N__49533\
        );

    \pid_alt.error_i_acumm_prereg_esr_17_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25664\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51405\,
            ce => \N__25560\,
            sr => \N__49533\
        );

    \pid_alt.error_i_acumm_prereg_esr_20_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25640\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51405\,
            ce => \N__25560\,
            sr => \N__49533\
        );

    \pid_alt.error_i_acumm_prereg_esr_16_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25601\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51405\,
            ce => \N__25560\,
            sr => \N__49533\
        );

    \Commands_frame_decoder.state_RNIBV7S_2_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25486\,
            in2 => \_gnd_net_\,
            in3 => \N__49767\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIT4CP1_14_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__25865\,
            in1 => \N__25853\,
            in2 => \N__25844\,
            in3 => \N__25832\,
            lcout => \pid_alt.N_551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIFCSD1_0_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__32841\,
            in1 => \N__31986\,
            in2 => \N__31178\,
            in3 => \N__49747\,
            lcout => \pid_alt.state_RNIFCSD1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26780\,
            in2 => \_gnd_net_\,
            in3 => \N__49033\,
            lcout => \dron_frame_decoder_1.N_755_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_7_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36616\,
            lcout => \dron_frame_decoder_1.drone_altitude_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51364\,
            ce => \N__33462\,
            sr => \N__49554\
        );

    \Commands_frame_decoder.state_RNIC08S_3_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25787\,
            in2 => \_gnd_net_\,
            in3 => \N__49768\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI36DT_4_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28097\,
            in2 => \_gnd_net_\,
            in3 => \N__49773\,
            lcout => \dron_frame_decoder_1.N_747_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIG6P4_4_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27125\,
            lcout => \drone_H_disp_side_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIJ9P4_7_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27104\,
            lcout => \drone_H_disp_side_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIH7P4_5_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27119\,
            lcout => \drone_H_disp_side_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_axb_2_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27137\,
            lcout => \pid_side.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_axb_3_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27131\,
            lcout => \pid_side.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_4_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__25966\,
            in1 => \N__27611\,
            in2 => \N__26719\,
            in3 => \N__40401\,
            lcout => alt_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51336\,
            ce => 'H',
            sr => \N__49581\
        );

    \Commands_frame_decoder.state_RNIF38S_6_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__26712\,
            in1 => \N__27610\,
            in2 => \_gnd_net_\,
            in3 => \N__49771\,
            lcout => \Commands_frame_decoder.state_RNIF38SZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNICP2N1_0_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25922\,
            in2 => \_gnd_net_\,
            in3 => \N__50795\,
            lcout => \pid_alt.N_850_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25892\,
            lcout => \uart_drone_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_0__0__0_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25898\,
            lcout => \uart_drone_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51536\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_2__0__0_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25886\,
            lcout => \uart_drone_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_ctle_14_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27176\,
            in2 => \_gnd_net_\,
            in3 => \N__49752\,
            lcout => \scaler_4.debug_CH3_20A_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_data_valid_RNO_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27219\,
            in2 => \_gnd_net_\,
            in3 => \N__27255\,
            lcout => \Commands_frame_decoder.count_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26069\,
            in2 => \N__26084\,
            in3 => \N__26083\,
            lcout => \Commands_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_0\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26063\,
            in2 => \_gnd_net_\,
            in3 => \N__26057\,
            lcout => \Commands_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_0\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_1\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26054\,
            in2 => \_gnd_net_\,
            in3 => \N__26048\,
            lcout => \Commands_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_1\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_2\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26045\,
            in2 => \_gnd_net_\,
            in3 => \N__26039\,
            lcout => \Commands_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_2\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_3\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26036\,
            in2 => \_gnd_net_\,
            in3 => \N__26024\,
            lcout => \Commands_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_3\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_4\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26021\,
            in2 => \_gnd_net_\,
            in3 => \N__26009\,
            lcout => \Commands_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_4\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_5\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26006\,
            in2 => \_gnd_net_\,
            in3 => \N__25994\,
            lcout => \Commands_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_5\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_6\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_7_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26261\,
            in2 => \_gnd_net_\,
            in3 => \N__26249\,
            lcout => \Commands_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_6\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_7\,
            clk => \N__51509\,
            ce => 'H',
            sr => \N__26462\
        );

    \Commands_frame_decoder.WDT_8_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26246\,
            in2 => \_gnd_net_\,
            in3 => \N__26234\,
            lcout => \Commands_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_8\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_9_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26230\,
            in2 => \_gnd_net_\,
            in3 => \N__26216\,
            lcout => \Commands_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_8\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_9\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26213\,
            in2 => \_gnd_net_\,
            in3 => \N__26201\,
            lcout => \Commands_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_9\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_10\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_11_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26198\,
            in2 => \_gnd_net_\,
            in3 => \N__26183\,
            lcout => \Commands_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_10\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_11\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_12_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26180\,
            in2 => \_gnd_net_\,
            in3 => \N__26165\,
            lcout => \Commands_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_11\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_12\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_13_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26161\,
            in2 => \_gnd_net_\,
            in3 => \N__26147\,
            lcout => \Commands_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_12\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_13\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_14_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26144\,
            in2 => \_gnd_net_\,
            in3 => \N__26126\,
            lcout => \Commands_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_13\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_14\,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \Commands_frame_decoder.WDT_15_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26114\,
            in2 => \_gnd_net_\,
            in3 => \N__26123\,
            lcout => \Commands_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51499\,
            ce => 'H',
            sr => \N__26458\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28937\,
            in2 => \N__28974\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26399\,
            in2 => \N__26393\,
            in3 => \N__26384\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26381\,
            in2 => \N__26375\,
            in3 => \N__26366\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26363\,
            in2 => \N__26357\,
            in3 => \N__26348\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26345\,
            in2 => \N__26339\,
            in3 => \N__26330\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26327\,
            in2 => \N__26315\,
            in3 => \N__26306\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26303\,
            in2 => \N__26297\,
            in3 => \N__26279\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26276\,
            in2 => \_gnd_net_\,
            in3 => \N__26264\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26477\,
            in2 => \N__48128\,
            in3 => \N__26468\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26465\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.un1_state57_i_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27535\,
            in2 => \_gnd_net_\,
            in3 => \N__49755\,
            lcout => \Commands_frame_decoder.un1_state57_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28756\,
            in1 => \N__27406\,
            in2 => \N__28856\,
            in3 => \N__39576\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__29007\,
            in1 => \N__28968\,
            in2 => \_gnd_net_\,
            in3 => \N__28938\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26423\,
            in2 => \N__26438\,
            in3 => \N__26437\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_0\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26417\,
            in2 => \_gnd_net_\,
            in3 => \N__26411\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_0\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_1\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26408\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_1\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_2\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26612\,
            in2 => \_gnd_net_\,
            in3 => \N__26606\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_2\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_3\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_4_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26602\,
            in2 => \_gnd_net_\,
            in3 => \N__26588\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_3\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_4\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26585\,
            in2 => \_gnd_net_\,
            in3 => \N__26573\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_4\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_5\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26570\,
            in2 => \_gnd_net_\,
            in3 => \N__26558\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_5\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_6\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_7_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26555\,
            in2 => \_gnd_net_\,
            in3 => \N__26543\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_6\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_7\,
            clk => \N__51464\,
            ce => 'H',
            sr => \N__26633\
        );

    \dron_frame_decoder_1.WDT_8_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26540\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_8\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_9_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26525\,
            in2 => \_gnd_net_\,
            in3 => \N__26513\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_8\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_9\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26510\,
            in2 => \_gnd_net_\,
            in3 => \N__26498\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_9\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_10\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_11_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26495\,
            in2 => \_gnd_net_\,
            in3 => \N__26480\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_10\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_11\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_12_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26678\,
            in2 => \_gnd_net_\,
            in3 => \N__26663\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_11\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_12\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_13_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26659\,
            in2 => \_gnd_net_\,
            in3 => \N__26645\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_12\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_13\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_14_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27784\,
            in2 => \_gnd_net_\,
            in3 => \N__26642\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_13\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_14\,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \dron_frame_decoder_1.WDT_15_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27803\,
            in2 => \_gnd_net_\,
            in3 => \N__26639\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51448\,
            ce => 'H',
            sr => \N__26623\
        );

    \uart_pc.data_1_4_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28773\,
            in1 => \N__27419\,
            in2 => \N__29081\,
            in3 => \N__40194\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36919\,
            in2 => \_gnd_net_\,
            in3 => \N__37009\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48426\,
            in1 => \N__27749\,
            in2 => \N__26636\,
            in3 => \N__36759\,
            lcout => \dron_frame_decoder_1.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29210\,
            in2 => \_gnd_net_\,
            in3 => \N__49759\,
            lcout => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0TLI1_4_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__28052\,
            in1 => \N__26765\,
            in2 => \N__49796\,
            in3 => \N__28120\,
            lcout => \dron_frame_decoder_1.N_763_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI3T3K1_7_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28051\,
            in1 => \N__26764\,
            in2 => \N__28078\,
            in3 => \N__28119\,
            lcout => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_rdy_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31054\,
            in2 => \_gnd_net_\,
            in3 => \N__29879\,
            lcout => uart_drone_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51420\,
            ce => 'H',
            sr => \N__49525\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_2_0_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29206\,
            in2 => \_gnd_net_\,
            in3 => \N__37112\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_2_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_2_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36609\,
            in1 => \N__36848\,
            in2 => \N__26768\,
            in3 => \N__42570\,
            lcout => \dron_frame_decoder_1.N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI7Q6K_5_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27998\,
            in2 => \_gnd_net_\,
            in3 => \N__29195\,
            lcout => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_2_0_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__28050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27752\,
            lcout => \dron_frame_decoder_1.state_ns_i_i_0_a2_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNITC181_2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__29239\,
            in1 => \N__29196\,
            in2 => \N__27839\,
            in3 => \N__49751\,
            lcout => \dron_frame_decoder_1.N_723_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_4_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__26745\,
            in1 => \N__27603\,
            in2 => \N__26998\,
            in3 => \N__40369\,
            lcout => xy_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51390\,
            ce => 'H',
            sr => \N__49540\
        );

    \Commands_frame_decoder.state_7_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27601\,
            in1 => \N__26991\,
            in2 => \N__26720\,
            in3 => \N__26916\,
            lcout => \Commands_frame_decoder.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51390\,
            ce => 'H',
            sr => \N__49540\
        );

    \Commands_frame_decoder.state_RNIG48S_7_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__26990\,
            in1 => \N__27600\,
            in2 => \_gnd_net_\,
            in3 => \N__49756\,
            lcout => \Commands_frame_decoder.state_RNIG48SZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_8_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27602\,
            in1 => \N__26974\,
            in2 => \N__26999\,
            in3 => \N__26917\,
            lcout => \Commands_frame_decoder.stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51390\,
            ce => 'H',
            sr => \N__49540\
        );

    \Commands_frame_decoder.state_9_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__26918\,
            in1 => \N__26936\,
            in2 => \N__26975\,
            in3 => \N__27604\,
            lcout => \Commands_frame_decoder.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51390\,
            ce => 'H',
            sr => \N__49540\
        );

    \Commands_frame_decoder.state_RNII68S_9_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__49757\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26927\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNILP1J_9_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26935\,
            in2 => \_gnd_net_\,
            in3 => \N__27599\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_10_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26811\,
            in2 => \N__26921\,
            in3 => \N__26915\,
            lcout => \Commands_frame_decoder.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51390\,
            ce => 'H',
            sr => \N__49540\
        );

    \pid_side.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49868\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34708\,
            in2 => \_gnd_net_\,
            in3 => \N__26789\,
            lcout => \pid_side.un1_pid_prereg_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_1\,
            carryout => \pid_side.un1_pid_prereg_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50107\,
            in2 => \_gnd_net_\,
            in3 => \N__26786\,
            lcout => \pid_side.un1_pid_prereg_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_2\,
            carryout => \pid_side.un1_pid_prereg_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28381\,
            in2 => \_gnd_net_\,
            in3 => \N__26783\,
            lcout => \pid_side.un1_pid_prereg_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_3\,
            carryout => \pid_side.un1_pid_prereg_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30865\,
            in2 => \N__48129\,
            in3 => \N__27026\,
            lcout => \pid_side.un1_pid_prereg_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_4\,
            carryout => \pid_side.un1_pid_prereg_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28348\,
            in2 => \N__48131\,
            in3 => \N__27023\,
            lcout => \pid_side.un1_pid_prereg_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_5\,
            carryout => \pid_side.un1_pid_prereg_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30361\,
            in2 => \N__48130\,
            in3 => \N__27020\,
            lcout => \pid_side.un1_pid_prereg_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_6\,
            carryout => \pid_side.un1_pid_prereg_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28450\,
            in2 => \N__48132\,
            in3 => \N__27017\,
            lcout => \pid_side.un1_pid_prereg_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_7\,
            carryout => \pid_side.un1_pid_prereg_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48136\,
            in2 => \N__27907\,
            in3 => \N__27014\,
            lcout => \pid_side.un1_pid_prereg_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29405\,
            in2 => \N__48191\,
            in3 => \N__27011\,
            lcout => \pid_side.un1_pid_prereg_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_9\,
            carryout => \pid_side.un1_pid_prereg_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28420\,
            in2 => \_gnd_net_\,
            in3 => \N__27008\,
            lcout => \pid_side.un1_pid_prereg_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_10\,
            carryout => \pid_side.un1_pid_prereg_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28709\,
            in2 => \N__48190\,
            in3 => \N__27005\,
            lcout => \pid_side.un1_pid_prereg_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_11\,
            carryout => \pid_side.un1_pid_prereg_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30832\,
            in2 => \_gnd_net_\,
            in3 => \N__27002\,
            lcout => \pid_side.un1_pid_prereg_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_12\,
            carryout => \pid_side.un1_pid_prereg_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28234\,
            in2 => \_gnd_net_\,
            in3 => \N__27071\,
            lcout => \pid_side.un1_pid_prereg_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_13\,
            carryout => \pid_side.un1_pid_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28267\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \pid_side.un1_pid_prereg_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_14\,
            carryout => \pid_side.un1_pid_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30922\,
            in2 => \_gnd_net_\,
            in3 => \N__27065\,
            lcout => \pid_side.un1_pid_prereg_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_15\,
            carryout => \pid_side.un1_pid_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28189\,
            in2 => \_gnd_net_\,
            in3 => \N__27062\,
            lcout => \pid_side.un1_pid_prereg_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \pid_side.un1_pid_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28657\,
            in2 => \_gnd_net_\,
            in3 => \N__27059\,
            lcout => \pid_side.un1_pid_prereg_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_17\,
            carryout => \pid_side.un1_pid_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28306\,
            in2 => \_gnd_net_\,
            in3 => \N__27056\,
            lcout => \pid_side.un1_pid_prereg_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_18\,
            carryout => \pid_side.un1_pid_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28146\,
            in2 => \_gnd_net_\,
            in3 => \N__27053\,
            lcout => \pid_side.un1_pid_prereg_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_side.un1_pid_prereg_cry_19\,
            carryout => \pid_side.un1_pid_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_21_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27050\,
            lcout => \pid_side.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51354\,
            ce => \N__41891\,
            sr => \N__49563\
        );

    \Commands_frame_decoder.source_CH2data_ess_7_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40006\,
            lcout => side_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51344\,
            ce => \N__27037\,
            sr => \N__49571\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_0_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42605\,
            lcout => \drone_H_disp_side_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36803\,
            lcout => \drone_H_disp_side_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_2_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37114\,
            lcout => \drone_H_disp_side_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_3_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37034\,
            lcout => \drone_H_disp_side_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_4_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36959\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_5_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36877\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_6_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48436\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_7_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36628\,
            lcout => \dron_frame_decoder_1.drone_H_disp_side_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51337\,
            ce => \N__27098\,
            sr => \N__49582\
        );

    \Commands_frame_decoder.source_alt_ki_7_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40005\,
            in2 => \_gnd_net_\,
            in3 => \N__50801\,
            lcout => alt_ki_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51329\,
            ce => \N__38848\,
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_1__0__0_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27290\,
            lcout => \uart_pc_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_0__0__0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27296\,
            lcout => \uart_pc_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51534\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27284\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27278\,
            lcout => \uart_pc_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.Q_0__0_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27272\,
            lcout => \debug_CH2_18A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__27613\,
            in1 => \N__27266\,
            in2 => \N__27229\,
            in3 => \N__49795\,
            lcout => \Commands_frame_decoder.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_4_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__27193\,
            in1 => \N__28982\,
            in2 => \N__36730\,
            in3 => \N__28949\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51500\,
            ce => 'H',
            sr => \N__49507\
        );

    \uart_pc.data_5_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__28730\,
            in2 => \N__39821\,
            in3 => \N__40041\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__39284\,
            in1 => \N__28829\,
            in2 => \N__28741\,
            in3 => \N__27389\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40299\,
            in2 => \_gnd_net_\,
            in3 => \N__39581\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27605\,
            in1 => \N__40040\,
            in2 => \N__27443\,
            in3 => \N__39283\,
            lcout => \Commands_frame_decoder.N_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__40643\,
            in1 => \N__28791\,
            in2 => \_gnd_net_\,
            in3 => \N__48993\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_4_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__28792\,
            in1 => \N__27358\,
            in2 => \N__27362\,
            in3 => \N__40300\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_4_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29057\,
            in1 => \N__40650\,
            in2 => \N__27359\,
            in3 => \N__40758\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51478\,
            ce => 'H',
            sr => \N__40524\
        );

    \uart_pc.data_Aux_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__30068\,
            in1 => \N__27334\,
            in2 => \N__40676\,
            in3 => \N__40757\,
            lcout => \uart_pc.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51478\,
            ce => 'H',
            sr => \N__40524\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29000\,
            in2 => \N__27323\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27307\,
            in2 => \N__29008\,
            in3 => \N__27314\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_7_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27715\,
            in2 => \N__27311\,
            in3 => \N__27299\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_8_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27700\,
            in2 => \N__27719\,
            in3 => \N__27707\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_9_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27685\,
            in2 => \N__27704\,
            in3 => \N__27692\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_10_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27670\,
            in2 => \N__27689\,
            in3 => \N__27677\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_11_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27655\,
            in2 => \N__27674\,
            in3 => \N__27662\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_12_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27643\,
            in2 => \N__27659\,
            in3 => \N__27647\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__51465\,
            ce => \N__28916\,
            sr => \N__49514\
        );

    \scaler_4.source_data_1_esr_13_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27644\,
            in2 => \N__27632\,
            in3 => \N__27623\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__51449\,
            ce => \N__28911\,
            sr => \N__49517\
        );

    \scaler_4.source_data_1_esr_14_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27620\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51449\,
            ce => \N__28911\,
            sr => \N__49517\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__31042\,
            in1 => \N__29874\,
            in2 => \_gnd_net_\,
            in3 => \N__49022\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29875\,
            in1 => \_gnd_net_\,
            in2 => \N__27617\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.data_rdyc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_i_i_0_a2_2_4_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36749\,
            in1 => \N__36908\,
            in2 => \N__48408\,
            in3 => \N__36996\,
            lcout => \dron_frame_decoder_1.N_412_4\,
            ltout => \dron_frame_decoder_1.N_412_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27806\,
            in3 => \N__27942\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_0_0_a2_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__27802\,
            in1 => \N__29220\,
            in2 => \N__27785\,
            in3 => \N__27764\,
            lcout => \dron_frame_decoder_1.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_1_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28053\,
            in1 => \N__27750\,
            in2 => \N__27947\,
            in3 => \N__29211\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.N_177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__28007\,
            in1 => \N__27751\,
            in2 => \N__27755\,
            in3 => \N__27855\,
            lcout => \dron_frame_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51421\,
            ce => 'H',
            sr => \N__49526\
        );

    \dron_frame_decoder_1.state_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__27725\,
            in1 => \N__27964\,
            in2 => \N__27834\,
            in3 => \N__27854\,
            lcout => \dron_frame_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51421\,
            ce => 'H',
            sr => \N__49526\
        );

    \dron_frame_decoder_1.source_data_valid_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__28054\,
            in1 => \N__32802\,
            in2 => \_gnd_net_\,
            in3 => \N__29212\,
            lcout => \debug_CH1_0A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51421\,
            ce => 'H',
            sr => \N__49526\
        );

    \dron_frame_decoder_1.state_RNI1H181_5_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__29204\,
            in1 => \N__27999\,
            in2 => \N__28121\,
            in3 => \N__49754\,
            lcout => \dron_frame_decoder_1.N_739_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_4_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__28000\,
            in1 => \N__28118\,
            in2 => \N__29222\,
            in3 => \N__27870\,
            lcout => \dron_frame_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51406\,
            ce => 'H',
            sr => \N__49534\
        );

    \dron_frame_decoder_1.state_RNI6P6K_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28114\,
            in2 => \_gnd_net_\,
            in3 => \N__29203\,
            lcout => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4\,
            ltout => \dron_frame_decoder_1.state_RNI6P6KZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_7_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__27872\,
            in1 => \_gnd_net_\,
            in2 => \N__28082\,
            in3 => \N__28077\,
            lcout => \dron_frame_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51406\,
            ce => 'H',
            sr => \N__49534\
        );

    \dron_frame_decoder_1.state_6_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__28058\,
            in1 => \N__29205\,
            in2 => \N__28079\,
            in3 => \N__27871\,
            lcout => \dron_frame_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51406\,
            ce => 'H',
            sr => \N__49534\
        );

    \dron_frame_decoder_1.state_RNO_0_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__28025\,
            in1 => \N__27976\,
            in2 => \N__28016\,
            in3 => \N__27963\,
            lcout => \dron_frame_decoder_1.N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_5_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__29314\,
            in1 => \N__28001\,
            in2 => \_gnd_net_\,
            in3 => \N__27875\,
            lcout => \dron_frame_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51391\,
            ce => 'H',
            sr => \N__49541\
        );

    \dron_frame_decoder_1.state_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27873\,
            in1 => \N__27980\,
            in2 => \N__27946\,
            in3 => \N__27965\,
            lcout => \dron_frame_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51391\,
            ce => 'H',
            sr => \N__49541\
        );

    \pid_side.pid_prereg_9_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__27920\,
            in1 => \N__27908\,
            in2 => \N__50047\,
            in3 => \N__34559\,
            lcout => \pid_side.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51391\,
            ce => 'H',
            sr => \N__49541\
        );

    \dron_frame_decoder_1.state_2_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__27874\,
            in1 => \N__27835\,
            in2 => \N__29243\,
            in3 => \N__29213\,
            lcout => \dron_frame_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51391\,
            ce => 'H',
            sr => \N__49541\
        );

    \pid_side.pid_prereg_8_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__28457\,
            in1 => \N__28451\,
            in2 => \N__50022\,
            in3 => \N__34593\,
            lcout => \pid_side.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51365\,
            ce => 'H',
            sr => \N__49555\
        );

    \pid_side.pid_prereg_11_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__28424\,
            in1 => \N__28394\,
            in2 => \N__50020\,
            in3 => \N__34431\,
            lcout => \pid_side.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51365\,
            ce => 'H',
            sr => \N__49555\
        );

    \pid_side.pid_prereg_4_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__28388\,
            in1 => \N__28382\,
            in2 => \N__50021\,
            in3 => \N__38230\,
            lcout => \pid_side.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51365\,
            ce => 'H',
            sr => \N__49555\
        );

    \pid_side.pid_prereg_6_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__49985\,
            in1 => \N__28352\,
            in2 => \N__34204\,
            in3 => \N__28322\,
            lcout => \pid_side.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51365\,
            ce => 'H',
            sr => \N__49555\
        );

    \pid_side.pid_prereg_19_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__28316\,
            in1 => \N__50027\,
            in2 => \N__28310\,
            in3 => \N__29344\,
            lcout => \pid_side.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51355\,
            ce => 'H',
            sr => \N__49564\
        );

    \pid_side.pid_prereg_15_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__28274\,
            in1 => \N__28244\,
            in2 => \N__50044\,
            in3 => \N__34804\,
            lcout => \pid_side.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51355\,
            ce => 'H',
            sr => \N__49564\
        );

    \pid_side.pid_prereg_14_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__28238\,
            in1 => \N__28205\,
            in2 => \N__34790\,
            in3 => \N__50023\,
            lcout => \pid_side.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51355\,
            ce => 'H',
            sr => \N__49564\
        );

    \pid_side.pid_prereg_17_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__28199\,
            in1 => \N__28193\,
            in2 => \N__50046\,
            in3 => \N__29357\,
            lcout => \pid_side.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51345\,
            ce => 'H',
            sr => \N__49572\
        );

    \pid_side.pid_prereg_20_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__50035\,
            in1 => \N__28154\,
            in2 => \N__29330\,
            in3 => \N__28148\,
            lcout => \pid_side.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51345\,
            ce => 'H',
            sr => \N__49572\
        );

    \pid_side.pid_prereg_12_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__28708\,
            in1 => \N__28676\,
            in2 => \N__50045\,
            in3 => \N__37841\,
            lcout => \pid_side.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51345\,
            ce => 'H',
            sr => \N__49572\
        );

    \pid_side.pid_prereg_18_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__50034\,
            in1 => \N__28670\,
            in2 => \N__28664\,
            in3 => \N__29369\,
            lcout => \pid_side.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51345\,
            ce => 'H',
            sr => \N__49572\
        );

    \pid_alt.error_d_reg_prev_esr_RNISPHM_15_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__28631\,
            in1 => \N__28613\,
            in2 => \_gnd_net_\,
            in3 => \N__28583\,
            lcout => \pid_alt.error_d_reg_prev_esr_RNISPHMZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_axb_8_l_ofx_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__29300\,
            in1 => \_gnd_net_\,
            in2 => \N__28505\,
            in3 => \N__29542\,
            lcout => \pid_side.error_axb_8_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_axb_7_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28501\,
            in2 => \_gnd_net_\,
            in3 => \N__29299\,
            lcout => \pid_side.error_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_2_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28478\,
            lcout => \pid_front.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_2_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37113\,
            lcout => \drone_H_disp_front_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51330\,
            ce => \N__42509\,
            sr => \N__49590\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37022\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_front_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51330\,
            ce => \N__42509\,
            sr => \N__49590\
        );

    \pid_side.error_axb_1_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28472\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_RNO_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31177\,
            in2 => \_gnd_net_\,
            in3 => \N__49776\,
            lcout => \pid_alt.state_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32018\,
            lcout => pid_altitude_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51490\,
            ce => \N__28811\,
            sr => \N__49503\
        );

    \uart_pc.state_RNO_0_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__32146\,
            in1 => \N__40705\,
            in2 => \_gnd_net_\,
            in3 => \N__49777\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__29795\,
            in1 => \N__31100\,
            in2 => \N__28805\,
            in3 => \N__31265\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__48988\,
            in1 => \N__31261\,
            in2 => \N__31110\,
            in3 => \N__29789\,
            lcout => \uart_pc.N_143\,
            ltout => \uart_pc.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__29696\,
            in1 => \N__29750\,
            in2 => \N__28802\,
            in3 => \N__48989\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__29028\,
            in1 => \N__31010\,
            in2 => \N__30953\,
            in3 => \N__49780\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__31334\,
            in1 => \N__31306\,
            in2 => \N__31109\,
            in3 => \N__29788\,
            lcout => \uart_pc.data_rdyc_1\,
            ltout => \uart_pc.data_rdyc_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIMQ8T1_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28778\,
            in3 => \N__48987\,
            lcout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__32958\,
            in1 => \N__31009\,
            in2 => \N__29030\,
            in3 => \N__49779\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__29029\,
            in1 => \N__33100\,
            in2 => \N__29012\,
            in3 => \N__33023\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_5_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29009\,
            in1 => \N__28981\,
            in2 => \_gnd_net_\,
            in3 => \N__28948\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51451\,
            ce => \N__28912\,
            sr => \N__49511\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__29998\,
            in1 => \N__30052\,
            in2 => \_gnd_net_\,
            in3 => \N__29952\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__29953\,
            in1 => \_gnd_net_\,
            in2 => \N__30056\,
            in3 => \N__29999\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIEAGS_4_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__29791\,
            in1 => \N__30140\,
            in2 => \_gnd_net_\,
            in3 => \N__49758\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__40749\,
            in1 => \N__29039\,
            in2 => \N__28873\,
            in3 => \N__40694\,
            lcout => \uart_pc.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51436\,
            ce => 'H',
            sr => \N__40528\
        );

    \uart_pc.data_Aux_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29900\,
            in1 => \N__40691\,
            in2 => \N__28852\,
            in3 => \N__40748\,
            lcout => \uart_pc.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51436\,
            ce => 'H',
            sr => \N__40528\
        );

    \uart_pc.data_Aux_3_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__28835\,
            in1 => \N__40692\,
            in2 => \N__28828\,
            in3 => \N__40750\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51436\,
            ce => 'H',
            sr => \N__40528\
        );

    \uart_pc.data_Aux_5_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__29045\,
            in1 => \N__40693\,
            in2 => \N__29074\,
            in3 => \N__40751\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51436\,
            ce => 'H',
            sr => \N__40528\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__29990\,
            in1 => \N__30038\,
            in2 => \_gnd_net_\,
            in3 => \N__29941\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__29942\,
            in1 => \_gnd_net_\,
            in2 => \N__30046\,
            in3 => \N__29991\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__29989\,
            in1 => \N__30037\,
            in2 => \_gnd_net_\,
            in3 => \N__29940\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_esr_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29893\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51407\,
            ce => \N__29284\,
            sr => \N__29266\
        );

    \uart_drone.data_esr_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30262\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51407\,
            ce => \N__29284\,
            sr => \N__29266\
        );

    \uart_drone.data_esr_5_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30224\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51407\,
            ce => \N__29284\,
            sr => \N__29266\
        );

    \uart_drone.data_esr_7_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30197\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51407\,
            ce => \N__29284\,
            sr => \N__29266\
        );

    \uart_drone.data_esr_3_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30248\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51393\,
            ce => \N__29291\,
            sr => \N__29267\
        );

    \uart_drone.data_esr_4_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30236\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51393\,
            ce => \N__29291\,
            sr => \N__29267\
        );

    \uart_drone.data_esr_1_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30275\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51393\,
            ce => \N__29291\,
            sr => \N__29267\
        );

    \uart_drone.data_esr_6_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51393\,
            ce => \N__29291\,
            sr => \N__29267\
        );

    \pid_alt.source_pid_1_10_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__31854\,
            in1 => \N__32016\,
            in2 => \N__32492\,
            in3 => \N__29144\,
            lcout => throttle_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51379\,
            ce => 'H',
            sr => \N__31774\
        );

    \pid_alt.source_pid_1_6_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__31855\,
            in1 => \N__29450\,
            in2 => \N__32672\,
            in3 => \N__32017\,
            lcout => throttle_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51379\,
            ce => 'H',
            sr => \N__31774\
        );

    \pid_alt.source_pid_1_8_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__32015\,
            in1 => \N__31856\,
            in2 => \N__37794\,
            in3 => \N__29105\,
            lcout => throttle_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51379\,
            ce => 'H',
            sr => \N__31774\
        );

    \dron_frame_decoder_1.state_RNI4N6K_2_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29238\,
            in2 => \_gnd_net_\,
            in3 => \N__29221\,
            lcout => \dron_frame_decoder_1.state_RNI4N6KZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIT3KA1_10_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29139\,
            in1 => \N__30180\,
            in2 => \N__31807\,
            in3 => \N__29097\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIFQKS1_11_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32046\,
            in2 => \N__29108\,
            in3 => \N__29448\,
            lcout => \pid_alt.N_530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNINTJA1_11_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32047\,
            in1 => \N__30181\,
            in2 => \N__31574\,
            in3 => \N__29098\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_i_a5_1_10_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIFBU82_6_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31803\,
            in1 => \N__30490\,
            in2 => \N__29453\,
            in3 => \N__29449\,
            lcout => \pid_alt.un1_reset_i_a5_1_10_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIEKJA1_1_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30610\,
            in1 => \N__31495\,
            in2 => \N__30543\,
            in3 => \N__31528\,
            lcout => \pid_alt.un1_reset_i_a5_0_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNI8LUI1_6_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34586\,
            in1 => \N__34560\,
            in2 => \N__34200\,
            in3 => \N__34247\,
            lcout => \pid_side.un1_reset_i_a5_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_10_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__34249\,
            in1 => \N__29417\,
            in2 => \N__49978\,
            in3 => \N__29404\,
            lcout => \pid_side.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51347\,
            ce => 'H',
            sr => \N__49556\
        );

    \pid_side.pid_prereg_RNIUDBG1_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34400\,
            in1 => \N__34193\,
            in2 => \N__34594\,
            in3 => \N__34561\,
            lcout => OPEN,
            ltout => \pid_side.un1_reset_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNIHJND2_10_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__34248\,
            in1 => \_gnd_net_\,
            in2 => \N__29372\,
            in3 => \N__34430\,
            lcout => \pid_side.N_531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNIT3QQ1_17_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29368\,
            in1 => \N__29356\,
            in2 => \N__29345\,
            in3 => \N__29326\,
            lcout => \pid_side.m7_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI14DT_2_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29315\,
            in2 => \_gnd_net_\,
            in3 => \N__49770\,
            lcout => \dron_frame_decoder_1.N_731_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_11_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37010\,
            lcout => \drone_H_disp_side_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51317\,
            ce => \N__29580\,
            sr => \N__49591\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_12_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36934\,
            lcout => \drone_H_disp_side_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51317\,
            ce => \N__29580\,
            sr => \N__49591\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_13_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36844\,
            lcout => \drone_H_disp_side_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51317\,
            ce => \N__29580\,
            sr => \N__49591\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_14_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48433\,
            lcout => \drone_H_disp_side_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51317\,
            ce => \N__29580\,
            sr => \N__49591\
        );

    \dron_frame_decoder_1.source_H_disp_side_esr_RNIV6RD_12_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_side_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_3_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29510\,
            lcout => \pid_front.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_3_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39373\,
            in2 => \_gnd_net_\,
            in3 => \N__50798\,
            lcout => xy_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51310\,
            ce => \N__39031\,
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29465\,
            lcout => \uart_drone_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__29759\,
            in1 => \N__48910\,
            in2 => \N__29692\,
            in3 => \N__29825\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__29717\,
            in1 => \N__29647\,
            in2 => \N__29722\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31332\,
            in2 => \_gnd_net_\,
            in3 => \N__29753\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31303\,
            in2 => \_gnd_net_\,
            in3 => \N__29744\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31098\,
            in2 => \_gnd_net_\,
            in3 => \N__29741\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__31099\,
            in1 => \N__31304\,
            in2 => \N__30152\,
            in3 => \N__32172\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__29738\,
            in1 => \N__29820\,
            in2 => \N__29690\,
            in3 => \N__48970\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__29721\,
            in1 => \N__29819\,
            in2 => \N__29689\,
            in3 => \N__48969\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__31260\,
            in1 => \N__30139\,
            in2 => \N__29732\,
            in3 => \N__29790\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29723\,
            in2 => \_gnd_net_\,
            in3 => \N__29648\,
            lcout => OPEN,
            ltout => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__48967\,
            in1 => \N__29691\,
            in2 => \N__29651\,
            in3 => \N__29821\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__33153\,
            in1 => \N__33004\,
            in2 => \N__33091\,
            in3 => \N__32463\,
            lcout => \uart_drone.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.Q_0__0_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29849\,
            lcout => \debug_CH0_16A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__33005\,
            in1 => \N__32912\,
            in2 => \N__32967\,
            in3 => \N__33075\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => \uart_drone.timer_Count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__32438\,
            in1 => \N__32342\,
            in2 => \N__29840\,
            in3 => \N__48968\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__30137\,
            in1 => \N__31108\,
            in2 => \N__32189\,
            in3 => \N__31293\,
            lcout => OPEN,
            ltout => \uart_pc.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__48966\,
            in1 => \N__29834\,
            in2 => \N__29837\,
            in3 => \N__32188\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__31292\,
            in1 => \N__40575\,
            in2 => \N__31112\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.N_144_1\,
            ltout => \uart_pc.N_144_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_4_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__30138\,
            in1 => \N__48965\,
            in2 => \N__29828\,
            in3 => \N__29818\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110011"
        )
    port map (
            in0 => \N__31291\,
            in1 => \N__29787\,
            in2 => \N__31111\,
            in3 => \N__30136\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29983\,
            in1 => \N__30030\,
            in2 => \_gnd_net_\,
            in3 => \N__29933\,
            lcout => \uart_pc.N_152\,
            ltout => \uart_pc.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30088\,
            in2 => \N__30155\,
            in3 => \N__30144\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_9_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__31414\,
            in1 => \N__31391\,
            in2 => \N__46170\,
            in3 => \N__35641\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51408\,
            ce => 'H',
            sr => \N__49522\
        );

    \uart_pc.bit_Count_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001001010000"
        )
    port map (
            in0 => \N__30097\,
            in1 => \N__40585\,
            in2 => \N__29951\,
            in3 => \N__30151\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51408\,
            ce => 'H',
            sr => \N__49522\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29936\,
            in2 => \_gnd_net_\,
            in3 => \N__30096\,
            lcout => OPEN,
            ltout => \uart_pc.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__30077\,
            in1 => \N__29988\,
            in2 => \N__30101\,
            in3 => \N__30036\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51408\,
            ce => 'H',
            sr => \N__49522\
        );

    \uart_pc.bit_Count_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__29954\,
            in1 => \N__30098\,
            in2 => \N__30045\,
            in3 => \N__30076\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51408\,
            ce => 'H',
            sr => \N__49522\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29934\,
            in1 => \N__29984\,
            in2 => \_gnd_net_\,
            in3 => \N__30031\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__30032\,
            in1 => \_gnd_net_\,
            in2 => \N__29997\,
            in3 => \N__29935\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__31021\,
            in1 => \N__30161\,
            in2 => \N__29894\,
            in3 => \N__31238\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31234\,
            in1 => \N__30274\,
            in2 => \N__31047\,
            in3 => \N__30335\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__31586\,
            in1 => \N__31025\,
            in2 => \N__30263\,
            in3 => \N__31239\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31235\,
            in1 => \N__30247\,
            in2 => \N__31048\,
            in3 => \N__30326\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__30320\,
            in1 => \N__30235\,
            in2 => \N__31046\,
            in3 => \N__31240\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__30223\,
            in2 => \N__31049\,
            in3 => \N__30698\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__30560\,
            in1 => \N__31026\,
            in2 => \N__30212\,
            in3 => \N__31241\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \uart_drone.data_Aux_7_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__31237\,
            in1 => \N__30196\,
            in2 => \N__31050\,
            in3 => \N__32096\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51394\,
            ce => 'H',
            sr => \N__33122\
        );

    \pid_alt.source_pid_1_9_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__31853\,
            in1 => \N__32030\,
            in2 => \N__31415\,
            in3 => \N__30185\,
            lcout => throttle_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51380\,
            ce => 'H',
            sr => \N__31778\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__31724\,
            in1 => \N__31654\,
            in2 => \_gnd_net_\,
            in3 => \N__34535\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__34537\,
            in1 => \_gnd_net_\,
            in2 => \N__31663\,
            in3 => \N__31725\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__34538\,
            in1 => \_gnd_net_\,
            in2 => \N__31664\,
            in3 => \N__31726\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31727\,
            in1 => \N__31661\,
            in2 => \_gnd_net_\,
            in3 => \N__34536\,
            lcout => \uart_drone.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_13_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__30410\,
            in1 => \N__30451\,
            in2 => \_gnd_net_\,
            in3 => \N__30505\,
            lcout => throttle_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51367\,
            ce => \N__31598\,
            sr => \N__31769\
        );

    \pid_alt.source_pid_1_esr_12_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__30506\,
            in1 => \N__30548\,
            in2 => \N__30460\,
            in3 => \N__30409\,
            lcout => throttle_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51367\,
            ce => \N__31598\,
            sr => \N__31769\
        );

    \pid_alt.source_pid_1_esr_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__31852\,
            in1 => \_gnd_net_\,
            in2 => \N__30674\,
            in3 => \N__30658\,
            lcout => throttle_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51367\,
            ce => \N__31598\,
            sr => \N__31769\
        );

    \pid_alt.source_pid_1_esr_4_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__31851\,
            in2 => \N__30614\,
            in3 => \N__30670\,
            lcout => throttle_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51367\,
            ce => \N__31598\,
            sr => \N__31769\
        );

    \pid_alt.pid_prereg_esr_RNIG5AU_0_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30499\,
            in1 => \N__30638\,
            in2 => \_gnd_net_\,
            in3 => \N__31563\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_i_a5_0_6_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI2R305_0_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30314\,
            in1 => \N__30308\,
            in2 => \N__30278\,
            in3 => \N__30685\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_i_a5_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI1RJPB_10_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__30719\,
            in1 => \N__30713\,
            in2 => \N__30704\,
            in3 => \N__30399\,
            lcout => OPEN,
            ltout => \pid_alt.pid_prereg_esr_RNI1RJPBZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI65QMC_24_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30459\,
            in1 => \N__32023\,
            in2 => \N__30701\,
            in3 => \N__48961\,
            lcout => \pid_alt.pid_prereg_esr_RNI65QMCZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__31662\,
            in1 => \N__34525\,
            in2 => \_gnd_net_\,
            in3 => \N__31714\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIJ6482_24_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30492\,
            in1 => \N__30458\,
            in2 => \_gnd_net_\,
            in3 => \N__30686\,
            lcout => \pid_alt.N_535\,
            ltout => \pid_alt.N_535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI70AB5_4_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__31833\,
            in1 => \N__30657\,
            in2 => \N__30617\,
            in3 => \N__30609\,
            lcout => \pid_alt.N_472_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46157\,
            in2 => \_gnd_net_\,
            in3 => \N__49760\,
            lcout => \ppm_encoder_1.pid_altitude_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__31640\,
            in1 => \N__31703\,
            in2 => \_gnd_net_\,
            in3 => \N__34514\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIHKIA2_12_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__30536\,
            in1 => \N__30491\,
            in2 => \N__30461\,
            in3 => \N__30408\,
            lcout => \pid_alt.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_7_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__30377\,
            in1 => \N__30368\,
            in2 => \N__49977\,
            in3 => \N__34401\,
            lcout => \pid_side.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \pid_side.state_0_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49926\,
            in1 => \N__32831\,
            in2 => \_gnd_net_\,
            in3 => \N__35867\,
            lcout => \pid_side.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \pid_side.pid_prereg_3_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__49930\,
            in1 => \N__50114\,
            in2 => \N__35787\,
            in3 => \N__30932\,
            lcout => \pid_side.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \pid_side.pid_prereg_16_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__30923\,
            in1 => \N__30890\,
            in2 => \N__49975\,
            in3 => \N__34753\,
            lcout => \pid_side.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \pid_side.pid_prereg_5_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__30878\,
            in1 => \N__30869\,
            in2 => \N__49976\,
            in3 => \N__38117\,
            lcout => \pid_side.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \ppm_encoder_1.rudder_6_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__46194\,
            in1 => \N__31211\,
            in2 => \_gnd_net_\,
            in3 => \N__38775\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51338\,
            ce => 'H',
            sr => \N__49565\
        );

    \pid_side.state_1_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51323\,
            ce => 'H',
            sr => \N__49583\
        );

    \pid_side.pid_prereg_13_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__30839\,
            in1 => \N__30809\,
            in2 => \N__50039\,
            in3 => \N__38284\,
            lcout => \pid_side.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51318\,
            ce => 'H',
            sr => \N__49592\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_1_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39641\,
            in2 => \_gnd_net_\,
            in3 => \N__50799\,
            lcout => xy_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51314\,
            ce => \N__39027\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_xy_kp_e_0_6_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40013\,
            in2 => \_gnd_net_\,
            in3 => \N__50800\,
            lcout => xy_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51314\,
            ce => \N__39027\,
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_1_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__42802\,
            in1 => \N__48785\,
            in2 => \_gnd_net_\,
            in3 => \N__32216\,
            lcout => \pid_front.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51311\,
            ce => 'H',
            sr => \N__49600\
        );

    \pid_front.state_RNIPKTD_0_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__42726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49769\,
            lcout => \pid_front.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIH1EN_0_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31163\,
            in2 => \_gnd_net_\,
            in3 => \N__49753\,
            lcout => \pid_alt.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__31101\,
            in1 => \N__31310\,
            in2 => \N__32135\,
            in3 => \N__32156\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__30943\,
            in1 => \N__31011\,
            in2 => \_gnd_net_\,
            in3 => \N__49778\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__32362\,
            in1 => \N__33081\,
            in2 => \N__30956\,
            in3 => \N__33171\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__48977\,
            in1 => \N__32423\,
            in2 => \N__32417\,
            in3 => \N__32339\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__32335\,
            in2 => \N__32415\,
            in3 => \N__48980\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32385\,
            in2 => \_gnd_net_\,
            in3 => \N__32117\,
            lcout => OPEN,
            ltout => \uart_drone.timer_Count_RNO_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__32405\,
            in1 => \N__32334\,
            in2 => \N__31337\,
            in3 => \N__48979\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31333\,
            in2 => \_gnd_net_\,
            in3 => \N__31305\,
            lcout => \uart_pc.N_126_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33006\,
            in2 => \_gnd_net_\,
            in3 => \N__32464\,
            lcout => \uart_drone.N_126_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__32908\,
            in1 => \N__32936\,
            in2 => \N__32341\,
            in3 => \N__48978\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__32907\,
            in2 => \N__32105\,
            in3 => \N__33158\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31204\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32245\,
            in2 => \_gnd_net_\,
            in3 => \N__31187\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32269\,
            in2 => \_gnd_net_\,
            in3 => \N__31184\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34978\,
            in2 => \_gnd_net_\,
            in3 => \N__31181\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34045\,
            in3 => \N__31370\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32638\,
            in2 => \_gnd_net_\,
            in3 => \N__31367\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32299\,
            in2 => \_gnd_net_\,
            in3 => \N__31364\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32584\,
            in2 => \N__48043\,
            in3 => \N__31361\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31358\,
            in2 => \_gnd_net_\,
            in3 => \N__31349\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51392\,
            ce => \N__36693\,
            sr => \N__49527\
        );

    \ppm_encoder_1.un1_throttle_cry_0_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44034\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35517\,
            in2 => \N__48040\,
            in3 => \N__31346\,
            lcout => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_0\,
            carryout => \ppm_encoder_1.un1_throttle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32544\,
            in2 => \_gnd_net_\,
            in3 => \N__31343\,
            lcout => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_1\,
            carryout => \ppm_encoder_1.un1_throttle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32733\,
            in2 => \N__48041\,
            in3 => \N__31340\,
            lcout => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_2\,
            carryout => \ppm_encoder_1.un1_throttle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46438\,
            in2 => \_gnd_net_\,
            in3 => \N__31430\,
            lcout => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_3\,
            carryout => \ppm_encoder_1.un1_throttle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32701\,
            in3 => \N__31427\,
            lcout => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_4\,
            carryout => \ppm_encoder_1.un1_throttle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32670\,
            in2 => \N__48042\,
            in3 => \N__31424\,
            lcout => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_5\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45534\,
            in2 => \_gnd_net_\,
            in3 => \N__31421\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37795\,
            in2 => \_gnd_net_\,
            in3 => \N__31418\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31407\,
            in2 => \_gnd_net_\,
            in3 => \N__31382\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32490\,
            in2 => \_gnd_net_\,
            in3 => \N__31379\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32616\,
            in2 => \_gnd_net_\,
            in3 => \N__31376\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32752\,
            in2 => \_gnd_net_\,
            in3 => \N__31373\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47885\,
            in2 => \N__41512\,
            in3 => \N__31604\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31601\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51366\,
            ce => \N__36698\,
            sr => \N__49542\
        );

    \pid_alt.state_RNIRQ15D_1_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32014\,
            in2 => \_gnd_net_\,
            in3 => \N__31768\,
            lcout => \pid_alt.N_72_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46667\,
            in1 => \N__31742\,
            in2 => \_gnd_net_\,
            in3 => \N__38657\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31641\,
            in1 => \N__31713\,
            in2 => \_gnd_net_\,
            in3 => \N__34517\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31442\,
            in1 => \N__31570\,
            in2 => \N__44038\,
            in3 => \N__32028\,
            lcout => throttle_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \pid_alt.source_pid_1_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__32025\,
            in1 => \N__31443\,
            in2 => \N__31535\,
            in3 => \N__35521\,
            lcout => throttle_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \pid_alt.source_pid_1_2_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__31444\,
            in1 => \N__31499\,
            in2 => \N__32546\,
            in3 => \N__32029\,
            lcout => throttle_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \pid_alt.source_pid_1_3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__32026\,
            in1 => \N__31465\,
            in2 => \N__32735\,
            in3 => \N__31445\,
            lcout => throttle_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \pid_alt.source_pid_1_11_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__32024\,
            in1 => \N__31842\,
            in2 => \N__32618\,
            in3 => \N__32054\,
            lcout => throttle_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \pid_alt.source_pid_1_7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__32027\,
            in1 => \N__31843\,
            in2 => \N__45544\,
            in3 => \N__31808\,
            lcout => throttle_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51346\,
            ce => 'H',
            sr => \N__31770\
        );

    \uart_drone.state_RNI62411_4_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__33095\,
            in1 => \N__33027\,
            in2 => \N__32896\,
            in3 => \N__33172\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39152\,
            in1 => \N__38806\,
            in2 => \_gnd_net_\,
            in3 => \N__46788\,
            lcout => \ppm_encoder_1.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46787\,
            in1 => \N__35621\,
            in2 => \_gnd_net_\,
            in3 => \N__38429\,
            lcout => \ppm_encoder_1.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI63LK2_3_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000100"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__34466\,
            in2 => \N__32092\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => \uart_drone.un1_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__34468\,
            in1 => \N__34516\,
            in2 => \N__31733\,
            in3 => \N__31701\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51331\,
            ce => 'H',
            sr => \N__49573\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31700\,
            in1 => \N__31626\,
            in2 => \_gnd_net_\,
            in3 => \N__34502\,
            lcout => \uart_drone.N_152\,
            ltout => \uart_drone.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011001000100"
        )
    port map (
            in0 => \N__34467\,
            in1 => \N__34515\,
            in2 => \N__31730\,
            in3 => \N__32898\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51331\,
            ce => 'H',
            sr => \N__49573\
        );

    \uart_drone.bit_Count_2_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__31702\,
            in1 => \N__31627\,
            in2 => \N__31673\,
            in3 => \N__34448\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51331\,
            ce => 'H',
            sr => \N__49573\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32085\,
            in1 => \N__33096\,
            in2 => \_gnd_net_\,
            in3 => \N__33028\,
            lcout => \uart_drone.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32066\,
            in1 => \N__33679\,
            in2 => \N__35731\,
            in3 => \N__36235\,
            lcout => front_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51322\,
            ce => 'H',
            sr => \N__33533\
        );

    \pid_front.source_pid_1_1_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33680\,
            in1 => \N__32067\,
            in2 => \N__36196\,
            in3 => \N__32222\,
            lcout => front_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51322\,
            ce => 'H',
            sr => \N__33533\
        );

    \pid_front.source_pid_1_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32068\,
            in1 => \N__33681\,
            in2 => \N__39250\,
            in3 => \N__36401\,
            lcout => front_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51322\,
            ce => 'H',
            sr => \N__33533\
        );

    \pid_front.source_pid_1_3_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__38900\,
            in1 => \N__32069\,
            in2 => \N__33686\,
            in3 => \N__36147\,
            lcout => front_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51322\,
            ce => 'H',
            sr => \N__33533\
        );

    \pid_front.pid_prereg_RNI9EOL_10_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33401\,
            in1 => \N__34891\,
            in2 => \_gnd_net_\,
            in3 => \N__33730\,
            lcout => \pid_front.N_532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIH2151_21_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__34854\,
            in1 => \N__48537\,
            in2 => \_gnd_net_\,
            in3 => \N__33412\,
            lcout => \pid_front.N_533\,
            ltout => \pid_front.N_533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIC5I03_4_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__38937\,
            in1 => \N__33572\,
            in2 => \N__32072\,
            in3 => \N__38973\,
            lcout => \pid_front.N_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIE0SA_1_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__34853\,
            in1 => \N__38936\,
            in2 => \_gnd_net_\,
            in3 => \N__32221\,
            lcout => OPEN,
            ltout => \pid_front.un1_reset_i_a5_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNISBN11_2_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32228\,
            in1 => \N__33678\,
            in2 => \N__32231\,
            in3 => \N__36397\,
            lcout => \pid_front.un1_reset_i_a5_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_RNIJ92F_0_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__38899\,
            in1 => \N__36454\,
            in2 => \N__38975\,
            in3 => \N__36236\,
            lcout => \pid_front.un1_reset_i_a5_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNI75JF_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__36452\,
            in1 => \N__36396\,
            in2 => \N__33685\,
            in3 => \N__32217\,
            lcout => \pid_front.un1_reset_i_a5_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIQBDL1_12_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__36453\,
            in1 => \N__34642\,
            in2 => \N__48536\,
            in3 => \N__34847\,
            lcout => \pid_front.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_1_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36789\,
            lcout => \drone_H_disp_front_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51309\,
            ce => \N__42519\,
            sr => \N__49601\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_8_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42601\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51306\,
            ce => \N__48344\,
            sr => \N__49611\
        );

    \uart_pc.state_RNO_0_2_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110010"
        )
    port map (
            in0 => \N__32130\,
            in1 => \N__40700\,
            in2 => \N__32179\,
            in3 => \N__49774\,
            lcout => \uart_pc.state_srsts_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_1_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__49775\,
            in1 => \N__32150\,
            in2 => \N__40711\,
            in3 => \N__32131\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__32384\,
            in1 => \N__32116\,
            in2 => \N__32387\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32465\,
            in2 => \_gnd_net_\,
            in3 => \N__32441\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33022\,
            in2 => \_gnd_net_\,
            in3 => \N__32429\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32426\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__48957\,
            in1 => \N__32416\,
            in2 => \N__32340\,
            in3 => \N__32386\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33076\,
            in1 => \N__48956\,
            in2 => \N__32363\,
            in3 => \N__33157\,
            lcout => \uart_drone.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_0_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42671\,
            in1 => \N__32834\,
            in2 => \_gnd_net_\,
            in3 => \N__33663\,
            lcout => \pid_front.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51423\,
            ce => 'H',
            sr => \N__49528\
        );

    \ppm_encoder_1.rudder_12_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32300\,
            in1 => \N__32285\,
            in2 => \N__46188\,
            in3 => \N__34140\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51423\,
            ce => 'H',
            sr => \N__49528\
        );

    \ppm_encoder_1.rudder_8_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__32279\,
            in1 => \N__32273\,
            in2 => \N__37605\,
            in3 => \N__46140\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51423\,
            ce => 'H',
            sr => \N__49528\
        );

    \ppm_encoder_1.rudder_7_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32255\,
            in1 => \N__32249\,
            in2 => \N__46189\,
            in3 => \N__45954\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51423\,
            ce => 'H',
            sr => \N__49528\
        );

    \ppm_encoder_1.rudder_11_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32639\,
            in1 => \N__32624\,
            in2 => \N__46187\,
            in3 => \N__35268\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51423\,
            ce => 'H',
            sr => \N__49528\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__46786\,
            in1 => \N__49781\,
            in2 => \N__46666\,
            in3 => \N__44914\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_3_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__36125\,
            in1 => \N__36152\,
            in2 => \N__41971\,
            in3 => \N__46365\,
            lcout => \ppm_encoder_1.elevatorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51395\,
            ce => 'H',
            sr => \N__49543\
        );

    \pid_front.state_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42695\,
            lcout => \pid_front.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51395\,
            ce => 'H',
            sr => \N__49543\
        );

    \ppm_encoder_1.throttle_11_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32617\,
            in1 => \N__32591\,
            in2 => \N__46388\,
            in3 => \N__34001\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51395\,
            ce => 'H',
            sr => \N__49543\
        );

    \ppm_encoder_1.rudder_13_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__32585\,
            in1 => \N__32561\,
            in2 => \N__41691\,
            in3 => \N__46366\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51395\,
            ce => 'H',
            sr => \N__49543\
        );

    \ppm_encoder_1.throttle_2_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32552\,
            in1 => \N__32545\,
            in2 => \N__46389\,
            in3 => \N__37737\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51395\,
            ce => 'H',
            sr => \N__49543\
        );

    \ppm_encoder_1.ppm_output_reg_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110010011110100"
        )
    port map (
            in0 => \N__42128\,
            in1 => \N__42233\,
            in2 => \N__32515\,
            in3 => \N__42104\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.throttle_10_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__32498\,
            in1 => \N__32491\,
            in2 => \N__46304\,
            in3 => \N__35619\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.throttle_12_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__32765\,
            in1 => \N__46242\,
            in2 => \N__34109\,
            in3 => \N__32759\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.throttle_3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__32741\,
            in1 => \N__32734\,
            in2 => \N__46305\,
            in3 => \N__42016\,
            lcout => \ppm_encoder_1.throttleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.throttle_5_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__32708\,
            in1 => \N__46243\,
            in2 => \N__38017\,
            in3 => \N__32702\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.throttle_6_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__32678\,
            in1 => \N__32671\,
            in2 => \N__46306\,
            in3 => \N__38802\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51381\,
            ce => 'H',
            sr => \N__49548\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__43766\,
            in1 => \N__40895\,
            in2 => \_gnd_net_\,
            in3 => \N__34142\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__43880\,
            in1 => \_gnd_net_\,
            in2 => \N__32645\,
            in3 => \N__41207\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_2_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46766\,
            in1 => \N__39214\,
            in2 => \_gnd_net_\,
            in3 => \N__37741\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46631\,
            in2 => \N__32642\,
            in3 => \N__37718\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_3_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46765\,
            in1 => \N__41970\,
            in2 => \_gnd_net_\,
            in3 => \N__42015\,
            lcout => \ppm_encoder_1.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_13_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__33386\,
            in1 => \N__33347\,
            in2 => \_gnd_net_\,
            in3 => \N__33320\,
            lcout => \pid_alt.error_i_acummZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51368\,
            ce => \N__33263\,
            sr => \N__33226\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38558\,
            in1 => \N__33110\,
            in2 => \_gnd_net_\,
            in3 => \N__46632\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__32895\,
            in1 => \N__33173\,
            in2 => \_gnd_net_\,
            in3 => \N__49765\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.state_RNI26LH_1_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42694\,
            in1 => \N__32832\,
            in2 => \_gnd_net_\,
            in3 => \N__33657\,
            lcout => \pid_front.state_ns_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38016\,
            in1 => \N__46767\,
            in2 => \_gnd_net_\,
            in3 => \N__39098\,
            lcout => \ppm_encoder_1.N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__32894\,
            in1 => \N__33104\,
            in2 => \N__33035\,
            in3 => \N__32968\,
            lcout => OPEN,
            ltout => \uart_drone.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__32969\,
            in1 => \N__32932\,
            in2 => \N__32915\,
            in3 => \N__49026\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.state_RNIQ7UK_1_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__50012\,
            in1 => \N__32833\,
            in2 => \_gnd_net_\,
            in3 => \N__35897\,
            lcout => OPEN,
            ltout => \pid_side.state_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.state_RNINK4U_1_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33473\,
            in3 => \N__49025\,
            lcout => \pid_side.state_RNINK4UZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.state_RNIL5IF_0_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__49766\,
            in1 => \_gnd_net_\,
            in2 => \N__50040\,
            in3 => \_gnd_net_\,
            lcout => \pid_side.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_0_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42571\,
            lcout => drone_altitude_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51348\,
            ce => \N__33469\,
            sr => \N__49574\
        );

    \pid_front.pid_prereg_esr_RNIQ3AH3_21_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__33656\,
            in1 => \N__49024\,
            in2 => \N__48535\,
            in3 => \N__33488\,
            lcout => OPEN,
            ltout => \pid_front.un1_reset_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNI2A6A6_2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__34643\,
            in1 => \N__33425\,
            in2 => \N__33416\,
            in3 => \N__33413\,
            lcout => \pid_front.pid_prereg_RNI2A6A6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIEQ7C_6_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34924\,
            in1 => \N__42640\,
            in2 => \N__36521\,
            in3 => \N__36484\,
            lcout => \pid_front.un1_reset_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_6_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__36485\,
            in1 => \N__39171\,
            in2 => \N__33598\,
            in3 => \N__33661\,
            lcout => front_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.source_pid_1_7_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__36520\,
            in1 => \N__33593\,
            in2 => \N__45601\,
            in3 => \N__33664\,
            lcout => front_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.source_pid_1_8_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__42641\,
            in1 => \N__37491\,
            in2 => \N__33599\,
            in3 => \N__33662\,
            lcout => front_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.source_pid_1_9_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__34925\,
            in1 => \N__33597\,
            in2 => \N__36090\,
            in3 => \N__33665\,
            lcout => front_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.source_pid_1_10_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__33588\,
            in1 => \N__33659\,
            in2 => \N__38465\,
            in3 => \N__33731\,
            lcout => front_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.source_pid_1_11_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__33660\,
            in1 => \N__33589\,
            in2 => \N__36333\,
            in3 => \N__34892\,
            lcout => front_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51332\,
            ce => 'H',
            sr => \N__33519\
        );

    \pid_front.state_RNIVITE6_1_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33658\,
            in2 => \_gnd_net_\,
            in3 => \N__33510\,
            lcout => \pid_front.state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.source_pid_1_esr_5_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__33574\,
            in1 => \N__33553\,
            in2 => \_gnd_net_\,
            in3 => \N__38938\,
            lcout => front_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51324\,
            ce => \N__33542\,
            sr => \N__33526\
        );

    \pid_front.source_pid_1_esr_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__38939\,
            in1 => \N__33573\,
            in2 => \N__33554\,
            in3 => \N__38974\,
            lcout => front_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51324\,
            ce => \N__33542\,
            sr => \N__33526\
        );

    \pid_front.source_pid_1_esr_12_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__36455\,
            in2 => \N__48542\,
            in3 => \N__34640\,
            lcout => front_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51324\,
            ce => \N__33542\,
            sr => \N__33526\
        );

    \pid_front.source_pid_1_esr_13_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__34641\,
            in1 => \N__34856\,
            in2 => \_gnd_net_\,
            in3 => \N__48538\,
            lcout => front_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51324\,
            ce => \N__33542\,
            sr => \N__33526\
        );

    \pid_front.pid_prereg_RNI86SO2_1_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36206\,
            in1 => \N__33494\,
            in2 => \N__33743\,
            in3 => \N__34633\,
            lcout => \pid_front.N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_1_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33479\,
            lcout => \pid_front.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIO5UD_6_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36478\,
            in1 => \N__42639\,
            in2 => \N__34917\,
            in3 => \N__33717\,
            lcout => OPEN,
            ltout => \pid_front.un1_reset_i_a5_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNIPQGQ_7_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__34877\,
            in2 => \N__33746\,
            in3 => \N__36510\,
            lcout => \pid_front.un1_reset_i_a5_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_10_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__48266\,
            in1 => \N__50459\,
            in2 => \N__42771\,
            in3 => \N__33723\,
            lcout => \pid_front.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51307\,
            ce => 'H',
            sr => \N__49613\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIOBV3_8_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33701\,
            lcout => \drone_H_disp_front_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33863\,
            in1 => \N__33887\,
            in2 => \N__33839\,
            in3 => \N__33764\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33788\,
            in1 => \N__33809\,
            in2 => \N__33959\,
            in3 => \N__35240\,
            lcout => \reset_module_System.reset6_15\,
            ltout => \reset_module_System.reset6_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__33692\,
            in1 => \N__35211\,
            in2 => \N__33695\,
            in3 => \N__35018\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35055\,
            in2 => \_gnd_net_\,
            in3 => \N__35126\,
            lcout => \reset_module_System.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35125\,
            in2 => \N__35057\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35239\,
            in2 => \_gnd_net_\,
            in3 => \N__33812\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33808\,
            in2 => \_gnd_net_\,
            in3 => \N__33797\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35138\,
            in2 => \_gnd_net_\,
            in3 => \N__33794\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35150\,
            in2 => \_gnd_net_\,
            in3 => \N__33791\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33787\,
            in2 => \_gnd_net_\,
            in3 => \N__33776\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35177\,
            in2 => \_gnd_net_\,
            in3 => \N__33773\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35189\,
            in2 => \_gnd_net_\,
            in3 => \N__33770\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__51481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35164\,
            in2 => \_gnd_net_\,
            in3 => \N__33767\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33760\,
            in2 => \_gnd_net_\,
            in3 => \N__33749\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33883\,
            in2 => \_gnd_net_\,
            in3 => \N__33872\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35068\,
            in2 => \_gnd_net_\,
            in3 => \N__33869\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33899\,
            in2 => \_gnd_net_\,
            in3 => \N__33866\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33859\,
            in2 => \_gnd_net_\,
            in3 => \N__33848\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33923\,
            in2 => \_gnd_net_\,
            in3 => \N__33845\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35090\,
            in2 => \_gnd_net_\,
            in3 => \N__33842\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__51469\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33832\,
            in2 => \_gnd_net_\,
            in3 => \N__33821\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__51454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35104\,
            in2 => \_gnd_net_\,
            in3 => \N__33818\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__51454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33935\,
            in3 => \N__33815\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__51454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33955\,
            in2 => \_gnd_net_\,
            in3 => \N__33941\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__51454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33938\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51454\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33931\,
            in1 => \N__33922\,
            in2 => \N__33911\,
            in3 => \N__33898\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNICBN01_6_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40425\,
            in1 => \N__45140\,
            in2 => \_gnd_net_\,
            in3 => \N__44919\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43375\,
            in1 => \N__37163\,
            in2 => \N__43241\,
            in3 => \N__35405\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51438\,
            ce => 'H',
            sr => \N__49535\
        );

    \ppm_encoder_1.init_pulses_RNIDCN01_0_7_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44920\,
            in1 => \_gnd_net_\,
            in2 => \N__45158\,
            in3 => \N__40962\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__40963\,
            in1 => \N__43871\,
            in2 => \N__45964\,
            in3 => \N__43782\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__43870\,
            in1 => \N__40426\,
            in2 => \N__43784\,
            in3 => \N__38780\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_8_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__43223\,
            in1 => \N__43376\,
            in2 => \N__35396\,
            in3 => \N__37148\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51438\,
            ce => 'H',
            sr => \N__49535\
        );

    \ppm_encoder_1.rudder_10_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__34049\,
            in1 => \N__34022\,
            in2 => \N__41148\,
            in3 => \N__46311\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51424\,
            ce => 'H',
            sr => \N__49544\
        );

    \ppm_encoder_1.init_pulses_6_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43366\,
            in1 => \N__37190\,
            in2 => \N__43238\,
            in3 => \N__35291\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51424\,
            ce => 'H',
            sr => \N__49544\
        );

    \ppm_encoder_1.elevator_0_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__46310\,
            in1 => \N__35735\,
            in2 => \_gnd_net_\,
            in3 => \N__44003\,
            lcout => \ppm_encoder_1.elevatorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51424\,
            ce => 'H',
            sr => \N__49544\
        );

    \ppm_encoder_1.throttle_RNII0PT2_11_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__33999\,
            in1 => \N__35269\,
            in2 => \N__45842\,
            in3 => \N__45933\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIC22D6_11_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__35375\,
            in1 => \_gnd_net_\,
            in2 => \N__34010\,
            in3 => \N__34007\,
            lcout => \ppm_encoder_1.elevator_RNIC22D6Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI24LH2_11_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__33969\,
            in1 => \N__33981\,
            in2 => \N__45368\,
            in3 => \N__45500\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46745\,
            in1 => \N__34000\,
            in2 => \_gnd_net_\,
            in3 => \N__33970\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46589\,
            in2 => \N__33986\,
            in3 => \N__33982\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_11_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__33983\,
            in1 => \N__34231\,
            in2 => \N__46367\,
            in3 => \N__34364\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51410\,
            ce => 'H',
            sr => \N__49549\
        );

    \ppm_encoder_1.elevator_11_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__33971\,
            in1 => \N__46321\,
            in2 => \N__36302\,
            in3 => \N__36335\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51410\,
            ce => 'H',
            sr => \N__49549\
        );

    \ppm_encoder_1.throttle_RNIK2PT2_12_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__34107\,
            in1 => \N__34141\,
            in2 => \N__45935\,
            in3 => \N__45839\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIH72D6_12_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35422\,
            in2 => \N__34118\,
            in3 => \N__34115\,
            lcout => \ppm_encoder_1.elevator_RNIH72D6Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI46LH2_12_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__34065\,
            in1 => \N__45477\,
            in2 => \N__34085\,
            in3 => \N__45366\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34067\,
            in1 => \N__34108\,
            in2 => \_gnd_net_\,
            in3 => \N__46782\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46630\,
            in1 => \_gnd_net_\,
            in2 => \N__34088\,
            in3 => \N__34083\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__34084\,
            in1 => \N__37820\,
            in2 => \N__46307\,
            in3 => \N__34352\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51396\,
            ce => 'H',
            sr => \N__49557\
        );

    \ppm_encoder_1.elevator_12_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__34066\,
            in1 => \N__46244\,
            in2 => \N__36284\,
            in3 => \N__36260\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51396\,
            ce => 'H',
            sr => \N__49557\
        );

    \ppm_encoder_1.un1_aileron_cry_0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46026\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_0_THRU_LUT4_0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35977\,
            in2 => \N__47883\,
            in3 => \N__34052\,
            lcout => \ppm_encoder_1.un1_aileron_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_0\,
            carryout => \ppm_encoder_1.un1_aileron_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_1_THRU_LUT4_0_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35929\,
            in2 => \_gnd_net_\,
            in3 => \N__34169\,
            lcout => \ppm_encoder_1.un1_aileron_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_1\,
            carryout => \ppm_encoder_1.un1_aileron_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_2_THRU_LUT4_0_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38615\,
            in2 => \N__47884\,
            in3 => \N__34166\,
            lcout => \ppm_encoder_1.un1_aileron_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_2\,
            carryout => \ppm_encoder_1.un1_aileron_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_3_THRU_LUT4_0_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46868\,
            in2 => \_gnd_net_\,
            in3 => \N__34163\,
            lcout => \ppm_encoder_1.un1_aileron_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_3\,
            carryout => \ppm_encoder_1.un1_aileron_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_4_THRU_LUT4_0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38579\,
            in2 => \_gnd_net_\,
            in3 => \N__34160\,
            lcout => \ppm_encoder_1.un1_aileron_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_4\,
            carryout => \ppm_encoder_1.un1_aileron_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_5_THRU_LUT4_0_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47842\,
            in2 => \N__38698\,
            in3 => \N__34157\,
            lcout => \ppm_encoder_1.un1_aileron_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_5\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45654\,
            in2 => \_gnd_net_\,
            in3 => \N__34154\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37542\,
            in2 => \_gnd_net_\,
            in3 => \N__34151\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38514\,
            in2 => \_gnd_net_\,
            in3 => \N__34148\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36036\,
            in2 => \_gnd_net_\,
            in3 => \N__34145\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34224\,
            in2 => \_gnd_net_\,
            in3 => \N__34355\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37819\,
            in2 => \_gnd_net_\,
            in3 => \N__34343\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47990\,
            in2 => \N__41621\,
            in3 => \N__34340\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34337\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51369\,
            ce => \N__36697\,
            sr => \N__49575\
        );

    \pid_alt.error_cry_0_c_inv_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__47989\,
            in1 => \N__34273\,
            in2 => \_gnd_net_\,
            in3 => \N__34296\,
            lcout => \pid_alt.drone_altitude_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_10_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__38170\,
            in1 => \N__35886\,
            in2 => \N__36041\,
            in3 => \N__34259\,
            lcout => side_order_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.source_pid_1_11_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__35887\,
            in1 => \N__38171\,
            in2 => \N__34232\,
            in3 => \N__34439\,
            lcout => side_order_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.source_pid_1_6_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__38172\,
            in1 => \N__35888\,
            in2 => \N__38697\,
            in3 => \N__34208\,
            lcout => side_order_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.source_pid_1_7_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__35889\,
            in1 => \N__38173\,
            in2 => \N__45658\,
            in3 => \N__34406\,
            lcout => side_order_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.source_pid_1_8_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__38174\,
            in1 => \N__35890\,
            in2 => \N__37552\,
            in3 => \N__34601\,
            lcout => side_order_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.source_pid_1_9_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__35891\,
            in1 => \N__38175\,
            in2 => \N__38524\,
            in3 => \N__34568\,
            lcout => side_order_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51357\,
            ce => 'H',
            sr => \N__38073\
        );

    \pid_side.state_RNI34HSI_1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35885\,
            in2 => \_gnd_net_\,
            in3 => \N__38060\,
            lcout => \pid_side.state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNIOB8E3_2_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34664\,
            in1 => \N__35896\,
            in2 => \N__34655\,
            in3 => \N__35956\,
            lcout => \pid_side.un1_reset_i_a5_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIH97T2_21_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38361\,
            in1 => \N__36007\,
            in2 => \_gnd_net_\,
            in3 => \N__38302\,
            lcout => \pid_side.N_534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34472\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNILTAI1_0_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38246\,
            in1 => \N__35783\,
            in2 => \N__38147\,
            in3 => \N__41919\,
            lcout => \pid_side.un1_reset_i_a5_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNITODS2_7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__34432\,
            in1 => \N__34402\,
            in2 => \N__38314\,
            in3 => \N__34376\,
            lcout => \pid_side.un1_reset_i_a5_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50072\,
            lcout => \pid_front.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51339\,
            ce => \N__48481\,
            sr => \N__49598\
        );

    \pid_side.pid_prereg_RNI7QS63_14_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34805\,
            in1 => \N__34789\,
            in2 => \N__34772\,
            in3 => \N__34757\,
            lcout => \pid_side.N_563\,
            ltout => \pid_side.N_563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNIGPS29_1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34739\,
            in1 => \N__34721\,
            in2 => \N__34733\,
            in3 => \N__34730\,
            lcout => OPEN,
            ltout => \pid_side.N_311_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNIQG8J9_21_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__38360\,
            in1 => \N__35878\,
            in2 => \N__34724\,
            in3 => \N__49023\,
            lcout => \pid_side.un1_reset_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNIN87D1_1_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37842\,
            in1 => \N__35948\,
            in2 => \N__35877\,
            in3 => \N__49831\,
            lcout => \pid_side.un1_reset_i_a5_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__50019\,
            in1 => \N__34715\,
            in2 => \N__34682\,
            in3 => \N__35949\,
            lcout => \pid_side.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51333\,
            ce => 'H',
            sr => \N__49602\
        );

    \pid_side.pid_prereg_RNI2JR61_1_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__38138\,
            in1 => \N__38315\,
            in2 => \_gnd_net_\,
            in3 => \N__49830\,
            lcout => \pid_side.un1_reset_i_a5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_RNI39UK1_0_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35788\,
            in1 => \N__41920\,
            in2 => \N__38258\,
            in3 => \N__37843\,
            lcout => \pid_side.un1_reset_i_a5_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_RNI3CC11_14_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__36356\,
            in1 => \N__34609\,
            in2 => \N__34961\,
            in3 => \N__36416\,
            lcout => \pid_front.N_569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_14_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__50543\,
            in1 => \N__47768\,
            in2 => \N__42817\,
            in3 => \N__34610\,
            lcout => \pid_front.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51325\,
            ce => 'H',
            sr => \N__49606\
        );

    \pid_front.pid_prereg_RNID03J_17_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34951\,
            in1 => \N__36532\,
            in2 => \N__34940\,
            in3 => \N__36544\,
            lcout => \pid_front.m7_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_9_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__36092\,
            in1 => \N__36062\,
            in2 => \N__46397\,
            in3 => \N__35695\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \N__49614\
        );

    \pid_front.pid_prereg_18_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42800\,
            in1 => \N__48590\,
            in2 => \N__50264\,
            in3 => \N__34952\,
            lcout => \pid_front.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \N__49614\
        );

    \pid_front.pid_prereg_19_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42801\,
            in1 => \N__48575\,
            in2 => \N__51911\,
            in3 => \N__34939\,
            lcout => \pid_front.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \N__49614\
        );

    \pid_front.pid_prereg_9_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__47591\,
            in1 => \N__48743\,
            in2 => \N__34923\,
            in3 => \N__42776\,
            lcout => \pid_front.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51312\,
            ce => 'H',
            sr => \N__49617\
        );

    \pid_front.pid_prereg_11_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__51797\,
            in1 => \N__48251\,
            in2 => \N__42805\,
            in3 => \N__34884\,
            lcout => \pid_front.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51312\,
            ce => 'H',
            sr => \N__49617\
        );

    \pid_front.pid_prereg_13_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__51863\,
            in1 => \N__47783\,
            in2 => \N__34841\,
            in3 => \N__42775\,
            lcout => \pid_front.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51312\,
            ce => 'H',
            sr => \N__49617\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_15_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36620\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \drone_H_disp_front_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51308\,
            ce => \N__48354\,
            sr => \N__49620\
        );

    \reset_module_System.reset_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__35223\,
            in1 => \N__35207\,
            in2 => \_gnd_net_\,
            in3 => \N__35015\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__35212\,
            in1 => \N__35246\,
            in2 => \N__35228\,
            in3 => \N__35017\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__35016\,
            in1 => \N__35224\,
            in2 => \N__35213\,
            in3 => \N__35056\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35188\,
            in1 => \N__35176\,
            in2 => \N__35165\,
            in3 => \N__35149\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35137\,
            in2 => \_gnd_net_\,
            in3 => \N__35124\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35108\,
            in1 => \N__35089\,
            in2 => \N__35078\,
            in3 => \N__35075\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__35069\,
            in1 => \N__35054\,
            in2 => \N__35030\,
            in3 => \N__35027\,
            lcout => \reset_module_System.reset6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_9_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__35000\,
            in1 => \N__34985\,
            in2 => \N__46390\,
            in3 => \N__35664\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51482\,
            ce => 'H',
            sr => \N__49529\
        );

    \ppm_encoder_1.init_pulses_11_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__43353\,
            in1 => \N__43237\,
            in2 => \N__37286\,
            in3 => \N__35348\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51470\,
            ce => 'H',
            sr => \N__49536\
        );

    \ppm_encoder_1.init_pulses_RNIOTJT_11_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__35283\,
            in1 => \N__45144\,
            in2 => \_gnd_net_\,
            in3 => \N__44931\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIOTJT_0_11_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44932\,
            in1 => \_gnd_net_\,
            in2 => \N__45159\,
            in3 => \N__35284\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35285\,
            in1 => \N__43753\,
            in2 => \_gnd_net_\,
            in3 => \N__35273\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41203\,
            in2 => \N__35249\,
            in3 => \N__43869\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_12_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__43236\,
            in1 => \N__43354\,
            in2 => \N__37274\,
            in3 => \N__35330\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51470\,
            ce => 'H',
            sr => \N__49536\
        );

    \ppm_encoder_1.init_pulses_16_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43350\,
            in1 => \N__37247\,
            in2 => \N__43242\,
            in3 => \N__35471\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51455\,
            ce => 'H',
            sr => \N__49545\
        );

    \ppm_encoder_1.init_pulses_RNIT2KT_16_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__45180\,
            in1 => \N__45136\,
            in2 => \_gnd_net_\,
            in3 => \N__44917\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_17_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43351\,
            in1 => \N__37232\,
            in2 => \N__43243\,
            in3 => \N__35447\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51455\,
            ce => 'H',
            sr => \N__49545\
        );

    \ppm_encoder_1.init_pulses_RNIU3KT_0_17_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__44244\,
            in1 => \N__45135\,
            in2 => \_gnd_net_\,
            in3 => \N__44916\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIU3KT_17_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44918\,
            in1 => \_gnd_net_\,
            in2 => \N__45157\,
            in3 => \N__44245\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_18_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__43221\,
            in1 => \N__37220\,
            in2 => \N__43373\,
            in3 => \N__35432\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51455\,
            ce => 'H',
            sr => \N__49545\
        );

    \ppm_encoder_1.init_pulses_2_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__43352\,
            in1 => \N__43222\,
            in2 => \N__37214\,
            in3 => \N__35309\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51455\,
            ce => 'H',
            sr => \N__49545\
        );

    \ppm_encoder_1.init_pulses_RNI87N01_2_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40911\,
            in1 => \N__45134\,
            in2 => \_gnd_net_\,
            in3 => \N__44915\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNINSH16_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42045\,
            in2 => \N__37655\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37921\,
            in2 => \N__37910\,
            in3 => \N__35312\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37687\,
            in2 => \N__37673\,
            in3 => \N__35303\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41996\,
            in2 => \N__41939\,
            in3 => \N__35300\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40789\,
            in2 => \N__38033\,
            in3 => \N__35297\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44122\,
            in2 => \N__37982\,
            in3 => \N__35294\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38743\,
            in2 => \N__38723\,
            in3 => \N__35408\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45727\,
            in2 => \N__45707\,
            in3 => \N__35399\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44077\,
            in2 => \N__37571\,
            in3 => \N__35384\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44146\,
            in2 => \N__35486\,
            in3 => \N__35381\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35587\,
            in2 => \N__35573\,
            in3 => \N__35378\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35371\,
            in2 => \N__35357\,
            in3 => \N__35339\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35336\,
            in2 => \N__35423\,
            in3 => \N__35321\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41659\,
            in2 => \N__41645\,
            in3 => \N__35318\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41851\,
            in2 => \N__41837\,
            in3 => \N__35315\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37409\,
            in2 => \N__37361\,
            in3 => \N__35474\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44597\,
            in2 => \_gnd_net_\,
            in3 => \N__35462\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35459\,
            in3 => \N__35438\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__40859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35435\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_1_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46795\,
            in1 => \N__37947\,
            in2 => \_gnd_net_\,
            in3 => \N__37893\,
            lcout => \ppm_encoder_1.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNINSJT_10_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41166\,
            in1 => \N__45148\,
            in2 => \_gnd_net_\,
            in3 => \N__44909\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPUJT_12_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44910\,
            in1 => \_gnd_net_\,
            in2 => \N__45160\,
            in3 => \N__40887\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR0KT_14_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__37445\,
            in1 => \N__45152\,
            in2 => \_gnd_net_\,
            in3 => \N__44911\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__43881\,
            in1 => \N__44105\,
            in2 => \N__37613\,
            in3 => \N__43728\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46663\,
            in1 => \N__35546\,
            in2 => \_gnd_net_\,
            in3 => \N__37966\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_1_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37967\,
            in1 => \N__35540\,
            in2 => \N__46308\,
            in3 => \N__35978\,
            lcout => \ppm_encoder_1.aileronZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51397\,
            ce => 'H',
            sr => \N__49576\
        );

    \ppm_encoder_1.elevator_1_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__36167\,
            in1 => \N__36197\,
            in2 => \N__37952\,
            in3 => \N__46255\,
            lcout => \ppm_encoder_1.elevatorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51397\,
            ce => 'H',
            sr => \N__49576\
        );

    \ppm_encoder_1.throttle_1_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__35534\,
            in1 => \N__35522\,
            in2 => \N__46309\,
            in3 => \N__37894\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51397\,
            ce => 'H',
            sr => \N__49576\
        );

    \ppm_encoder_1.aileron_2_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__37714\,
            in1 => \N__46248\,
            in2 => \N__35930\,
            in3 => \N__35495\,
            lcout => \ppm_encoder_1.aileronZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51397\,
            ce => 'H',
            sr => \N__49576\
        );

    \ppm_encoder_1.elevator_RNIGN7O2_9_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__35701\,
            in1 => \N__38485\,
            in2 => \N__45498\,
            in3 => \N__45367\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIV9PO6_9_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__44150\,
            in1 => \_gnd_net_\,
            in2 => \N__35489\,
            in3 => \N__35627\,
            lcout => \ppm_encoder_1.throttle_RNIV9PO6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46665\,
            in1 => \N__35681\,
            in2 => \_gnd_net_\,
            in3 => \N__38486\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35648\,
            in1 => \N__46807\,
            in2 => \_gnd_net_\,
            in3 => \N__35702\,
            lcout => \ppm_encoder_1.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__35666\,
            in1 => \N__43711\,
            in2 => \N__43886\,
            in3 => \N__44177\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__44498\,
            in1 => \_gnd_net_\,
            in2 => \N__35675\,
            in3 => \N__35672\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51382\,
            ce => \N__44410\,
            sr => \N__49584\
        );

    \ppm_encoder_1.throttle_RNI04QV2_9_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__35665\,
            in1 => \N__35647\,
            in2 => \N__45832\,
            in3 => \N__45897\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__43710\,
            in1 => \N__43882\,
            in2 => \_gnd_net_\,
            in3 => \N__41416\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGUOT2_10_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__35620\,
            in1 => \N__41149\,
            in2 => \N__45841\,
            in3 => \N__45905\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI7T1D6_10_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35594\,
            in2 => \N__35576\,
            in3 => \N__35561\,
            lcout => \ppm_encoder_1.elevator_RNI7T1D6Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI02LH2_10_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__38424\,
            in1 => \N__36018\,
            in2 => \N__45494\,
            in3 => \N__45353\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46664\,
            in1 => \N__35555\,
            in2 => \_gnd_net_\,
            in3 => \N__36019\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_10_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__36020\,
            in1 => \N__46256\,
            in2 => \N__36050\,
            in3 => \N__36037\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51370\,
            ce => 'H',
            sr => \N__49593\
        );

    \pid_side.pid_prereg_esr_RNIAA5MI_21_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__38389\,
            in1 => \N__36008\,
            in2 => \N__35993\,
            in3 => \N__35984\,
            lcout => \pid_side.pid_prereg_esr_RNIAA5MIZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__35747\,
            in1 => \N__35892\,
            in2 => \N__46030\,
            in3 => \N__41921\,
            lcout => side_order_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51358\,
            ce => 'H',
            sr => \N__38075\
        );

    \pid_side.source_pid_1_1_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35893\,
            in1 => \N__35748\,
            in2 => \N__49835\,
            in3 => \N__35976\,
            lcout => side_order_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51358\,
            ce => 'H',
            sr => \N__38075\
        );

    \pid_side.source_pid_1_2_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__35749\,
            in1 => \N__35894\,
            in2 => \N__35928\,
            in3 => \N__35957\,
            lcout => side_order_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51358\,
            ce => 'H',
            sr => \N__38075\
        );

    \pid_side.source_pid_1_3_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35895\,
            in1 => \N__35750\,
            in2 => \N__35792\,
            in3 => \N__38614\,
            lcout => side_order_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51358\,
            ce => 'H',
            sr => \N__38075\
        );

    \pid_side.pid_prereg_esr_RNIIK254_21_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__38388\,
            in1 => \N__38316\,
            in2 => \N__38370\,
            in3 => \N__37855\,
            lcout => \pid_side.N_291\,
            ltout => \pid_side.N_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_RNISEFQ7_4_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__38256\,
            in1 => \N__38123\,
            in2 => \N__35753\,
            in3 => \N__38191\,
            lcout => \pid_side.N_451_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_0_c_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35727\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_0_THRU_LUT4_0_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36192\,
            in2 => \N__48084\,
            in3 => \N__36158\,
            lcout => \ppm_encoder_1.un1_elevator_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_0\,
            carryout => \ppm_encoder_1.un1_elevator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_1_THRU_LUT4_0_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39246\,
            in2 => \_gnd_net_\,
            in3 => \N__36155\,
            lcout => \ppm_encoder_1.un1_elevator_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_1\,
            carryout => \ppm_encoder_1.un1_elevator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_2_THRU_LUT4_0_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36148\,
            in2 => \N__48085\,
            in3 => \N__36110\,
            lcout => \ppm_encoder_1.un1_elevator_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_2\,
            carryout => \ppm_encoder_1.un1_elevator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_3_THRU_LUT4_0_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46831\,
            in2 => \_gnd_net_\,
            in3 => \N__36107\,
            lcout => \ppm_encoder_1.un1_elevator_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_3\,
            carryout => \ppm_encoder_1.un1_elevator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_4_THRU_LUT4_0_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39127\,
            in2 => \_gnd_net_\,
            in3 => \N__36104\,
            lcout => \ppm_encoder_1.un1_elevator_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_4\,
            carryout => \ppm_encoder_1.un1_elevator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_5_THRU_LUT4_0_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39172\,
            in2 => \N__48086\,
            in3 => \N__36101\,
            lcout => \ppm_encoder_1.un1_elevator_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_5\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45597\,
            in2 => \_gnd_net_\,
            in3 => \N__36098\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37498\,
            in2 => \_gnd_net_\,
            in3 => \N__36095\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36091\,
            in2 => \_gnd_net_\,
            in3 => \N__36341\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38464\,
            in2 => \_gnd_net_\,
            in3 => \N__36338\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36334\,
            in2 => \_gnd_net_\,
            in3 => \N__36287\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36277\,
            in2 => \_gnd_net_\,
            in3 => \N__36245\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41560\,
            in2 => \N__48087\,
            in3 => \N__36242\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36239\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51340\,
            ce => \N__36692\,
            sr => \N__49607\
        );

    \pid_front.pid_prereg_esr_RNI5QBD_0_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38955\,
            in1 => \N__38886\,
            in2 => \N__38925\,
            in3 => \N__36231\,
            lcout => \pid_front.un1_reset_i_a5_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_4_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36970\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51326\,
            ce => \N__42526\,
            sr => \N__49615\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_5_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36880\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51326\,
            ce => \N__42526\,
            sr => \N__49615\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_6_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48448\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51326\,
            ce => \N__42526\,
            sr => \N__49615\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_7_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36605\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51326\,
            ce => \N__42526\,
            sr => \N__49615\
        );

    \pid_front.pid_prereg_17_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__42791\,
            in1 => \N__47729\,
            in2 => \N__36548\,
            in3 => \N__51569\,
            lcout => \pid_front.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51319\,
            ce => 'H',
            sr => \N__49618\
        );

    \pid_front.pid_prereg_20_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42798\,
            in1 => \N__48560\,
            in2 => \N__51722\,
            in3 => \N__36533\,
            lcout => \pid_front.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51319\,
            ce => 'H',
            sr => \N__49618\
        );

    \pid_front.pid_prereg_7_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__42799\,
            in1 => \N__50417\,
            in2 => \N__36516\,
            in3 => \N__47612\,
            lcout => \pid_front.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51319\,
            ce => 'H',
            sr => \N__49618\
        );

    \pid_front.pid_prereg_6_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__47627\,
            in1 => \N__50312\,
            in2 => \N__42816\,
            in3 => \N__36477\,
            lcout => \pid_front.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51319\,
            ce => 'H',
            sr => \N__49618\
        );

    \pid_front.pid_prereg_12_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__51767\,
            in1 => \N__47798\,
            in2 => \N__42815\,
            in3 => \N__36440\,
            lcout => \pid_front.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51319\,
            ce => 'H',
            sr => \N__49618\
        );

    \pid_front.pid_prereg_16_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__47741\,
            in1 => \N__50345\,
            in2 => \N__42804\,
            in3 => \N__36415\,
            lcout => \pid_front.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51316\,
            ce => 'H',
            sr => \N__49621\
        );

    \pid_front.pid_prereg_2_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42764\,
            in1 => \N__48709\,
            in2 => \N__47699\,
            in3 => \N__36386\,
            lcout => \pid_front.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51316\,
            ce => 'H',
            sr => \N__49621\
        );

    \pid_front.pid_prereg_15_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__47753\,
            in1 => \N__51827\,
            in2 => \N__42803\,
            in3 => \N__36355\,
            lcout => \pid_front.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51316\,
            ce => 'H',
            sr => \N__49621\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_10_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37129\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51313\,
            ce => \N__48355\,
            sr => \N__49623\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_11_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37048\,
            lcout => \drone_H_disp_front_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51313\,
            ce => \N__48355\,
            sr => \N__49623\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_12_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36971\,
            lcout => \drone_H_disp_front_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51313\,
            ce => \N__48355\,
            sr => \N__49623\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_13_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36884\,
            lcout => \drone_H_disp_front_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51313\,
            ce => \N__48355\,
            sr => \N__49623\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_9_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36809\,
            lcout => \dron_frame_decoder_1.drone_H_disp_front_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51313\,
            ce => \N__48355\,
            sr => \N__49623\
        );

    \ppm_encoder_1.rudder_esr_4_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36731\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51503\,
            ce => \N__36688\,
            sr => \N__49530\
        );

    \ppm_encoder_1.rudder_esr_5_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36713\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51503\,
            ce => \N__36688\,
            sr => \N__49530\
        );

    \ppm_encoder_1.init_pulses_RNI4Q625_0_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41288\,
            in2 => \N__37346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37388\,
            in2 => \_gnd_net_\,
            in3 => \N__36635\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40484\,
            in2 => \N__40442\,
            in3 => \N__37202\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40826\,
            in3 => \N__37199\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40769\,
            in2 => \_gnd_net_\,
            in3 => \N__37196\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40478\,
            in2 => \_gnd_net_\,
            in3 => \N__37193\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40490\,
            in2 => \N__40412\,
            in3 => \N__37178\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37175\,
            in2 => \_gnd_net_\,
            in3 => \N__37151\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37376\,
            in2 => \_gnd_net_\,
            in3 => \N__37136\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37370\,
            in3 => \N__37133\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37622\,
            in2 => \_gnd_net_\,
            in3 => \N__37295\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37292\,
            in2 => \_gnd_net_\,
            in3 => \N__37277\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40865\,
            in2 => \_gnd_net_\,
            in3 => \N__37265\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40496\,
            in2 => \N__40451\,
            in3 => \N__37262\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37304\,
            in2 => \_gnd_net_\,
            in3 => \N__37259\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44054\,
            in2 => \_gnd_net_\,
            in3 => \N__37256\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37253\,
            in2 => \_gnd_net_\,
            in3 => \N__37241\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37238\,
            in2 => \_gnd_net_\,
            in3 => \N__37226\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__45240\,
            in1 => \N__44835\,
            in2 => \N__45133\,
            in3 => \N__37223\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIEDN01_0_8_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44833\,
            in1 => \_gnd_net_\,
            in2 => \N__45089\,
            in3 => \N__44101\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFEN01_0_9_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__44170\,
            in1 => \N__45028\,
            in2 => \_gnd_net_\,
            in3 => \N__44834\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI1AEO1_15_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__45029\,
            in1 => \N__44202\,
            in2 => \N__44912\,
            in3 => \N__41443\,
            lcout => \ppm_encoder_1.init_pulses_RNI1AEO1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_0_3_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45024\,
            in2 => \_gnd_net_\,
            in3 => \N__44832\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNILVE13_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__44839\,
            in1 => \N__41409\,
            in2 => \N__37349\,
            in3 => \N__41345\,
            lcout => \ppm_encoder_1.init_pulses_RNILVE13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43358\,
            in1 => \N__37334\,
            in2 => \N__43239\,
            in3 => \N__37325\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51456\,
            ce => 'H',
            sr => \N__49558\
        );

    \ppm_encoder_1.init_pulses_RNIQVJT_13_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__40464\,
            in1 => \_gnd_net_\,
            in2 => \N__45131\,
            in3 => \N__44899\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_14_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43359\,
            in1 => \N__37319\,
            in2 => \N__43240\,
            in3 => \N__37310\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51456\,
            ce => 'H',
            sr => \N__49558\
        );

    \ppm_encoder_1.init_pulses_RNIR0KT_0_14_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__44898\,
            in1 => \N__45078\,
            in2 => \_gnd_net_\,
            in3 => \N__37440\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__37441\,
            in1 => \N__43757\,
            in2 => \N__43852\,
            in3 => \N__41467\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__41693\,
            in1 => \N__43835\,
            in2 => \N__43776\,
            in3 => \N__40465\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__43175\,
            in1 => \N__37424\,
            in2 => \N__43374\,
            in3 => \N__37415\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51456\,
            ce => 'H',
            sr => \N__49558\
        );

    \ppm_encoder_1.init_pulses_0_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__43176\,
            in1 => \N__42032\,
            in2 => \N__41381\,
            in3 => \N__43361\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51439\,
            ce => 'H',
            sr => \N__49566\
        );

    \ppm_encoder_1.init_pulses_RNI65N01_0_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41405\,
            in1 => \N__45052\,
            in2 => \_gnd_net_\,
            in3 => \N__44858\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQ_3_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__44861\,
            in1 => \_gnd_net_\,
            in2 => \N__45122\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI58QQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_1_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43360\,
            in1 => \N__37403\,
            in2 => \N__43220\,
            in3 => \N__37394\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51439\,
            ce => 'H',
            sr => \N__49566\
        );

    \ppm_encoder_1.init_pulses_RNI76N01_1_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44859\,
            in1 => \_gnd_net_\,
            in2 => \N__45121\,
            in3 => \N__40941\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI76N01_0_1_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40942\,
            in1 => \N__45051\,
            in2 => \_gnd_net_\,
            in3 => \N__44857\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__43177\,
            in1 => \N__37640\,
            in2 => \N__37631\,
            in3 => \N__43362\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51439\,
            ce => 'H',
            sr => \N__49566\
        );

    \ppm_encoder_1.init_pulses_RNINSJT_0_10_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41167\,
            in1 => \N__45056\,
            in2 => \_gnd_net_\,
            in3 => \N__44860\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIU1QV2_8_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__37755\,
            in1 => \N__37606\,
            in2 => \N__45932\,
            in3 => \N__45829\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIQ4PO6_8_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44078\,
            in2 => \N__37574\,
            in3 => \N__37562\,
            lcout => \ppm_encoder_1.throttle_RNIQ4PO6Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIEL7O2_8_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__37458\,
            in1 => \N__37512\,
            in2 => \N__45361\,
            in3 => \N__45476\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__37460\,
            in1 => \N__37756\,
            in2 => \N__46813\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46601\,
            in2 => \N__37556\,
            in3 => \N__37513\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_8_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__37514\,
            in1 => \N__37553\,
            in2 => \N__46387\,
            in3 => \N__37526\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51425\,
            ce => 'H',
            sr => \N__49577\
        );

    \ppm_encoder_1.elevator_8_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__37459\,
            in1 => \N__37502\,
            in2 => \N__46396\,
            in3 => \N__37472\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51425\,
            ce => 'H',
            sr => \N__49577\
        );

    \ppm_encoder_1.throttle_8_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__37799\,
            in1 => \N__37757\,
            in2 => \N__37769\,
            in3 => \N__46386\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51425\,
            ce => 'H',
            sr => \N__49577\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111011100"
        )
    port map (
            in0 => \N__45156\,
            in1 => \N__49784\,
            in2 => \N__44930\,
            in3 => \N__41723\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110000000"
        )
    port map (
            in0 => \N__43701\,
            in1 => \N__46806\,
            in2 => \N__46662\,
            in3 => \N__41261\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__41262\,
            in1 => \N__49783\,
            in2 => \N__37745\,
            in3 => \N__44786\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__46642\,
            in1 => \N__44900\,
            in2 => \N__49797\,
            in3 => \N__41746\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIKGMK2_2_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37742\,
            in1 => \N__37710\,
            in2 => \N__45360\,
            in3 => \N__45802\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIPVQ05_2_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001111"
        )
    port map (
            in0 => \N__37694\,
            in1 => \N__39207\,
            in2 => \N__37676\,
            in3 => \N__45454\,
            lcout => \ppm_encoder_1.elevator_RNIPVQ05Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__37661\,
            in1 => \N__49785\,
            in2 => \N__40993\,
            in3 => \N__44787\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIHNQ05_0_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__44011\,
            in1 => \N__45453\,
            in2 => \N__42059\,
            in3 => \N__41699\,
            lcout => \ppm_encoder_1.elevator_RNIHNQ05Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41720\,
            in2 => \_gnd_net_\,
            in3 => \N__41741\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__44668\,
            in1 => \N__41113\,
            in2 => \N__43739\,
            in3 => \N__49015\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI077O2_1_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__37965\,
            in1 => \N__45314\,
            in2 => \N__37951\,
            in3 => \N__45440\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIUINC6_1_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101111"
        )
    port map (
            in0 => \N__45890\,
            in1 => \N__37871\,
            in2 => \N__37928\,
            in3 => \N__37925\,
            lcout => \ppm_encoder_1.throttle_RNIUINC6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__37865\,
            in1 => \N__49014\,
            in2 => \N__41117\,
            in3 => \N__44669\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7D_0_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__41721\,
            in1 => \_gnd_net_\,
            in2 => \N__41747\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHO7DZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEES71_1_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37895\,
            in1 => \N__42175\,
            in2 => \N__37874\,
            in3 => \N__44667\,
            lcout => \ppm_encoder_1.throttle_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_2_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37864\,
            in2 => \_gnd_net_\,
            in3 => \N__40983\,
            lcout => \ppm_encoder_1.N_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.source_pid_1_esr_12_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__38318\,
            in1 => \N__38398\,
            in2 => \N__38375\,
            in3 => \N__37856\,
            lcout => side_order_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51383\,
            ce => \N__38090\,
            sr => \N__38074\
        );

    \pid_side.source_pid_1_esr_13_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__38399\,
            in1 => \N__38371\,
            in2 => \_gnd_net_\,
            in3 => \N__38317\,
            lcout => side_order_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51383\,
            ce => \N__38090\,
            sr => \N__38074\
        );

    \pid_side.source_pid_1_esr_4_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__38142\,
            in1 => \N__38200\,
            in2 => \N__38180\,
            in3 => \N__38257\,
            lcout => side_order_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51383\,
            ce => \N__38090\,
            sr => \N__38074\
        );

    \pid_side.source_pid_1_esr_5_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__38201\,
            in1 => \N__38179\,
            in2 => \_gnd_net_\,
            in3 => \N__38143\,
            lcout => side_order_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51383\,
            ce => \N__38090\,
            sr => \N__38074\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNI9NSB1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41263\,
            in1 => \N__41087\,
            in2 => \N__41367\,
            in3 => \N__44666\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIVRTU2_4_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__45785\,
            in1 => \N__46415\,
            in2 => \N__38039\,
            in3 => \N__41041\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFISN6_4_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40793\,
            in2 => \N__38036\,
            in3 => \N__46889\,
            lcout => \ppm_encoder_1.elevator_RNIFISN6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNI1UTU2_5_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__38018\,
            in1 => \N__43642\,
            in2 => \N__45813\,
            in3 => \N__45889\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8F7O2_5_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__39087\,
            in1 => \N__45423\,
            in2 => \N__38550\,
            in3 => \N__45310\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKNSN6_5_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44126\,
            in2 => \N__37991\,
            in3 => \N__37988\,
            lcout => \ppm_encoder_1.elevator_RNIKNSN6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIQTPV2_6_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__38807\,
            in1 => \N__38776\,
            in2 => \N__45840\,
            in3 => \N__45898\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGQOO6_6_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38750\,
            in2 => \N__38726\,
            in3 => \N__38708\,
            lcout => \ppm_encoder_1.throttle_RNIGQOO6Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAH7O2_6_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__39144\,
            in1 => \N__45422\,
            in2 => \N__38653\,
            in3 => \N__45309\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__38652\,
            in1 => \N__46328\,
            in2 => \N__38702\,
            in3 => \N__38669\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51371\,
            ce => 'H',
            sr => \N__49603\
        );

    \ppm_encoder_1.aileron_3_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__38630\,
            in1 => \N__38613\,
            in2 => \N__46374\,
            in3 => \N__42277\,
            lcout => \ppm_encoder_1.aileronZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.aileron_5_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__38594\,
            in1 => \N__38578\,
            in2 => \N__38554\,
            in3 => \N__46340\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.aileron_9_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__38525\,
            in1 => \N__38498\,
            in2 => \N__46375\,
            in3 => \N__38479\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.elevator_10_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__38460\,
            in1 => \N__38435\,
            in2 => \N__38428\,
            in3 => \N__46341\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.elevator_2_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__46332\,
            in1 => \N__39251\,
            in2 => \N__39215\,
            in3 => \N__39221\,
            lcout => \ppm_encoder_1.elevatorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.elevator_6_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__39185\,
            in1 => \N__39148\,
            in2 => \N__39179\,
            in3 => \N__46342\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \ppm_encoder_1.elevator_5_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__46333\,
            in1 => \N__39128\,
            in2 => \N__39097\,
            in3 => \N__39104\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51359\,
            ce => 'H',
            sr => \N__49608\
        );

    \Commands_frame_decoder.source_xy_kp_1_e_0_4_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40255\,
            in2 => \_gnd_net_\,
            in3 => \N__50797\,
            lcout => xy_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51349\,
            ce => \N__39032\,
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_4_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42814\,
            in1 => \N__48626\,
            in2 => \N__47663\,
            in3 => \N__38961\,
            lcout => \pid_front.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51341\,
            ce => 'H',
            sr => \N__49616\
        );

    \pid_front.pid_prereg_5_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__42810\,
            in1 => \N__48671\,
            in2 => \N__47645\,
            in3 => \N__38924\,
            lcout => \pid_front.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51334\,
            ce => 'H',
            sr => \N__49619\
        );

    \pid_front.pid_prereg_3_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__42809\,
            in1 => \N__50384\,
            in2 => \N__47681\,
            in3 => \N__38892\,
            lcout => \pid_front.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51334\,
            ce => 'H',
            sr => \N__49619\
        );

    \Commands_frame_decoder.source_alt_ki_6_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40139\,
            in2 => \_gnd_net_\,
            in3 => \N__50796\,
            lcout => alt_ki_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51327\,
            ce => \N__38855\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI4D23_13_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43468\,
            lcout => \drone_H_disp_front_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIK7V3_4_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39794\,
            lcout => \drone_H_disp_front_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIL8V3_5_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39788\,
            lcout => \drone_H_disp_front_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIM9V3_6_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39782\,
            lcout => \drone_H_disp_front_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNINAV3_7_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39776\,
            lcout => \drone_H_disp_front_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH3data_esr_0_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39760\,
            lcout => front_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_1_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39651\,
            lcout => front_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_2_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39512\,
            lcout => front_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_3_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39363\,
            lcout => front_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_4_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40403\,
            lcout => front_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_5_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40256\,
            lcout => front_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_esr_6_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40140\,
            lcout => front_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \Commands_frame_decoder.source_CH3data_ess_7_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39993\,
            lcout => front_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51320\,
            ce => \N__39884\,
            sr => \N__49624\
        );

    \pid_front.error_axb_7_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__39853\,
            in1 => \N__39844\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pid_front.error_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI1A23_10_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39866\,
            lcout => \drone_H_disp_front_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNIPCV3_9_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39860\,
            lcout => \drone_H_disp_front_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_axb_8_l_ofx_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__39854\,
            in1 => \N__39845\,
            in2 => \_gnd_net_\,
            in3 => \N__43518\,
            lcout => \pid_front.error_axb_8_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_6_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39836\,
            in1 => \N__40707\,
            in2 => \N__39811\,
            in3 => \N__40759\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51504\,
            ce => 'H',
            sr => \N__40532\
        );

    \uart_pc.data_Aux_7_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__40760\,
            in1 => \N__40543\,
            in2 => \N__40712\,
            in3 => \N__40589\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51504\,
            ce => 'H',
            sr => \N__40532\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__44926\,
            in1 => \_gnd_net_\,
            in2 => \N__41344\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQNZ0Z02\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_0_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41337\,
            in2 => \_gnd_net_\,
            in3 => \N__44925\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41372\,
            in2 => \_gnd_net_\,
            in3 => \N__42182\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_1_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41325\,
            in2 => \_gnd_net_\,
            in3 => \N__44848\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBAN01_0_5_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__44849\,
            in1 => \N__43903\,
            in2 => \_gnd_net_\,
            in3 => \N__45124\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9QBU2_13_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__41441\,
            in1 => \N__41326\,
            in2 => \N__40472\,
            in3 => \N__44853\,
            lcout => \ppm_encoder_1.init_pulses_RNI9QBU2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIN1F13_2_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__41327\,
            in1 => \N__40924\,
            in2 => \N__44913\,
            in3 => \N__41439\,
            lcout => \ppm_encoder_1.init_pulses_RNIN1F13Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIR5F13_6_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41440\,
            in1 => \N__41328\,
            in2 => \N__44933\,
            in3 => \N__40433\,
            lcout => \ppm_encoder_1.init_pulses_RNIR5F13Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011011110"
        )
    port map (
            in0 => \N__44852\,
            in1 => \N__49782\,
            in2 => \N__46582\,
            in3 => \N__45127\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPUJT_0_12_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__45125\,
            in1 => \N__40888\,
            in2 => \_gnd_net_\,
            in3 => \N__44850\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__44851\,
            in1 => \N__41442\,
            in2 => \N__45253\,
            in3 => \N__45126\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_3_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43308\,
            in1 => \N__40847\,
            in2 => \N__43219\,
            in3 => \N__40838\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51483\,
            ce => 'H',
            sr => \N__49559\
        );

    \ppm_encoder_1.init_pulses_RNI98N01_0_3_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110001101100"
        )
    port map (
            in0 => \N__44842\,
            in1 => \N__41221\,
            in2 => \N__45090\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI98N01_3_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41220\,
            in1 => \N__45031\,
            in2 => \_gnd_net_\,
            in3 => \N__44841\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_4_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__40814\,
            in1 => \N__40802\,
            in2 => \N__43244\,
            in3 => \N__43309\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51483\,
            ce => 'H',
            sr => \N__49559\
        );

    \ppm_encoder_1.init_pulses_RNIA9N01_4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__41052\,
            in1 => \N__45030\,
            in2 => \_gnd_net_\,
            in3 => \N__44840\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIA9N01_0_4_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44843\,
            in1 => \_gnd_net_\,
            in2 => \N__45091\,
            in3 => \N__41053\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__41054\,
            in1 => \N__43839\,
            in2 => \N__43783\,
            in3 => \N__41042\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_5_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__41018\,
            in1 => \N__43178\,
            in2 => \N__41006\,
            in3 => \N__43310\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51483\,
            ce => 'H',
            sr => \N__49559\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__46752\,
            in1 => \N__41270\,
            in2 => \_gnd_net_\,
            in3 => \N__42219\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI63RK_3_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41077\,
            in2 => \_gnd_net_\,
            in3 => \N__40994\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDCN01_7_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40967\,
            in2 => \N__40946\,
            in3 => \N__44896\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010001"
        )
    port map (
            in0 => \N__41192\,
            in1 => \N__43831\,
            in2 => \N__43777\,
            in3 => \N__40943\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__46754\,
            in1 => \N__43762\,
            in2 => \N__46645\,
            in3 => \N__45085\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_RNI33GU_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__42220\,
            in1 => \_gnd_net_\,
            in2 => \N__41276\,
            in3 => \N__46753\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__43832\,
            in1 => \N__43761\,
            in2 => \N__40928\,
            in3 => \N__40925\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIRDT63_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44897\,
            in1 => \N__45211\,
            in2 => \_gnd_net_\,
            in3 => \N__41323\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__41447\,
            in1 => \N__41324\,
            in2 => \N__41417\,
            in3 => \N__44846\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQ1_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__45023\,
            in1 => \N__41081\,
            in2 => \N__41274\,
            in3 => \N__41368\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIGLOQZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02_2_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41291\,
            in3 => \N__44844\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNIFQN02Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_RNICJ561_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41083\,
            in1 => \N__43954\,
            in2 => \N__41275\,
            in3 => \N__42221\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_153_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49764\,
            in2 => \_gnd_net_\,
            in3 => \N__44845\,
            lcout => \ppm_encoder_1.N_1818_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001011"
        )
    port map (
            in0 => \N__41225\,
            in1 => \N__43834\,
            in2 => \N__41202\,
            in3 => \N__43749\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__43833\,
            in1 => \N__41168\,
            in2 => \N__43772\,
            in3 => \N__41150\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_rep1_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__44847\,
            in1 => \N__49010\,
            in2 => \N__41107\,
            in3 => \N__41082\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIM4PT2_13_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__41692\,
            in1 => \N__45924\,
            in2 => \N__41486\,
            in3 => \N__45830\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIMC2D6_13_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__41663\,
            in1 => \_gnd_net_\,
            in2 => \N__41648\,
            in3 => \N__41630\,
            lcout => \ppm_encoder_1.elevator_RNIMC2D6Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI68LH2_13_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__41529\,
            in1 => \N__41580\,
            in2 => \N__45362\,
            in3 => \N__45478\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41484\,
            in1 => \N__46805\,
            in2 => \_gnd_net_\,
            in3 => \N__41530\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46583\,
            in1 => \_gnd_net_\,
            in2 => \N__41624\,
            in3 => \N__41581\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_13_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__41582\,
            in1 => \N__46376\,
            in2 => \N__41620\,
            in3 => \N__41594\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51440\,
            ce => 'H',
            sr => \N__49585\
        );

    \ppm_encoder_1.elevator_13_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__41531\,
            in1 => \N__41570\,
            in2 => \N__46394\,
            in3 => \N__41546\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51440\,
            ce => 'H',
            sr => \N__49585\
        );

    \ppm_encoder_1.throttle_13_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__41485\,
            in1 => \N__41519\,
            in2 => \N__46395\,
            in3 => \N__41495\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51440\,
            ce => 'H',
            sr => \N__49585\
        );

    \ppm_encoder_1.throttle_esr_RNIATV93_14_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__41815\,
            in1 => \N__41468\,
            in2 => \N__45831\,
            in3 => \N__45925\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIVU947_14_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41858\,
            in2 => \N__41840\,
            in3 => \N__41822\,
            lcout => \ppm_encoder_1.aileron_esr_RNIVU947Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIQ0MS2_14_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__41779\,
            in2 => \N__45499\,
            in3 => \N__45352\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46814\,
            in1 => \N__41816\,
            in2 => \_gnd_net_\,
            in3 => \N__41798\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46643\,
            in1 => \_gnd_net_\,
            in2 => \N__41783\,
            in3 => \N__41780\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44473\,
            in2 => \N__41765\,
            in3 => \N__41762\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51426\,
            ce => \N__44408\,
            sr => \N__49594\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47501\,
            in1 => \N__44188\,
            in2 => \N__47474\,
            in3 => \N__41753\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__41745\,
            in1 => \N__41722\,
            in2 => \N__44725\,
            in3 => \N__42174\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIGCMK2_0_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__43979\,
            in1 => \N__45993\,
            in2 => \N__41702\,
            in3 => \N__45304\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_0\,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111010000"
        )
    port map (
            in0 => \N__45448\,
            in1 => \N__44012\,
            in2 => \N__42062\,
            in3 => \N__42058\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__44722\,
            in1 => \N__46644\,
            in2 => \N__49799\,
            in3 => \N__43953\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110010"
        )
    port map (
            in0 => \N__44723\,
            in1 => \N__45161\,
            in2 => \N__49798\,
            in3 => \N__42217\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIMIMK2_3_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__42020\,
            in1 => \N__42278\,
            in2 => \N__45338\,
            in3 => \N__45786\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIT3R05_3_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \N__41995\,
            in1 => \N__41975\,
            in2 => \N__41942\,
            in3 => \N__45447\,
            lcout => \ppm_encoder_1.elevator_RNIT3R05Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.pid_prereg_esr_0_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48296\,
            lcout => \pid_side.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51399\,
            ce => \N__41890\,
            sr => \N__49604\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI78NT_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__42173\,
            in1 => \N__43946\,
            in2 => \N__42218\,
            in3 => \N__42420\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__47173\,
            in1 => \_gnd_net_\,
            in2 => \N__41861\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42419\,
            in2 => \_gnd_net_\,
            in3 => \N__42086\,
            lcout => \ppm_encoder_1.PPM_STATE_53_d\,
            ltout => \ppm_encoder_1.PPM_STATE_53_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__43944\,
            in1 => \N__42204\,
            in2 => \N__42236\,
            in3 => \N__42171\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47174\,
            in2 => \_gnd_net_\,
            in3 => \N__42421\,
            lcout => \ppm_encoder_1.N_134_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43945\,
            in1 => \N__42205\,
            in2 => \N__44724\,
            in3 => \N__42172\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42829\,
            in1 => \N__42068\,
            in2 => \N__42854\,
            in3 => \N__47086\,
            lcout => \ppm_encoder_1.N_232\,
            ltout => \ppm_encoder_1.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__49038\,
            in1 => \N__47163\,
            in2 => \N__42146\,
            in3 => \N__42423\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42830\,
            in1 => \N__47087\,
            in2 => \N__42395\,
            in3 => \N__42853\,
            lcout => \ppm_encoder_1.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__42424\,
            in1 => \N__42112\,
            in2 => \N__47172\,
            in3 => \N__42097\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51384\,
            ce => 'H',
            sr => \N__49609\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__42113\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42425\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51384\,
            ce => 'H',
            sr => \N__49609\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__47364\,
            in1 => \N__46977\,
            in2 => \N__46958\,
            in3 => \N__42087\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__46978\,
            in1 => \N__47365\,
            in2 => \N__46954\,
            in3 => \N__42422\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42359\,
            in1 => \N__47363\,
            in2 => \N__42341\,
            in3 => \N__46946\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42386\,
            in1 => \N__44490\,
            in2 => \_gnd_net_\,
            in3 => \N__42371\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51372\,
            ce => \N__44411\,
            sr => \N__49612\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44488\,
            in1 => \N__42242\,
            in2 => \_gnd_net_\,
            in3 => \N__42353\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51372\,
            ce => \N__44411\,
            sr => \N__49612\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43919\,
            in1 => \N__44489\,
            in2 => \_gnd_net_\,
            in3 => \N__42332\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51372\,
            ce => \N__44411\,
            sr => \N__49612\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42320\,
            in1 => \N__46976\,
            in2 => \N__42287\,
            in3 => \N__46995\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42314\,
            in1 => \N__42302\,
            in2 => \_gnd_net_\,
            in3 => \N__44491\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51372\,
            ce => \N__44411\,
            sr => \N__49612\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__42276\,
            in1 => \_gnd_net_\,
            in2 => \N__46655\,
            in3 => \N__42257\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47298\,
            in1 => \N__47320\,
            in2 => \N__47275\,
            in3 => \N__47341\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__42836\,
            in1 => \N__47547\,
            in2 => \N__42857\,
            in3 => \N__47244\,
            lcout => \ppm_encoder_1.N_139_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44826\,
            lcout => \ppm_encoder_1.N_1818_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47496\,
            in2 => \_gnd_net_\,
            in3 => \N__47523\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_RNI3C23_12_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43525\,
            lcout => \drone_H_disp_front_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47418\,
            in1 => \N__47442\,
            in2 => \N__47393\,
            in3 => \N__47466\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_8_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__47600\,
            in1 => \N__50495\,
            in2 => \N__42818\,
            in3 => \N__42630\,
            lcout => \pid_front.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51342\,
            ce => 'H',
            sr => \N__49622\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_0_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42610\,
            lcout => \drone_H_disp_front_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51335\,
            ce => \N__42527\,
            sr => \N__49625\
        );

    \pid_front.error_cry_0_c_inv_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42461\,
            in2 => \_gnd_net_\,
            in3 => \N__42472\,
            lcout => \pid_front.error_axb_0\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \pid_front.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_0_c_RNIC7KB_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42455\,
            in2 => \_gnd_net_\,
            in3 => \N__42428\,
            lcout => \pid_front.error_1\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_0\,
            carryout => \pid_front.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_1_c_RNIEALB_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43088\,
            in2 => \_gnd_net_\,
            in3 => \N__43064\,
            lcout => \pid_front.error_2\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_1\,
            carryout => \pid_front.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_2_c_RNIGDMB_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43061\,
            in2 => \_gnd_net_\,
            in3 => \N__43031\,
            lcout => \pid_front.error_3\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_2\,
            carryout => \pid_front.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_3_c_RNIABAG_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43028\,
            in2 => \N__43022\,
            in3 => \N__42998\,
            lcout => \pid_front.error_4\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_3\,
            carryout => \pid_front.error_cry_0_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_0_0_c_RNIOQKB_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42995\,
            in2 => \N__42989\,
            in3 => \N__42965\,
            lcout => \pid_front.error_5\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_0_0\,
            carryout => \pid_front.error_cry_1_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_1_0_c_RNIR0RF_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42962\,
            in2 => \N__42956\,
            in3 => \N__42932\,
            lcout => \pid_front.error_6\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_1_0\,
            carryout => \pid_front.error_cry_2_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_2_0_c_RNIU61K_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42929\,
            in2 => \N__42923\,
            in3 => \N__42899\,
            lcout => \pid_front.error_7\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_2_0\,
            carryout => \pid_front.error_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_3_0_c_RNI1D7O_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42896\,
            in2 => \N__42890\,
            in3 => \N__42860\,
            lcout => \pid_front.error_8\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \pid_front.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_4_c_RNILNBG_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43625\,
            in2 => \N__43619\,
            in3 => \N__43598\,
            lcout => \pid_front.error_9\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_4\,
            carryout => \pid_front.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_5_c_RNIVNFF_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43595\,
            in2 => \N__43586\,
            in3 => \N__43562\,
            lcout => \pid_front.error_10\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_5\,
            carryout => \pid_front.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_6_c_RNI3VJG_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43559\,
            in2 => \_gnd_net_\,
            in3 => \N__43538\,
            lcout => \pid_front.error_11\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_6\,
            carryout => \pid_front.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_7_c_RNIAPPM_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43535\,
            in2 => \N__43529\,
            in3 => \N__43484\,
            lcout => \pid_front.error_12\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_7\,
            carryout => \pid_front.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_8_c_RNIAC2E_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43481\,
            in2 => \N__43472\,
            in3 => \N__43436\,
            lcout => \pid_front.error_13\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_8\,
            carryout => \pid_front.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_9_c_RNIDG3E_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43433\,
            in2 => \N__48371\,
            in3 => \N__43409\,
            lcout => \pid_front.error_14\,
            ltout => OPEN,
            carryin => \pid_front.error_cry_9\,
            carryout => \pid_front.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_cry_10_c_RNINTDI_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__43406\,
            in1 => \N__48370\,
            in2 => \_gnd_net_\,
            in3 => \N__43394\,
            lcout => \pid_front.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_9_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43372\,
            in1 => \N__43256\,
            in2 => \N__43218\,
            in3 => \N__43100\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51493\,
            ce => 'H',
            sr => \N__49567\
        );

    \ppm_encoder_1.init_pulses_RNIFEN01_9_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__44163\,
            in1 => \N__45061\,
            in2 => \_gnd_net_\,
            in3 => \N__44922\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBAN01_5_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__43902\,
            in1 => \N__45060\,
            in2 => \_gnd_net_\,
            in3 => \N__44921\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIEDN01_8_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__44100\,
            in1 => \N__45062\,
            in2 => \_gnd_net_\,
            in3 => \N__44923\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIS1KT_15_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__44924\,
            in1 => \_gnd_net_\,
            in2 => \N__45123\,
            in3 => \N__44215\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_0_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__43978\,
            in1 => \N__46190\,
            in2 => \_gnd_net_\,
            in3 => \N__44042\,
            lcout => \ppm_encoder_1.throttleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51484\,
            ce => 'H',
            sr => \N__49578\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_0_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44010\,
            in1 => \N__43977\,
            in2 => \_gnd_net_\,
            in3 => \N__43958\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46538\,
            in2 => \N__43922\,
            in3 => \N__46001\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__43904\,
            in1 => \N__43840\,
            in2 => \N__43778\,
            in3 => \N__43646\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44501\,
            in1 => \N__46466\,
            in2 => \_gnd_net_\,
            in3 => \N__44357\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51471\,
            ce => \N__44404\,
            sr => \N__49586\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44348\,
            in1 => \N__44342\,
            in2 => \_gnd_net_\,
            in3 => \N__44503\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51471\,
            ce => \N__44404\,
            sr => \N__49586\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44499\,
            in1 => \N__44327\,
            in2 => \_gnd_net_\,
            in3 => \N__44315\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51471\,
            ce => \N__44404\,
            sr => \N__49586\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44500\,
            in1 => \N__44309\,
            in2 => \_gnd_net_\,
            in3 => \N__44300\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51471\,
            ce => \N__44404\,
            sr => \N__49586\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44288\,
            in1 => \N__44502\,
            in2 => \_gnd_net_\,
            in3 => \N__44276\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51471\,
            ce => \N__44404\,
            sr => \N__49586\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44260\,
            in1 => \N__47420\,
            in2 => \N__44230\,
            in3 => \N__47444\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_16_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__45182\,
            in1 => \N__44261\,
            in2 => \N__45221\,
            in3 => \N__44831\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51458\,
            ce => 'H',
            sr => \N__49595\
        );

    \ppm_encoder_1.pulses2count_17_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__44828\,
            in1 => \N__45218\,
            in2 => \N__44231\,
            in3 => \N__44252\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51458\,
            ce => 'H',
            sr => \N__49595\
        );

    \ppm_encoder_1.pulses2count_15_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__44216\,
            in1 => \N__44189\,
            in2 => \N__45220\,
            in3 => \N__44830\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51458\,
            ce => 'H',
            sr => \N__49595\
        );

    \ppm_encoder_1.pulses2count_18_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__44829\,
            in1 => \N__45254\,
            in2 => \N__45194\,
            in3 => \N__45219\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51458\,
            ce => 'H',
            sr => \N__49595\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45190\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIT2KT_0_16_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__45181\,
            in1 => \N__45132\,
            in2 => \_gnd_net_\,
            in3 => \N__44827\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44564\,
            in1 => \N__47276\,
            in2 => \N__44543\,
            in3 => \N__47300\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44492\,
            in1 => \N__44588\,
            in2 => \_gnd_net_\,
            in3 => \N__44579\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51441\,
            ce => \N__44409\,
            sr => \N__49599\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45683\,
            in1 => \N__44494\,
            in2 => \_gnd_net_\,
            in3 => \N__44558\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51441\,
            ce => \N__44409\,
            sr => \N__49599\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44493\,
            in1 => \N__44534\,
            in2 => \_gnd_net_\,
            in3 => \N__44522\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51441\,
            ce => \N__44409\,
            sr => \N__49599\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44516\,
            in1 => \_gnd_net_\,
            in2 => \N__44504\,
            in3 => \N__44420\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51441\,
            ce => \N__44409\,
            sr => \N__49599\
        );

    \ppm_encoder_1.throttle_RNISVPV2_7_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__45510\,
            in1 => \N__45965\,
            in2 => \N__45934\,
            in3 => \N__45803\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNILVOO6_7_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__45731\,
            in1 => \_gnd_net_\,
            in2 => \N__45710\,
            in3 => \N__45692\,
            lcout => \ppm_encoder_1.throttle_RNILVOO6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNICJ7O2_7_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__45570\,
            in1 => \N__45627\,
            in2 => \N__45339\,
            in3 => \N__45424\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46812\,
            in1 => \N__45511\,
            in2 => \_gnd_net_\,
            in3 => \N__45571\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46584\,
            in1 => \_gnd_net_\,
            in2 => \N__45686\,
            in3 => \N__45628\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__45629\,
            in1 => \N__45677\,
            in2 => \N__45662\,
            in3 => \N__46155\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51427\,
            ce => 'H',
            sr => \N__49605\
        );

    \ppm_encoder_1.elevator_7_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__45572\,
            in1 => \N__45617\,
            in2 => \N__46193\,
            in3 => \N__45605\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51427\,
            ce => 'H',
            sr => \N__49605\
        );

    \ppm_encoder_1.throttle_7_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__45560\,
            in1 => \N__45512\,
            in2 => \N__45545\,
            in3 => \N__46156\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51427\,
            ce => 'H',
            sr => \N__49605\
        );

    \ppm_encoder_1.elevator_RNI6D7O2_4_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__46677\,
            in1 => \N__46476\,
            in2 => \N__45452\,
            in3 => \N__45308\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_4_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__46478\,
            in1 => \N__46880\,
            in2 => \N__46191\,
            in3 => \N__46867\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51413\,
            ce => 'H',
            sr => \N__49610\
        );

    \ppm_encoder_1.elevator_4_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__46679\,
            in1 => \N__46151\,
            in2 => \N__46850\,
            in3 => \N__46835\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51413\,
            ce => 'H',
            sr => \N__49610\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46811\,
            in1 => \N__46413\,
            in2 => \_gnd_net_\,
            in3 => \N__46678\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46585\,
            in2 => \N__46481\,
            in3 => \N__46477\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_4_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__46457\,
            in1 => \N__46442\,
            in2 => \N__46192\,
            in3 => \N__46414\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51413\,
            ce => 'H',
            sr => \N__49610\
        );

    \ppm_encoder_1.aileron_0_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__46144\,
            in1 => \N__46031\,
            in2 => \_gnd_net_\,
            in3 => \N__45997\,
            lcout => \ppm_encoder_1.aileronZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51413\,
            ce => 'H',
            sr => \N__49610\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45977\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45971\,
            in2 => \N__48176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47126\,
            in2 => \N__48104\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46928\,
            in2 => \N__48173\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47054\,
            in2 => \N__48105\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47093\,
            in2 => \N__48174\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47021\,
            in2 => \N__48106\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46919\,
            in2 => \N__48175\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46910\,
            in2 => \N__48210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46898\,
            in2 => \N__48161\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47177\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47319\,
            in1 => \N__47150\,
            in2 => \N__47141\,
            in3 => \N__47340\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47120\,
            in1 => \N__47575\,
            in2 => \N__47108\,
            in3 => \N__47197\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__47222\,
            in1 => \N__46996\,
            in2 => \N__47201\,
            in3 => \N__47576\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47078\,
            in1 => \N__47221\,
            in2 => \N__47069\,
            in3 => \N__47246\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47525\,
            in1 => \N__47048\,
            in2 => \N__47036\,
            in3 => \N__47549\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_0_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46997\,
            in2 => \N__47014\,
            in3 => \N__47015\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_1_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46979\,
            in2 => \_gnd_net_\,
            in3 => \N__46961\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_2_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46953\,
            in2 => \_gnd_net_\,
            in3 => \N__47369\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_3_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47366\,
            in2 => \_gnd_net_\,
            in3 => \N__47345\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_4_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47342\,
            in2 => \_gnd_net_\,
            in3 => \N__47324\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_5_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47321\,
            in2 => \_gnd_net_\,
            in3 => \N__47303\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_6_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47299\,
            in2 => \_gnd_net_\,
            in3 => \N__47279\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_7_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47271\,
            in2 => \_gnd_net_\,
            in3 => \N__47249\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__51373\,
            ce => 'H',
            sr => \N__47714\
        );

    \ppm_encoder_1.counter_8_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47245\,
            in2 => \_gnd_net_\,
            in3 => \N__47225\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_9_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47220\,
            in2 => \_gnd_net_\,
            in3 => \N__47204\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_10_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47196\,
            in2 => \_gnd_net_\,
            in3 => \N__47180\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_11_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47574\,
            in2 => \_gnd_net_\,
            in3 => \N__47552\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_12_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47548\,
            in2 => \_gnd_net_\,
            in3 => \N__47528\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_13_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47524\,
            in2 => \_gnd_net_\,
            in3 => \N__47504\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_14_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47497\,
            in2 => \_gnd_net_\,
            in3 => \N__47477\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_15_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47467\,
            in2 => \_gnd_net_\,
            in3 => \N__47447\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__51360\,
            ce => 'H',
            sr => \N__47713\
        );

    \ppm_encoder_1.counter_16_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47443\,
            in2 => \_gnd_net_\,
            in3 => \N__47423\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__51350\,
            ce => 'H',
            sr => \N__47712\
        );

    \ppm_encoder_1.counter_17_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47419\,
            in2 => \_gnd_net_\,
            in3 => \N__47399\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__51350\,
            ce => 'H',
            sr => \N__47712\
        );

    \ppm_encoder_1.counter_18_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47391\,
            in2 => \_gnd_net_\,
            in3 => \N__47396\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51350\,
            ce => 'H',
            sr => \N__47712\
        );

    \pid_front.un1_pid_prereg_un1_pid_prereg_cry_1_c_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48784\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_22_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_1_THRU_LUT4_0_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48710\,
            in2 => \_gnd_net_\,
            in3 => \N__47684\,
            lcout => \pid_front.un1_pid_prereg_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_1\,
            carryout => \pid_front.un1_pid_prereg_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_2_THRU_LUT4_0_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50377\,
            in2 => \_gnd_net_\,
            in3 => \N__47666\,
            lcout => \pid_front.un1_pid_prereg_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_2\,
            carryout => \pid_front.un1_pid_prereg_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_3_THRU_LUT4_0_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48625\,
            in2 => \_gnd_net_\,
            in3 => \N__47648\,
            lcout => \pid_front.un1_pid_prereg_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_3\,
            carryout => \pid_front.un1_pid_prereg_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_4_THRU_LUT4_0_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48667\,
            in2 => \N__48207\,
            in3 => \N__47630\,
            lcout => \pid_front.un1_pid_prereg_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_4\,
            carryout => \pid_front.un1_pid_prereg_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_5_THRU_LUT4_0_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48165\,
            in2 => \N__50311\,
            in3 => \N__47615\,
            lcout => \pid_front.un1_pid_prereg_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_5\,
            carryout => \pid_front.un1_pid_prereg_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_6_THRU_LUT4_0_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48169\,
            in2 => \N__50416\,
            in3 => \N__47603\,
            lcout => \pid_front.un1_pid_prereg_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_6\,
            carryout => \pid_front.un1_pid_prereg_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_7_THRU_LUT4_0_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50491\,
            in2 => \N__48209\,
            in3 => \N__47594\,
            lcout => \pid_front.un1_pid_prereg_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_7\,
            carryout => \pid_front.un1_pid_prereg_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_8_THRU_LUT4_0_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48739\,
            in2 => \N__48208\,
            in3 => \N__47579\,
            lcout => \pid_front.un1_pid_prereg_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_9_THRU_LUT4_0_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50452\,
            in2 => \N__48232\,
            in3 => \N__48254\,
            lcout => \pid_front.un1_pid_prereg_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_9\,
            carryout => \pid_front.un1_pid_prereg_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_10_THRU_LUT4_0_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51796\,
            in2 => \_gnd_net_\,
            in3 => \N__48239\,
            lcout => \pid_front.un1_pid_prereg_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_10\,
            carryout => \pid_front.un1_pid_prereg_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_11_THRU_LUT4_0_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51760\,
            in2 => \N__48231\,
            in3 => \N__47786\,
            lcout => \pid_front.un1_pid_prereg_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_11\,
            carryout => \pid_front.un1_pid_prereg_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_12_THRU_LUT4_0_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51856\,
            in2 => \_gnd_net_\,
            in3 => \N__47771\,
            lcout => \pid_front.un1_pid_prereg_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_12\,
            carryout => \pid_front.un1_pid_prereg_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_13_THRU_LUT4_0_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50539\,
            in2 => \_gnd_net_\,
            in3 => \N__47756\,
            lcout => \pid_front.un1_pid_prereg_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_13\,
            carryout => \pid_front.un1_pid_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_14_THRU_LUT4_0_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51823\,
            in2 => \_gnd_net_\,
            in3 => \N__47744\,
            lcout => \pid_front.un1_pid_prereg_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_14\,
            carryout => \pid_front.un1_pid_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_15_THRU_LUT4_0_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50341\,
            in2 => \_gnd_net_\,
            in3 => \N__47732\,
            lcout => \pid_front.un1_pid_prereg_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_15\,
            carryout => \pid_front.un1_pid_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_16_THRU_LUT4_0_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51562\,
            in2 => \_gnd_net_\,
            in3 => \N__47717\,
            lcout => \pid_front.un1_pid_prereg_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \pid_front.un1_pid_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_17_THRU_LUT4_0_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50251\,
            in2 => \_gnd_net_\,
            in3 => \N__48578\,
            lcout => \pid_front.un1_pid_prereg_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_17\,
            carryout => \pid_front.un1_pid_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_18_THRU_LUT4_0_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51907\,
            in2 => \_gnd_net_\,
            in3 => \N__48563\,
            lcout => \pid_front.un1_pid_prereg_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_18\,
            carryout => \pid_front.un1_pid_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.un1_pid_prereg_cry_19_THRU_LUT4_0_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51711\,
            in2 => \_gnd_net_\,
            in3 => \N__48548\,
            lcout => \pid_front.un1_pid_prereg_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_front.un1_pid_prereg_cry_19\,
            carryout => \pid_front.un1_pid_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.pid_prereg_esr_21_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51712\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48545\,
            lcout => \pid_front.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51328\,
            ce => \N__48482\,
            sr => \N__49627\
        );

    \dron_frame_decoder_1.source_H_disp_front_esr_14_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48455\,
            lcout => \drone_H_disp_front_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51321\,
            ce => \N__48359\,
            sr => \N__49628\
        );

    \GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49746\,
            lcout => \GB_BUFFER_reset_system_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_side.error_p_reg_0_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48289\,
            in1 => \N__48308\,
            in2 => \_gnd_net_\,
            in3 => \N__50178\,
            lcout => \pid_side.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51460\,
            ce => 'H',
            sr => \N__50697\
        );

    \pid_side.error_p_reg_1_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50177\,
            in1 => \N__49854\,
            in2 => \_gnd_net_\,
            in3 => \N__48278\,
            lcout => \pid_side.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51460\,
            ce => 'H',
            sr => \N__50697\
        );

    \pid_side.error_p_reg_3_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50179\,
            in1 => \N__50095\,
            in2 => \_gnd_net_\,
            in3 => \N__50126\,
            lcout => \pid_side.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51460\,
            ce => 'H',
            sr => \N__50697\
        );

    \pid_front.error_p_reg_0_LC_20_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51658\,
            in1 => \N__50059\,
            in2 => \_gnd_net_\,
            in3 => \N__50081\,
            lcout => \pid_front.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51351\,
            ce => 'H',
            sr => \N__50690\
        );

    \pid_side.pid_prereg_1_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__50048\,
            in1 => \N__49867\,
            in2 => \_gnd_net_\,
            in3 => \N__49821\,
            lcout => \pid_side.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51415\,
            ce => 'H',
            sr => \N__49626\
        );

    \pid_front.state_RNIVIRQ_1_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49064\,
            in2 => \_gnd_net_\,
            in3 => \N__49046\,
            lcout => \pid_front.state_RNIVIRQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_front.error_p_reg_1_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51657\,
            in1 => \N__48774\,
            in2 => \_gnd_net_\,
            in3 => \N__48794\,
            lcout => \pid_front.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51361\,
            ce => 'H',
            sr => \N__50691\
        );

    \pid_front.error_p_reg_9_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51660\,
            in1 => \N__48738\,
            in2 => \_gnd_net_\,
            in3 => \N__48755\,
            lcout => \pid_front.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51375\,
            ce => 'H',
            sr => \N__50692\
        );

    \pid_front.error_p_reg_2_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51659\,
            in1 => \N__48702\,
            in2 => \_gnd_net_\,
            in3 => \N__48719\,
            lcout => \pid_front.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51375\,
            ce => 'H',
            sr => \N__50692\
        );

    \pid_front.error_p_reg_5_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__48660\,
            in1 => \_gnd_net_\,
            in2 => \N__51680\,
            in3 => \N__48683\,
            lcout => \pid_front.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51386\,
            ce => 'H',
            sr => \N__50693\
        );

    \pid_front.error_p_reg_4_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48612\,
            in1 => \N__51671\,
            in2 => \_gnd_net_\,
            in3 => \N__48638\,
            lcout => \pid_front.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51386\,
            ce => 'H',
            sr => \N__50693\
        );

    \pid_front.error_p_reg_14_LC_24_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50552\,
            in1 => \N__51665\,
            in2 => \_gnd_net_\,
            in3 => \N__50523\,
            lcout => \pid_front.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51416\,
            ce => 'H',
            sr => \N__50696\
        );

    \pid_front.error_p_reg_8_LC_24_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51663\,
            in1 => \N__50484\,
            in2 => \_gnd_net_\,
            in3 => \N__50504\,
            lcout => \pid_front.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51416\,
            ce => 'H',
            sr => \N__50696\
        );

    \pid_front.error_p_reg_10_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50468\,
            in1 => \N__51664\,
            in2 => \_gnd_net_\,
            in3 => \N__50445\,
            lcout => \pid_front.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51416\,
            ce => 'H',
            sr => \N__50696\
        );

    \pid_front.error_p_reg_7_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51662\,
            in1 => \N__50409\,
            in2 => \_gnd_net_\,
            in3 => \N__50426\,
            lcout => \pid_front.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51416\,
            ce => 'H',
            sr => \N__50696\
        );

    \pid_front.error_p_reg_3_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51661\,
            in1 => \N__50373\,
            in2 => \_gnd_net_\,
            in3 => \N__50390\,
            lcout => \pid_front.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51416\,
            ce => 'H',
            sr => \N__50696\
        );

    \pid_front.error_p_reg_16_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51668\,
            in1 => \N__50334\,
            in2 => \_gnd_net_\,
            in3 => \N__50354\,
            lcout => \pid_front.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_6_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__50292\,
            in1 => \N__51670\,
            in2 => \_gnd_net_\,
            in3 => \N__50318\,
            lcout => \pid_front.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_18_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50273\,
            in1 => \N__51676\,
            in2 => \_gnd_net_\,
            in3 => \N__50244\,
            lcout => \pid_front.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_19_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__51891\,
            in1 => \N__51669\,
            in2 => \_gnd_net_\,
            in3 => \N__51920\,
            lcout => \pid_front.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_13_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51667\,
            in1 => \N__51855\,
            in2 => \_gnd_net_\,
            in3 => \N__51872\,
            lcout => \pid_front.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_15_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51675\,
            in1 => \N__51822\,
            in2 => \_gnd_net_\,
            in3 => \N__51836\,
            lcout => \pid_front.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_11_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51666\,
            in1 => \N__51795\,
            in2 => \_gnd_net_\,
            in3 => \N__51803\,
            lcout => \pid_front.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_12_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51677\,
            in1 => \N__51776\,
            in2 => \_gnd_net_\,
            in3 => \N__51750\,
            lcout => \pid_front.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51401\,
            ce => 'H',
            sr => \N__50695\
        );

    \pid_front.error_p_reg_20_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51699\,
            in1 => \N__51731\,
            in2 => \_gnd_net_\,
            in3 => \N__51679\,
            lcout => \pid_front.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51387\,
            ce => 'H',
            sr => \N__50694\
        );

    \pid_front.error_p_reg_17_LC_24_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__51561\,
            in1 => \N__51678\,
            in2 => \_gnd_net_\,
            in3 => \N__51575\,
            lcout => \pid_front.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51387\,
            ce => 'H',
            sr => \N__50694\
        );
end \INTERFACE\;
