-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Apr 14 2019 14:18:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "Pc2drone" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of Pc2drone
entity Pc2drone is
port (
    uart_input_pc : in std_logic;
    debug_CH5_31B : out std_logic;
    debug_CH3_20A : out std_logic;
    debug_CH0_16A : out std_logic;
    uart_input_drone : in std_logic;
    ppm_output : out std_logic;
    debug_CH6_5B : out std_logic;
    debug_CH2_18A : out std_logic;
    debug_CH4_2A : out std_logic;
    debug_CH1_0A : out std_logic;
    clk_system : in std_logic);
end Pc2drone;

-- Architecture of Pc2drone
-- View name is \INTERFACE\
architecture \INTERFACE\ of Pc2drone is

signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \pid_alt.O_0_6\ : std_logic;
signal \pid_alt.O_0_14\ : std_logic;
signal \pid_alt.O_0_12\ : std_logic;
signal \pid_alt.O_0_21\ : std_logic;
signal \pid_alt.O_0_7\ : std_logic;
signal \pid_alt.O_0_17\ : std_logic;
signal \pid_alt.O_0_15\ : std_logic;
signal \pid_alt.O_0_16\ : std_logic;
signal \pid_alt.O_0_5\ : std_logic;
signal \pid_alt.O_0_22\ : std_logic;
signal \pid_alt.O_0_4\ : std_logic;
signal \pid_alt.O_0_10\ : std_logic;
signal \pid_alt.O_0_23\ : std_logic;
signal \pid_alt.O_0_11\ : std_logic;
signal \pid_alt.O_0_13\ : std_logic;
signal \pid_alt.O_0_24\ : std_logic;
signal \pid_alt.O_0_19\ : std_logic;
signal \pid_alt.O_0_20\ : std_logic;
signal \pid_alt.O_0_18\ : std_logic;
signal \pid_alt.O_0_9\ : std_logic;
signal \pid_alt.error_p_regZ0Z_15\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_13\ : std_logic;
signal \pid_alt.O_18\ : std_logic;
signal \pid_alt.error_p_regZ0Z_14\ : std_logic;
signal \pid_alt.O_23\ : std_logic;
signal \pid_alt.O_4\ : std_logic;
signal \pid_alt.O_17\ : std_logic;
signal \pid_alt.O_19\ : std_logic;
signal \pid_alt.O_20\ : std_logic;
signal \pid_alt.O_21\ : std_logic;
signal \pid_alt.O_22\ : std_logic;
signal \pid_alt.O_6\ : std_logic;
signal \pid_alt.O_24\ : std_logic;
signal \pid_alt.O_15\ : std_logic;
signal \pid_alt.error_p_regZ0Z_11\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_\ : std_logic;
signal \pid_alt.O_16\ : std_logic;
signal \pid_alt.error_p_regZ0Z_12\ : std_logic;
signal \pid_alt.O_14\ : std_logic;
signal \pid_alt.error_p_regZ0Z_10\ : std_logic;
signal \pid_alt.O_5\ : std_logic;
signal \pid_alt.O_7\ : std_logic;
signal \pid_alt.O_9\ : std_logic;
signal \pid_alt.O_8\ : std_logic;
signal \pid_alt.N_62_mux_cascade_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5\ : std_logic;
signal \pid_alt.N_37_cascade_\ : std_logic;
signal \pid_alt.N_62_mux\ : std_logic;
signal \pid_alt.N_37\ : std_logic;
signal \pid_alt.error_p_regZ0Z_1\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_2\ : std_logic;
signal \pid_alt.error_p_regZ0Z_17\ : std_logic;
signal \pid_alt.error_p_regZ0Z_5\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_\ : std_logic;
signal \pid_alt.error_p_regZ0Z_19\ : std_logic;
signal alt_ki_0 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_4\ : std_logic;
signal throttle_command_6 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7\ : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_13\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_5\ : std_logic;
signal \ppm_encoder_1.N_297_cascade_\ : std_logic;
signal scaler_2_data_5 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_10\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_14\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_9\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\ : std_logic;
signal throttle_command_9 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_9\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_9\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\ : std_logic;
signal \pid_alt.O_0_8\ : std_logic;
signal \pid_alt.error_p_regZ0Z_4\ : std_logic;
signal alt_kp_2 : std_logic;
signal alt_ki_4 : std_logic;
signal alt_ki_1 : std_logic;
signal alt_ki_2 : std_logic;
signal alt_ki_3 : std_logic;
signal alt_ki_5 : std_logic;
signal alt_ki_6 : std_logic;
signal \pid_alt.O_12\ : std_logic;
signal \pid_alt.error_p_regZ0Z_8\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_\ : std_logic;
signal \pid_alt.O_13\ : std_logic;
signal \pid_alt.error_p_regZ0Z_9\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pid_alt.error_1\ : std_logic;
signal \pid_alt.error_cry_0\ : std_logic;
signal \pid_alt.error_2\ : std_logic;
signal \pid_alt.error_cry_1\ : std_logic;
signal \pid_alt.error_3\ : std_logic;
signal \pid_alt.error_cry_2\ : std_logic;
signal \pid_alt.error_4\ : std_logic;
signal \pid_alt.error_cry_3\ : std_logic;
signal \pid_alt.error_5\ : std_logic;
signal \pid_alt.error_cry_4\ : std_logic;
signal \pid_alt.error_6\ : std_logic;
signal \pid_alt.error_cry_5\ : std_logic;
signal \pid_alt.error_7\ : std_logic;
signal \pid_alt.error_cry_6\ : std_logic;
signal \pid_alt.error_cry_7\ : std_logic;
signal \pid_alt.error_8\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pid_alt.error_9\ : std_logic;
signal \pid_alt.error_cry_8\ : std_logic;
signal \pid_alt.error_10\ : std_logic;
signal \pid_alt.error_cry_9\ : std_logic;
signal \pid_alt.error_11\ : std_logic;
signal \pid_alt.error_cry_10\ : std_logic;
signal \pid_alt.error_12\ : std_logic;
signal \pid_alt.error_cry_11\ : std_logic;
signal \pid_alt.error_13\ : std_logic;
signal \pid_alt.error_cry_12\ : std_logic;
signal \pid_alt.error_14\ : std_logic;
signal \pid_alt.error_cry_13\ : std_logic;
signal \pid_alt.error_cry_14\ : std_logic;
signal \pid_alt.error_15\ : std_logic;
signal \pid_alt.m35_e_2\ : std_logic;
signal \pid_alt.m35_e_2_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5\ : std_logic;
signal \pid_alt.m35_e_3\ : std_logic;
signal \pid_alt.m21_e_2_cascade_\ : std_logic;
signal \pid_alt.m21_e_0_cascade_\ : std_logic;
signal \pid_alt.m21_e_8\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_0\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8\ : std_logic;
signal \pid_alt.drone_altitude_i_0\ : std_logic;
signal drone_altitude_0 : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_\ : std_logic;
signal \pid_alt.N_9_0\ : std_logic;
signal \pid_alt.m21_e_9\ : std_logic;
signal \pid_alt.N_9_0_cascade_\ : std_logic;
signal \pid_alt.m21_e_10\ : std_logic;
signal \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_\ : std_logic;
signal \pid_alt.un1_reset_1_0_i\ : std_logic;
signal \pid_alt.un1_reset_1_0_i_cascade_\ : std_logic;
signal \pid_alt.N_60_i_0\ : std_logic;
signal \pid_alt.error_p_regZ0Z_0\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_0\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_1\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_2\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_3\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI91H61Z0Z_4\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_4\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_5\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_6\ : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_7\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_8\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_9\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_10\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_11\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_12\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_13\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_14\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14\ : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIKU581Z0Z_15\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_15\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIO2681Z0Z_16\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_16\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNID23KZ0Z_17\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIS6681Z0Z_17\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_17\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI0B681Z0Z_18\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_18\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIIU781Z0Z_19\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIH63KZ0Z_19\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_19\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI2G981Z0Z_20\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_20\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_21\ : std_logic;
signal \pid_alt.pid_preregZ0Z_14\ : std_logic;
signal \pid_alt.pid_preregZ0Z_19\ : std_logic;
signal \pid_alt.pid_preregZ0Z_20\ : std_logic;
signal \pid_alt.pid_preregZ0Z_21\ : std_logic;
signal \pid_alt.pid_preregZ0Z_16\ : std_logic;
signal \pid_alt.pid_preregZ0Z_15\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_\ : std_logic;
signal \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_17\ : std_logic;
signal \pid_alt.pid_preregZ0Z_18\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_2_3\ : std_logic;
signal \pid_alt.source_pid_9_0_0_4\ : std_logic;
signal throttle_command_5 : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_11\ : std_logic;
signal \ppm_encoder_1.N_303_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_11\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_11\ : std_logic;
signal throttle_command_11 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_7\ : std_logic;
signal \ppm_encoder_1.N_299_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_7\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\ : std_logic;
signal throttle_command_7 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_6\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_13\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_5\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_5\ : std_logic;
signal \ppm_encoder_1.throttle_RNIN3352Z0Z_0\ : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_5\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_4\ : std_logic;
signal \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_5\ : std_logic;
signal \ppm_encoder_1.throttle_RNIJII96Z0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_7\ : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal \ppm_encoder_1.throttle_RNITSI96Z0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_8\ : std_logic;
signal \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_9\ : std_logic;
signal \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_13\ : std_logic;
signal \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_12\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_13\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_15\ : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_18\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_16\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\ : std_logic;
signal \bfn_2_28_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_4\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_8\ : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_11\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_15\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_15\ : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_cry_17\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_18\ : std_logic;
signal alt_kp_3 : std_logic;
signal alt_kp_6 : std_logic;
signal alt_kp_5 : std_logic;
signal alt_kp_1 : std_logic;
signal alt_kp_0 : std_logic;
signal drone_altitude_15 : std_logic;
signal alt_command_2 : std_logic;
signal alt_command_3 : std_logic;
signal alt_command_1 : std_logic;
signal \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8\ : std_logic;
signal \Commands_frame_decoder.source_CH1data8_cascade_\ : std_logic;
signal alt_command_0 : std_logic;
signal drone_altitude_i_7 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_7\ : std_logic;
signal drone_altitude_i_8 : std_logic;
signal drone_altitude_i_9 : std_logic;
signal drone_altitude_i_10 : std_logic;
signal drone_altitude_i_11 : std_logic;
signal \pid_alt.error_axbZ0Z_1\ : std_logic;
signal drone_altitude_1 : std_logic;
signal \pid_alt.error_axbZ0Z_12\ : std_logic;
signal drone_altitude_12 : std_logic;
signal \pid_alt.error_axbZ0Z_13\ : std_logic;
signal drone_altitude_13 : std_logic;
signal \pid_alt.error_axbZ0Z_14\ : std_logic;
signal \pid_alt.error_axbZ0Z_2\ : std_logic;
signal \pid_alt.error_axbZ0Z_3\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_1\ : std_logic;
signal \pid_alt.error_i_regZ0Z_1\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_1\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_0\ : std_logic;
signal \pid_alt.error_i_regZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_2\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_2\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_1\ : std_logic;
signal \pid_alt.error_i_regZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_3\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_3\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_2\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_4\ : std_logic;
signal \pid_alt.error_i_regZ0Z_4\ : std_logic;
signal \pid_alt.error_i_acumm7lto4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_3\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_5\ : std_logic;
signal \pid_alt.error_i_regZ0Z_5\ : std_logic;
signal \pid_alt.error_i_acumm7lto5\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_4\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_5\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_7\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_6\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_7\ : std_logic;
signal \pid_alt.error_i_regZ0Z_8\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_8\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_8\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \pid_alt.error_i_regZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_9\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_9\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_8\ : std_logic;
signal \pid_alt.error_i_regZ0Z_10\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_10\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_10\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_9\ : std_logic;
signal \pid_alt.error_i_regZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_11\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_11\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_10\ : std_logic;
signal \pid_alt.error_i_regZ0Z_12\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_12\ : std_logic;
signal \pid_alt.error_i_acumm7lto12\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_11\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_13\ : std_logic;
signal \pid_alt.error_i_regZ0Z_13\ : std_logic;
signal \pid_alt.error_i_acumm7lto13\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_12\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_13\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_15\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_16\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_18\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_20\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_21\ : std_logic;
signal \pid_alt.state_0_g_0\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_0\ : std_logic;
signal \pid_alt.error_i_regZ0Z_0\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_0\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO\ : std_logic;
signal \pid_alt.error_i_regZ0Z_14\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_14\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_16\ : std_logic;
signal \pid_alt.error_i_regZ0Z_19\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_19\ : std_logic;
signal \pid_alt.error_p_regZ0Z_16\ : std_logic;
signal \pid_alt.error_i_regZ0Z_16\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIB03KZ0Z_16\ : std_logic;
signal \ppm_encoder_1.N_306\ : std_logic;
signal \dron_frame_decoder_1.N_194_4_cascade_\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_20\ : std_logic;
signal \pid_alt.m7_e_4\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO\ : std_logic;
signal \pid_alt.error_i_regZ0Z_15\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_15\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO\ : std_logic;
signal \pid_alt.error_i_regZ0Z_17\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_17\ : std_logic;
signal \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO\ : std_logic;
signal \pid_alt.error_i_acumm_preregZ0Z_18\ : std_logic;
signal \pid_alt.source_pid_9_0_tz_6\ : std_logic;
signal \pid_alt.source_pid_9_0_tz_6_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_8\ : std_logic;
signal \pid_alt.pid_preregZ0Z_11\ : std_logic;
signal \pid_alt.pid_preregZ0Z_9\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\ : std_logic;
signal \pid_alt.pid_preregZ0Z_6\ : std_logic;
signal \pid_alt.pid_preregZ0Z_0\ : std_logic;
signal \pid_alt.pid_preregZ0Z_10\ : std_logic;
signal \pid_alt.pid_preregZ0Z_7\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\ : std_logic;
signal \pid_alt.N_92_cascade_\ : std_logic;
signal \pid_alt.un1_reset_1_cascade_\ : std_logic;
signal \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\ : std_logic;
signal \pid_alt.un1_reset_0_i_cascade_\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_13\ : std_logic;
signal \bfn_3_22_0_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_14\ : std_logic;
signal \pid_alt.pid_preregZ0Z_3\ : std_logic;
signal \pid_alt.pid_preregZ0Z_13\ : std_logic;
signal \pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6\ : std_logic;
signal \pid_alt.N_88\ : std_logic;
signal \pid_alt.pid_preregZ0Z_4\ : std_logic;
signal \pid_alt.N_88_cascade_\ : std_logic;
signal \pid_alt.N_90\ : std_logic;
signal \pid_alt.pid_preregZ0Z_22\ : std_logic;
signal \pid_alt.pid_preregZ0Z_2\ : std_logic;
signal \pid_alt.N_90_cascade_\ : std_logic;
signal \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\ : std_logic;
signal \pid_alt.N_60_i_1\ : std_logic;
signal \pid_alt.un1_reset_0_i\ : std_logic;
signal \pid_alt.pid_preregZ0Z_5\ : std_logic;
signal \pid_alt.pid_preregZ0Z_12\ : std_logic;
signal \pid_alt.N_130\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_1\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIALN65Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_4_cascade_\ : std_logic;
signal \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNI5V123Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_3\ : std_logic;
signal \ppm_encoder_1.throttle_RNI82223Z0Z_3\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_10\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_9\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_10\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_7\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_8\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_2\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_6\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_16\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_4\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_4\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_4\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_1\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_11_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_10_5\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_14\ : std_logic;
signal \ppm_encoder_1.N_319_cascade_\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_12\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_2\ : std_logic;
signal alt_kp_7 : std_logic;
signal alt_kp_4 : std_logic;
signal \pid_alt.O_10\ : std_logic;
signal \pid_alt.error_p_regZ0Z_6\ : std_logic;
signal \pid_alt.error_i_regZ0Z_6\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_6\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7\ : std_logic;
signal \pid_alt.O_11\ : std_logic;
signal \pid_alt.N_422_0_g\ : std_logic;
signal \pid_alt.error_p_regZ0Z_7\ : std_logic;
signal \pid_alt.error_i_regZ0Z_7\ : std_logic;
signal \pid_alt.error_i_acummZ0Z_7\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_11\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_9\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_10\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_8\ : std_logic;
signal drone_altitude_14 : std_logic;
signal drone_altitude_2 : std_logic;
signal drone_altitude_3 : std_logic;
signal \pid_alt.error_i_regZ0Z_18\ : std_logic;
signal \pid_alt.error_p_regZ0Z_18\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNIF43KZ0Z_18\ : std_logic;
signal \pid_alt.error_i_regZ0Z_20\ : std_logic;
signal \pid_alt.error_p_regZ0Z_20\ : std_logic;
signal \pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20\ : std_logic;
signal \frame_decoder_CH2data_1\ : std_logic;
signal \frame_decoder_CH2data_2\ : std_logic;
signal \frame_decoder_CH2data_3\ : std_logic;
signal \frame_decoder_CH2data_4\ : std_logic;
signal \frame_decoder_CH2data_5\ : std_logic;
signal \frame_decoder_CH2data_6\ : std_logic;
signal \scaler_2.N_881_i_l_ofxZ0\ : std_logic;
signal \frame_decoder_CH2data_7\ : std_logic;
signal \scaler_2.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \scaler_2.un2_source_data_0\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\ : std_logic;
signal scaler_2_data_7 : std_logic;
signal \scaler_2.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\ : std_logic;
signal scaler_2_data_9 : std_logic;
signal \scaler_2.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\ : std_logic;
signal scaler_2_data_11 : std_logic;
signal \scaler_2.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\ : std_logic;
signal \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \scaler_2.un2_source_data_0_cry_9\ : std_logic;
signal scaler_2_data_14 : std_logic;
signal alt_ki_7 : std_logic;
signal \pid_alt.un1_pid_prereg_0_axb_1\ : std_logic;
signal \pid_alt.un1_pid_prereg_0_cry_0_THRU_CO\ : std_logic;
signal \pid_alt.pid_preregZ0Z_1\ : std_logic;
signal \N_423_g\ : std_logic;
signal \pid_alt.N_422_0\ : std_logic;
signal \pid_alt.state_1_0_0\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_11\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_7\ : std_logic;
signal throttle_command_10 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\ : std_logic;
signal throttle_command_13 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\ : std_logic;
signal throttle_command_2 : std_logic;
signal throttle_command_4 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\ : std_logic;
signal \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_12\ : std_logic;
signal \ppm_encoder_1.N_304_cascade_\ : std_logic;
signal scaler_2_data_12 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_12\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_12\ : std_logic;
signal throttle_command_12 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_12\ : std_logic;
signal \ppm_encoder_1.init_pulses_3_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_0_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_8\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\ : std_logic;
signal \ppm_encoder_1.throttle_RNIONI96Z0Z_8\ : std_logic;
signal \ppm_encoder_1.init_pulses_1_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.init_pulses_2_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.un2_throttle_iv_1_8\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_8\ : std_logic;
signal throttle_command_8 : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_8\ : std_logic;
signal scaler_2_data_8 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_4\ : std_logic;
signal \ppm_encoder_1.N_296\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_4\ : std_logic;
signal \ppm_encoder_1.N_227\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_0_11\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_10\ : std_logic;
signal \ppm_encoder_1.N_302_cascade_\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_145_17_cascade_\ : std_logic;
signal \ppm_encoder_1.N_145_17\ : std_logic;
signal \ppm_encoder_1.N_238_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_4\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_11\ : std_logic;
signal \ppm_encoder_1.N_300\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_8\ : std_logic;
signal \ppm_encoder_1.N_301\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_9\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_1\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_11\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_d_12\ : std_logic;
signal \ppm_encoder_1.un1_init_pulses_3_axb_16\ : std_logic;
signal \dron_frame_decoder_1.drone_altitude_4\ : std_logic;
signal drone_altitude_i_4 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_5\ : std_logic;
signal drone_altitude_i_5 : std_logic;
signal \dron_frame_decoder_1.drone_altitude_6\ : std_logic;
signal drone_altitude_i_6 : std_logic;
signal alt_command_4 : std_logic;
signal alt_command_5 : std_logic;
signal alt_command_6 : std_logic;
signal alt_command_7 : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\ : std_logic;
signal \frame_decoder_OFF2data_1\ : std_logic;
signal \frame_decoder_OFF2data_2\ : std_logic;
signal \frame_decoder_OFF2data_3\ : std_logic;
signal \frame_decoder_OFF2data_4\ : std_logic;
signal \frame_decoder_OFF2data_5\ : std_logic;
signal \frame_decoder_OFF2data_6\ : std_logic;
signal \frame_decoder_OFF2data_7\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\ : std_logic;
signal \dron_frame_decoder_1.state_RNO_1Z0Z_0\ : std_logic;
signal \dron_frame_decoder_1.N_194_4\ : std_logic;
signal \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\ : std_logic;
signal \dron_frame_decoder_1.state_RNO_0Z0Z_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_0\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_1\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3\ : std_logic;
signal \debug_CH1_0A_c\ : std_logic;
signal \pid_alt.N_60_i\ : std_logic;
signal \pid_alt.state_RNIFCSD1Z0Z_0\ : std_logic;
signal \frame_decoder_OFF2data_0\ : std_logic;
signal \frame_decoder_CH2data_0\ : std_logic;
signal scaler_2_data_4 : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\ : std_logic;
signal \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_13\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_13\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_8\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_8\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\ : std_logic;
signal scaler_2_data_10 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_10\ : std_logic;
signal scaler_2_data_13 : std_logic;
signal \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_10\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_elevator_cry_13\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_14\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\ : std_logic;
signal scaler_2_data_6 : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_6\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_6\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_13\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_13\ : std_logic;
signal throttle_command_0 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\ : std_logic;
signal throttle_command_1 : std_logic;
signal \ppm_encoder_1.throttleZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\ : std_logic;
signal throttle_command_3 : std_logic;
signal pid_altitude_dv : std_logic;
signal \ppm_encoder_1.throttleZ0Z_3\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_1\ : std_logic;
signal \ppm_encoder_1.N_140_0_cascade_\ : std_logic;
signal \ppm_encoder_1.N_145\ : std_logic;
signal ppm_output_c : std_logic;
signal \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_2\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_0\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_1\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\ : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_1\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_2\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_4\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_5\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_6\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_7\ : std_logic;
signal \bfn_5_28_0_\ : std_logic;
signal \ppm_encoder_1.counter24_0_data_tmp_8\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_10\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_10\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\ : std_logic;
signal \ppm_encoder_1.N_238\ : std_logic;
signal \ppm_encoder_1.counter24_0_N_2_THRU_CO\ : std_logic;
signal \ppm_encoder_1.PPM_STATEZ0Z_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_3\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\ : std_logic;
signal \bfn_5_29_0_\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_7\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_8\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_9\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_10\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_11\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_rudder_cry_13\ : std_logic;
signal \bfn_5_30_0_\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.state_RNIF38SZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.N_390_0\ : std_logic;
signal \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\ : std_logic;
signal \dron_frame_decoder_1.N_382_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_3_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0\ : std_logic;
signal \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\ : std_logic;
signal \GB_BUFFER_reset_system_g_THRU_CO\ : std_logic;
signal uart_drone_data_0 : std_logic;
signal uart_drone_data_1 : std_logic;
signal uart_drone_data_2 : std_logic;
signal uart_drone_data_3 : std_logic;
signal uart_drone_data_4 : std_logic;
signal uart_drone_data_5 : std_logic;
signal uart_drone_data_6 : std_logic;
signal uart_drone_data_7 : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \frame_decoder_CH4data_1\ : std_logic;
signal \frame_decoder_OFF4data_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_OFF4data_2\ : std_logic;
signal \frame_decoder_CH4data_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_CH4data_3\ : std_logic;
signal \frame_decoder_OFF4data_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_OFF4data_4\ : std_logic;
signal \frame_decoder_CH4data_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH4data_5\ : std_logic;
signal \frame_decoder_OFF4data_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH4data_6\ : std_logic;
signal \frame_decoder_OFF4data_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8\ : std_logic;
signal \scaler_4.N_905_i_l_ofxZ0\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_1_c_RNO_1\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal scaler_4_data_6 : std_logic;
signal \scaler_4.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\ : std_logic;
signal scaler_4_data_7 : std_logic;
signal \scaler_4.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\ : std_logic;
signal scaler_4_data_8 : std_logic;
signal \scaler_4.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\ : std_logic;
signal scaler_4_data_9 : std_logic;
signal \scaler_4.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\ : std_logic;
signal scaler_4_data_10 : std_logic;
signal \scaler_4.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\ : std_logic;
signal scaler_4_data_11 : std_logic;
signal \scaler_4.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\ : std_logic;
signal scaler_4_data_12 : std_logic;
signal \scaler_4.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\ : std_logic;
signal \scaler_4.un3_source_data_0_cry_8_c_RNIS918\ : std_logic;
signal scaler_4_data_13 : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \scaler_4.un2_source_data_0_cry_9\ : std_logic;
signal scaler_4_data_14 : std_logic;
signal \scaler_4.un2_source_data_0\ : std_logic;
signal \frame_decoder_OFF4data_0\ : std_logic;
signal \frame_decoder_CH4data_0\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_4\ : std_logic;
signal scaler_4_data_4 : std_logic;
signal \ppm_encoder_1.rudderZ0Z_4\ : std_logic;
signal scaler_4_data_5 : std_logic;
signal \ppm_encoder_1.rudderZ0Z_5\ : std_logic;
signal \ppm_encoder_1.pid_altitude_dv_0\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_7\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_12\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_11_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\ : std_logic;
signal \ppm_encoder_1.N_1014_0\ : std_logic;
signal \ppm_encoder_1.N_1014_i\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_0\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_1\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_2\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_1\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_3\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_2\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_4\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_3\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_5\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_4\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_5\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_7\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_6\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_7\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_8\ : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_9\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_8\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_10\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_9\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_11\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_10\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_11\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_12\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_13\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_14\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_15\ : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_16\ : std_logic;
signal \ppm_encoder_1.un1_counter_13_cry_17\ : std_logic;
signal \ppm_encoder_1.N_320_g\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_12\ : std_logic;
signal \ppm_encoder_1.rudderZ0Z_12\ : std_logic;
signal \uart_pc_sync.aux_2__0_Z0Z_0\ : std_logic;
signal \uart_pc_sync.aux_3__0_Z0Z_0\ : std_logic;
signal uart_input_drone_c : std_logic;
signal \uart_drone_sync.aux_0__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_1__0__0_0\ : std_logic;
signal \uart_drone_sync.aux_2__0__0_0\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_1_1_0\ : std_logic;
signal \Commands_frame_decoder.state_RNIQRI31Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.source_offset4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_8\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.source_CH4data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.source_CH2data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_4\ : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\ : std_logic;
signal \frame_decoder_OFF4data_7\ : std_logic;
signal \frame_decoder_CH4data_7\ : std_logic;
signal \scaler_4.un3_source_data_0_axb_7\ : std_logic;
signal \uart_drone.data_AuxZ0Z_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_2\ : std_logic;
signal \uart_drone.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.data_AuxZ0Z_5\ : std_logic;
signal \uart_drone.data_AuxZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \frame_decoder_CH3data_1\ : std_logic;
signal \frame_decoder_OFF3data_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_0\ : std_logic;
signal \frame_decoder_CH3data_2\ : std_logic;
signal \frame_decoder_OFF3data_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1\ : std_logic;
signal \frame_decoder_OFF3data_3\ : std_logic;
signal \frame_decoder_CH3data_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2\ : std_logic;
signal \frame_decoder_CH3data_4\ : std_logic;
signal \frame_decoder_OFF3data_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3\ : std_logic;
signal \frame_decoder_CH3data_5\ : std_logic;
signal \frame_decoder_OFF3data_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4\ : std_logic;
signal \frame_decoder_CH3data_6\ : std_logic;
signal \frame_decoder_OFF3data_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_axb_7\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8\ : std_logic;
signal \frame_decoder_OFF3data_7\ : std_logic;
signal \frame_decoder_CH3data_7\ : std_logic;
signal \scaler_3.N_893_i_l_ofxZ0\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_1_c_RNO_0\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal scaler_3_data_6 : std_logic;
signal \scaler_3.un2_source_data_0_cry_1\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\ : std_logic;
signal scaler_3_data_7 : std_logic;
signal \scaler_3.un2_source_data_0_cry_2\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_2_c_RNI780L\ : std_logic;
signal scaler_3_data_8 : std_logic;
signal \scaler_3.un2_source_data_0_cry_3\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\ : std_logic;
signal scaler_3_data_9 : std_logic;
signal \scaler_3.un2_source_data_0_cry_4\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\ : std_logic;
signal scaler_3_data_10 : std_logic;
signal \scaler_3.un2_source_data_0_cry_5\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\ : std_logic;
signal scaler_3_data_11 : std_logic;
signal \scaler_3.un2_source_data_0_cry_6\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\ : std_logic;
signal scaler_3_data_12 : std_logic;
signal \scaler_3.un2_source_data_0_cry_7\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_8\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\ : std_logic;
signal \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\ : std_logic;
signal scaler_3_data_13 : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \scaler_3.un2_source_data_0_cry_9\ : std_logic;
signal scaler_3_data_14 : std_logic;
signal \scaler_3.un2_source_data_0\ : std_logic;
signal scaler_3_data_5 : std_logic;
signal \debug_CH3_20A_c_0_g\ : std_logic;
signal \ppm_encoder_1.N_305\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_13\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\ : std_logic;
signal \ppm_encoder_1.throttleZ0Z_6\ : std_logic;
signal \ppm_encoder_1.elevatorZ0Z_6\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\ : std_logic;
signal \ppm_encoder_1.N_298_cascade_\ : std_logic;
signal \ppm_encoder_1.aileronZ0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_10_mux\ : std_logic;
signal \ppm_encoder_1.pulses2count_9_sn_N_7\ : std_logic;
signal \ppm_encoder_1.N_320\ : std_logic;
signal \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_14\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_16\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_16\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_17\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_17\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_18\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_18\ : std_logic;
signal \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_15\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_17\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_16\ : std_logic;
signal \ppm_encoder_1.counterZ0Z_18\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\ : std_logic;
signal \ppm_encoder_1.init_pulsesZ0Z_15\ : std_logic;
signal \ppm_encoder_1.CHOOSE_CHANNEL_159_d\ : std_logic;
signal \ppm_encoder_1.PPM_STATE_59_d\ : std_logic;
signal \ppm_encoder_1.pulses2countZ0Z_15\ : std_logic;
signal \uart_pc_sync.aux_1__0_Z0Z_0\ : std_logic;
signal uart_input_pc_c : std_logic;
signal \uart_pc_sync.aux_0__0_Z0Z_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_338\ : std_logic;
signal \Commands_frame_decoder.N_309_cascade_\ : std_logic;
signal uart_pc_data_7 : std_logic;
signal uart_pc_data_2 : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\ : std_logic;
signal uart_pc_data_5 : std_logic;
signal \Commands_frame_decoder.state_ns_0_a3_3_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.N_342\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.N_308_2\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_0\ : std_logic;
signal \Commands_frame_decoder.N_308_2_cascade_\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_1_0\ : std_logic;
signal \uart_drone.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_drone.stateZ0Z_0\ : std_logic;
signal uart_pc_data_0 : std_logic;
signal uart_pc_data_6 : std_logic;
signal \uart_drone.stateZ0Z_1\ : std_logic;
signal \uart_drone.state_srsts_i_0_2_cascade_\ : std_logic;
signal \uart_drone_sync.aux_3__0__0_0\ : std_logic;
signal uart_pc_data_3 : std_logic;
signal \Commands_frame_decoder.count_1_sqmuxa\ : std_logic;
signal \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\ : std_logic;
signal uart_pc_data_1 : std_logic;
signal \uart_pc.timer_Count_RNILR1B2Z0Z_2\ : std_logic;
signal uart_pc_data_4 : std_logic;
signal \uart_drone.data_Auxce_0_0_2\ : std_logic;
signal \uart_drone.data_Auxce_0_6\ : std_logic;
signal \uart_drone.data_Auxce_0_5\ : std_logic;
signal \uart_drone.data_Auxce_0_3\ : std_logic;
signal \uart_drone.timer_Count_RNIES9Q1Z0Z_2\ : std_logic;
signal \uart_drone.data_rdyc_1\ : std_logic;
signal \uart_drone.data_rdyc_1_0\ : std_logic;
signal \uart_pc.data_AuxZ0Z_6\ : std_logic;
signal \uart_pc.data_AuxZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\ : std_logic;
signal \uart_drone.data_Auxce_0_0_0\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT10lto13_1\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0\ : std_logic;
signal \dron_frame_decoder_1.WDT10lt14_0_cascade_\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\ : std_logic;
signal \dron_frame_decoder_1.stateZ0Z_2\ : std_logic;
signal \frame_decoder_OFF3data_0\ : std_logic;
signal \frame_decoder_CH3data_0\ : std_logic;
signal scaler_3_data_4 : std_logic;
signal \Commands_frame_decoder.source_offset3data_1_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.stateZ0Z_9\ : std_logic;
signal \bfn_10_11_0_\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_drone.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_4\ : std_logic;
signal uart_drone_data_rdy : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_2\ : std_logic;
signal \uart_drone.timer_CountZ1Z_2\ : std_logic;
signal \uart_drone.un1_state_2_0_a3_0\ : std_logic;
signal \Commands_frame_decoder.state_ns_i_a3_1_0_0\ : std_logic;
signal \uart_drone.N_126_li\ : std_logic;
signal \uart_drone.timer_Count_0_sqmuxa\ : std_logic;
signal \uart_drone.N_143_cascade_\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_3\ : std_logic;
signal \uart_pc.state_srsts_i_0_2\ : std_logic;
signal \uart_pc.N_145_cascade_\ : std_logic;
signal \uart_drone.timer_CountZ0Z_4\ : std_logic;
signal \uart_drone.timer_CountZ1Z_3\ : std_logic;
signal \uart_drone.N_145\ : std_logic;
signal \uart_drone.stateZ0Z_2\ : std_logic;
signal \uart_drone.N_144_1_cascade_\ : std_logic;
signal \uart_drone.N_144_1\ : std_logic;
signal \uart_drone.N_143\ : std_logic;
signal \uart_drone.stateZ0Z_4\ : std_logic;
signal \uart_pc.un1_state_2_0_cascade_\ : std_logic;
signal \uart_pc.data_AuxZ1Z_1\ : std_logic;
signal \uart_pc.data_Auxce_0_0_2\ : std_logic;
signal \uart_pc.data_AuxZ1Z_2\ : std_logic;
signal \uart_pc.data_AuxZ0Z_4\ : std_logic;
signal \uart_pc.data_AuxZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.WDT8lto13_1_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0_cascade_\ : std_logic;
signal \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\ : std_logic;
signal \Commands_frame_decoder.N_303_0\ : std_logic;
signal \Commands_frame_decoder.WDT8lt14_0\ : std_logic;
signal \Commands_frame_decoder.N_335\ : std_logic;
signal \Commands_frame_decoder.preinitZ0\ : std_logic;
signal \uart_pc.data_Auxce_0_6\ : std_logic;
signal \uart_pc.data_Auxce_0_1\ : std_logic;
signal \uart_pc.data_Auxce_0_0_4\ : std_logic;
signal \uart_drone.data_Auxce_0_1\ : std_logic;
signal \uart_pc.data_Auxce_0_5\ : std_logic;
signal \dron_frame_decoder_1.WDT10_0_i\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_0\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_1\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_0\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_2\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_1\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_3\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_2\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_4\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_3\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_5\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_4\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_5\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_7\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_6\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_7\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_8\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_9\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_8\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_10\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_9\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_11\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_10\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_12\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_11\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_12\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_14\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_13\ : std_logic;
signal \dron_frame_decoder_1.un1_WDT_cry_14\ : std_logic;
signal \dron_frame_decoder_1.WDTZ0Z_15\ : std_logic;
signal \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\ : std_logic;
signal \uart_pc.stateZ0Z_1\ : std_logic;
signal \uart_drone.timer_CountZ0Z_0\ : std_logic;
signal \uart_drone.timer_CountZ1Z_1\ : std_logic;
signal \uart_drone.timer_Count_RNO_0_0_1\ : std_logic;
signal \Commands_frame_decoder.CO0_cascade_\ : std_logic;
signal \Commands_frame_decoder.CO0\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_2\ : std_logic;
signal uart_pc_data_rdy : std_logic;
signal \Commands_frame_decoder.stateZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.count_RNIDLVE1Z0Z_2\ : std_logic;
signal \Commands_frame_decoder.countZ0Z_0\ : std_logic;
signal \uart_pc.stateZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.state_0_sqmuxa\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_0\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_1\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_0\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_2\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_1\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_3\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_2\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_4\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_3\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_5\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_4\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_5\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_7\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_6\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_7\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_8\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_9\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_8\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_10\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_9\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_11\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_10\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_12\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_11\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_12\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_14\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_13\ : std_logic;
signal \Commands_frame_decoder.un1_WDT_cry_14\ : std_logic;
signal \Commands_frame_decoder.WDTZ0Z_15\ : std_logic;
signal \Commands_frame_decoder.un1_state51_iZ0\ : std_logic;
signal \uart_pc.N_144_1\ : std_logic;
signal \uart_pc.data_rdyc_1\ : std_logic;
signal \uart_pc.stateZ0Z_3\ : std_logic;
signal \uart_pc.N_152\ : std_logic;
signal \uart_pc.CO0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_2\ : std_logic;
signal \uart_pc.bit_CountZ0Z_0\ : std_logic;
signal \uart_pc.un1_state_4_0\ : std_logic;
signal \uart_pc.un1_state_7_0\ : std_logic;
signal \uart_pc.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.data_AuxZ0Z_7\ : std_logic;
signal \debug_CH0_16A_c\ : std_logic;
signal \uart_drone.un1_state_2_0\ : std_logic;
signal \uart_drone.data_AuxZ0Z_4\ : std_logic;
signal \uart_drone.state_RNIOU0NZ0Z_4\ : std_logic;
signal \pid_alt.stateZ0Z_0\ : std_logic;
signal \pid_alt.state_0_0\ : std_logic;
signal \reset_module_System.reset6_15_cascade_\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \reset_module_System.countZ0Z_2\ : std_logic;
signal \reset_module_System.count_1_2\ : std_logic;
signal \reset_module_System.count_1_cry_1\ : std_logic;
signal \reset_module_System.countZ0Z_3\ : std_logic;
signal \reset_module_System.count_1_cry_2\ : std_logic;
signal \reset_module_System.count_1_cry_3\ : std_logic;
signal \reset_module_System.count_1_cry_4\ : std_logic;
signal \reset_module_System.countZ0Z_6\ : std_logic;
signal \reset_module_System.count_1_cry_5\ : std_logic;
signal \reset_module_System.count_1_cry_6\ : std_logic;
signal \reset_module_System.count_1_cry_7\ : std_logic;
signal \reset_module_System.count_1_cry_8\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \reset_module_System.count_1_cry_9\ : std_logic;
signal \reset_module_System.count_1_cry_10\ : std_logic;
signal \reset_module_System.count_1_cry_11\ : std_logic;
signal \reset_module_System.count_1_cry_12\ : std_logic;
signal \reset_module_System.count_1_cry_13\ : std_logic;
signal \reset_module_System.count_1_cry_14\ : std_logic;
signal \reset_module_System.count_1_cry_15\ : std_logic;
signal \reset_module_System.count_1_cry_16\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \reset_module_System.count_1_cry_17\ : std_logic;
signal \reset_module_System.count_1_cry_18\ : std_logic;
signal \reset_module_System.countZ0Z_20\ : std_logic;
signal \reset_module_System.count_1_cry_19\ : std_logic;
signal \reset_module_System.count_1_cry_20\ : std_logic;
signal \uart_pc.stateZ0Z_4\ : std_logic;
signal \uart_pc.state_srsts_0_0_0_cascade_\ : std_logic;
signal \uart_pc.stateZ0Z_0\ : std_logic;
signal \uart_pc.un1_state_2_0_a3_0\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_1\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_3\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_2\ : std_logic;
signal \uart_pc.un4_timer_Count_1_cry_3\ : std_logic;
signal \uart_pc.timer_CountZ1Z_3\ : std_logic;
signal \uart_pc.N_126_li\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_4\ : std_logic;
signal \uart_pc.timer_CountZ0Z_4\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_2\ : std_logic;
signal \uart_pc.timer_CountZ1Z_2\ : std_logic;
signal \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uart_pc.timer_CountZ1Z_1\ : std_logic;
signal \uart_pc.N_143\ : std_logic;
signal \uart_pc.timer_Count_0_sqmuxa\ : std_logic;
signal reset_system : std_logic;
signal \uart_pc.timer_CountZ0Z_0\ : std_logic;
signal \reset_module_System.countZ0Z_8\ : std_logic;
signal \reset_module_System.countZ0Z_7\ : std_logic;
signal \reset_module_System.countZ0Z_5\ : std_logic;
signal \reset_module_System.countZ0Z_9\ : std_logic;
signal \reset_module_System.countZ0Z_4\ : std_logic;
signal \reset_module_System.countZ0Z_18\ : std_logic;
signal \reset_module_System.countZ0Z_16\ : std_logic;
signal \reset_module_System.reset6_3_cascade_\ : std_logic;
signal \reset_module_System.reset6_13\ : std_logic;
signal \reset_module_System.countZ0Z_12\ : std_logic;
signal \reset_module_System.reset6_17_cascade_\ : std_logic;
signal \reset_module_System.reset6_19_cascade_\ : std_logic;
signal \reset_module_System.countZ0Z_0\ : std_logic;
signal \reset_module_System.reset6_15\ : std_logic;
signal \reset_module_System.count_1_1_cascade_\ : std_logic;
signal \reset_module_System.reset6_19\ : std_logic;
signal \reset_module_System.countZ0Z_1\ : std_logic;
signal \reset_module_System.countZ0Z_14\ : std_logic;
signal \reset_module_System.countZ0Z_11\ : std_logic;
signal \reset_module_System.countZ0Z_17\ : std_logic;
signal \reset_module_System.countZ0Z_10\ : std_logic;
signal \reset_module_System.reset6_14\ : std_logic;
signal \reset_module_System.countZ0Z_19\ : std_logic;
signal \reset_module_System.countZ0Z_15\ : std_logic;
signal \reset_module_System.countZ0Z_21\ : std_logic;
signal \reset_module_System.countZ0Z_13\ : std_logic;
signal \reset_module_System.reset6_11\ : std_logic;
signal \uart_pc.data_Auxce_0_3\ : std_logic;
signal \uart_pc.data_AuxZ0Z_3\ : std_logic;
signal \uart_drone.un1_state_7_0_cascade_\ : std_logic;
signal \uart_drone.un1_state_7_0\ : std_logic;
signal \uart_drone.CO0\ : std_logic;
signal \uart_drone.N_152\ : std_logic;
signal \uart_drone.un1_state_4_0\ : std_logic;
signal \uart_drone.stateZ0Z_3\ : std_logic;
signal \uart_drone.bit_CountZ0Z_2\ : std_logic;
signal \uart_drone.bit_CountZ0Z_1\ : std_logic;
signal \uart_drone.bit_CountZ0Z_0\ : std_logic;
signal \uart_drone.data_Auxce_0_0_4\ : std_logic;
signal \debug_CH3_20A_c\ : std_logic;
signal reset_system_g : std_logic;
signal \debug_CH3_20A_c_0\ : std_logic;
signal \uart_pc.data_Auxce_0_0_0\ : std_logic;
signal \debug_CH2_18A_c\ : std_logic;
signal \uart_pc.un1_state_2_0\ : std_logic;
signal \uart_pc.data_AuxZ1Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_system_c_g : std_logic;
signal \uart_pc.state_RNIEAGSZ0Z_4\ : std_logic;

signal clk_system_wire : std_logic;
signal uart_input_drone_wire : std_logic;
signal uart_input_pc_wire : std_logic;
signal \debug_CH2_18A_wire\ : std_logic;
signal \debug_CH0_16A_wire\ : std_logic;
signal \debug_CH6_5B_wire\ : std_logic;
signal \debug_CH1_0A_wire\ : std_logic;
signal \debug_CH5_31B_wire\ : std_logic;
signal \debug_CH4_2A_wire\ : std_logic;
signal ppm_output_wire : std_logic;
signal \debug_CH3_20A_wire\ : std_logic;
signal \pid_alt.un2_error_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    clk_system_wire <= clk_system;
    uart_input_drone_wire <= uart_input_drone;
    uart_input_pc_wire <= uart_input_pc;
    debug_CH2_18A <= \debug_CH2_18A_wire\;
    debug_CH0_16A <= \debug_CH0_16A_wire\;
    debug_CH6_5B <= \debug_CH6_5B_wire\;
    debug_CH1_0A <= \debug_CH1_0A_wire\;
    debug_CH5_31B <= \debug_CH5_31B_wire\;
    debug_CH4_2A <= \debug_CH4_2A_wire\;
    ppm_output <= ppm_output_wire;
    debug_CH3_20A <= \debug_CH3_20A_wire\;
    \pid_alt.un2_error_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_A_wire\ <= \N__14840\&\N__14867\&\N__14891\&\N__14915\&\N__14942\&\N__14969\&\N__14996\&\N__15023\&\N__14636\&\N__14666\&\N__14693\&\N__14722\&\N__14750\&\N__14777\&\N__14804\&\N__15362\;
    \pid_alt.un2_error_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__20501\&\N__16982\&\N__16970\&\N__20489\&\N__16772\&\N__14483\&\N__16958\&\N__16946\;
    \pid_alt.O_0_24\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_0_23\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_0_22\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_0_21\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_0_20\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_0_19\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_0_18\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_0_17\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_0_16\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_0_15\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_0_14\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_0_13\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_0_12\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_0_11\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_0_10\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_0_9\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_0_8\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_0_7\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_0_6\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_0_5\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_0_4\ <= \pid_alt.un2_error_mulonly_0_24_0_O_wire\(4);
    \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\ <= \N__14833\&\N__14860\&\N__14884\&\N__14908\&\N__14935\&\N__14965\&\N__14992\&\N__15019\&\N__14632\&\N__14662\&\N__14692\&\N__14723\&\N__14749\&\N__14776\&\N__14803\&\N__15358\;
    \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__21149\&\N__14567\&\N__14579\&\N__14471\&\N__14591\&\N__14606\&\N__14459\&\N__14144\;
    \pid_alt.O_24\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(24);
    \pid_alt.O_23\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(23);
    \pid_alt.O_22\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(22);
    \pid_alt.O_21\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(21);
    \pid_alt.O_20\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(20);
    \pid_alt.O_19\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(19);
    \pid_alt.O_18\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(18);
    \pid_alt.O_17\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(17);
    \pid_alt.O_16\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(16);
    \pid_alt.O_15\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(15);
    \pid_alt.O_14\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(14);
    \pid_alt.O_13\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(13);
    \pid_alt.O_12\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(12);
    \pid_alt.O_11\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(11);
    \pid_alt.O_10\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(10);
    \pid_alt.O_9\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(9);
    \pid_alt.O_8\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(8);
    \pid_alt.O_7\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(7);
    \pid_alt.O_6\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(6);
    \pid_alt.O_5\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(5);
    \pid_alt.O_4\ <= \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\(4);

    \pid_alt.un2_error_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28718\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28717\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_mulonly_0_24_0_O_wire\
        );

    \pid_alt.un2_error_1_mulonly_0_24_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28699\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28704\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pid_alt.un2_error_1_mulonly_0_24_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pid_alt.un2_error_1_mulonly_0_24_0_A_wire\,
            C => \pid_alt.un2_error_1_mulonly_0_24_0_C_wire\,
            B => \pid_alt.un2_error_1_mulonly_0_24_0_B_wire\,
            OHOLDTOP => '0',
            O => \pid_alt.un2_error_1_mulonly_0_24_0_O_wire\
        );

    \clk_system_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__37455\,
            GLOBALBUFFEROUTPUT => clk_system_c_g
        );

    \clk_system_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37457\,
            DIN => \N__37456\,
            DOUT => \N__37455\,
            PACKAGEPIN => clk_system_wire
        );

    \clk_system_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37457\,
            PADOUT => \N__37456\,
            PADIN => \N__37455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_drone_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37446\,
            DIN => \N__37445\,
            DOUT => \N__37444\,
            PACKAGEPIN => uart_input_drone_wire
        );

    \uart_input_drone_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37446\,
            PADOUT => \N__37445\,
            PADIN => \N__37444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_drone_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \uart_input_pc_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37437\,
            DIN => \N__37436\,
            DOUT => \N__37435\,
            PACKAGEPIN => uart_input_pc_wire
        );

    \uart_input_pc_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37437\,
            PADOUT => \N__37436\,
            PADIN => \N__37435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => uart_input_pc_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH2_18A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37428\,
            DIN => \N__37427\,
            DOUT => \N__37426\,
            PACKAGEPIN => \debug_CH2_18A_wire\
        );

    \debug_CH2_18A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37428\,
            PADOUT => \N__37427\,
            PADIN => \N__37426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH0_16A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37419\,
            DIN => \N__37418\,
            DOUT => \N__37417\,
            PACKAGEPIN => \debug_CH0_16A_wire\
        );

    \debug_CH0_16A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37419\,
            PADOUT => \N__37418\,
            PADIN => \N__37417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH6_5B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37410\,
            DIN => \N__37409\,
            DOUT => \N__37408\,
            PACKAGEPIN => \debug_CH6_5B_wire\
        );

    \debug_CH6_5B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37410\,
            PADOUT => \N__37409\,
            PADIN => \N__37408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH1_0A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37401\,
            DIN => \N__37400\,
            DOUT => \N__37399\,
            PACKAGEPIN => \debug_CH1_0A_wire\
        );

    \debug_CH1_0A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37401\,
            PADOUT => \N__37400\,
            PADIN => \N__37399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH5_31B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37392\,
            DIN => \N__37391\,
            DOUT => \N__37390\,
            PACKAGEPIN => \debug_CH5_31B_wire\
        );

    \debug_CH5_31B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37392\,
            PADOUT => \N__37391\,
            PADIN => \N__37390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH4_2A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37383\,
            DIN => \N__37382\,
            DOUT => \N__37381\,
            PACKAGEPIN => \debug_CH4_2A_wire\
        );

    \debug_CH4_2A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37383\,
            PADOUT => \N__37382\,
            PADIN => \N__37381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ppm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37374\,
            DIN => \N__37373\,
            DOUT => \N__37372\,
            PACKAGEPIN => ppm_output_wire
        );

    \ppm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37374\,
            PADOUT => \N__37373\,
            PADIN => \N__37372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24710\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \debug_CH3_20A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37365\,
            DIN => \N__37364\,
            DOUT => \N__37363\,
            PACKAGEPIN => \debug_CH3_20A_wire\
        );

    \debug_CH3_20A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37365\,
            PADOUT => \N__37364\,
            PADIN => \N__37363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36976\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__9045\ : CascadeMux
    port map (
            O => \N__37346\,
            I => \uart_drone.un1_state_7_0_cascade_\
        );

    \I__9044\ : CascadeMux
    port map (
            O => \N__37343\,
            I => \N__37340\
        );

    \I__9043\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__37337\,
            I => \uart_drone.un1_state_7_0\
        );

    \I__9041\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__37331\,
            I => \uart_drone.CO0\
        );

    \I__9039\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37322\
        );

    \I__9038\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37319\
        );

    \I__9037\ : InMux
    port map (
            O => \N__37326\,
            I => \N__37316\
        );

    \I__9036\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37313\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__37322\,
            I => \N__37310\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37307\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__37316\,
            I => \N__37304\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__37313\,
            I => \N__37299\
        );

    \I__9031\ : Span4Mux_h
    port map (
            O => \N__37310\,
            I => \N__37299\
        );

    \I__9030\ : Span4Mux_h
    port map (
            O => \N__37307\,
            I => \N__37296\
        );

    \I__9029\ : Odrv4
    port map (
            O => \N__37304\,
            I => \uart_drone.N_152\
        );

    \I__9028\ : Odrv4
    port map (
            O => \N__37299\,
            I => \uart_drone.N_152\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__37296\,
            I => \uart_drone.N_152\
        );

    \I__9026\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37283\
        );

    \I__9025\ : InMux
    port map (
            O => \N__37288\,
            I => \N__37278\
        );

    \I__9024\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37278\
        );

    \I__9023\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37275\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__37283\,
            I => \N__37272\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__37278\,
            I => \N__37267\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__37275\,
            I => \N__37267\
        );

    \I__9019\ : Span4Mux_v
    port map (
            O => \N__37272\,
            I => \N__37264\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__37267\,
            I => \N__37261\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__37264\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__9016\ : Odrv4
    port map (
            O => \N__37261\,
            I => \uart_drone.un1_state_4_0\
        );

    \I__9015\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37252\
        );

    \I__9014\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37248\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__37252\,
            I => \N__37244\
        );

    \I__9012\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37241\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__37248\,
            I => \N__37237\
        );

    \I__9010\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37233\
        );

    \I__9009\ : Span4Mux_v
    port map (
            O => \N__37244\,
            I => \N__37228\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__37241\,
            I => \N__37228\
        );

    \I__9007\ : CascadeMux
    port map (
            O => \N__37240\,
            I => \N__37223\
        );

    \I__9006\ : Span4Mux_h
    port map (
            O => \N__37237\,
            I => \N__37220\
        );

    \I__9005\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37217\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__37233\,
            I => \N__37212\
        );

    \I__9003\ : Span4Mux_h
    port map (
            O => \N__37228\,
            I => \N__37212\
        );

    \I__9002\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37209\
        );

    \I__9001\ : InMux
    port map (
            O => \N__37226\,
            I => \N__37204\
        );

    \I__9000\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37204\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__37220\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__37217\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__37212\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__37209\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__37204\,
            I => \uart_drone.stateZ0Z_3\
        );

    \I__8994\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37186\
        );

    \I__8993\ : InMux
    port map (
            O => \N__37192\,
            I => \N__37176\
        );

    \I__8992\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37176\
        );

    \I__8991\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37176\
        );

    \I__8990\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37176\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__37186\,
            I => \N__37171\
        );

    \I__8988\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37168\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37165\
        );

    \I__8986\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37162\
        );

    \I__8985\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37158\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__37171\,
            I => \N__37149\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__37168\,
            I => \N__37149\
        );

    \I__8982\ : Span4Mux_v
    port map (
            O => \N__37165\,
            I => \N__37149\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37149\
        );

    \I__8980\ : InMux
    port map (
            O => \N__37161\,
            I => \N__37146\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__37158\,
            I => \N__37143\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__37149\,
            I => \N__37140\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__37146\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__37143\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__37140\,
            I => \uart_drone.bit_CountZ0Z_2\
        );

    \I__8974\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37128\
        );

    \I__8973\ : CascadeMux
    port map (
            O => \N__37132\,
            I => \N__37123\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__37131\,
            I => \N__37120\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__37128\,
            I => \N__37114\
        );

    \I__8970\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37111\
        );

    \I__8969\ : InMux
    port map (
            O => \N__37126\,
            I => \N__37108\
        );

    \I__8968\ : InMux
    port map (
            O => \N__37123\,
            I => \N__37097\
        );

    \I__8967\ : InMux
    port map (
            O => \N__37120\,
            I => \N__37097\
        );

    \I__8966\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37097\
        );

    \I__8965\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37097\
        );

    \I__8964\ : InMux
    port map (
            O => \N__37117\,
            I => \N__37094\
        );

    \I__8963\ : Span4Mux_v
    port map (
            O => \N__37114\,
            I => \N__37087\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__37111\,
            I => \N__37087\
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__37108\,
            I => \N__37087\
        );

    \I__8960\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37082\
        );

    \I__8959\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37082\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__37097\,
            I => \N__37079\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__37094\,
            I => \N__37076\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__37087\,
            I => \N__37073\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__37082\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8954\ : Odrv12
    port map (
            O => \N__37079\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__37076\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__37073\,
            I => \uart_drone.bit_CountZ0Z_1\
        );

    \I__8951\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37052\
        );

    \I__8950\ : InMux
    port map (
            O => \N__37063\,
            I => \N__37052\
        );

    \I__8949\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37052\
        );

    \I__8948\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37052\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__37052\,
            I => \N__37047\
        );

    \I__8946\ : InMux
    port map (
            O => \N__37051\,
            I => \N__37044\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__37050\,
            I => \N__37038\
        );

    \I__8944\ : Span4Mux_v
    port map (
            O => \N__37047\,
            I => \N__37033\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37033\
        );

    \I__8942\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37030\
        );

    \I__8941\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37025\
        );

    \I__8940\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37022\
        );

    \I__8939\ : InMux
    port map (
            O => \N__37038\,
            I => \N__37019\
        );

    \I__8938\ : Span4Mux_h
    port map (
            O => \N__37033\,
            I => \N__37016\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__37013\
        );

    \I__8936\ : InMux
    port map (
            O => \N__37029\,
            I => \N__37010\
        );

    \I__8935\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37007\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__37025\,
            I => \N__37004\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__37022\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__37019\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__37016\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8930\ : Odrv12
    port map (
            O => \N__37013\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__37010\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__37007\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8927\ : Odrv12
    port map (
            O => \N__37004\,
            I => \uart_drone.bit_CountZ0Z_0\
        );

    \I__8926\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__36980\,
            I => \uart_drone.data_Auxce_0_0_4\
        );

    \I__8922\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36973\
        );

    \I__8921\ : IoInMux
    port map (
            O => \N__36976\,
            I => \N__36970\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__36973\,
            I => \N__36966\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__36970\,
            I => \N__36962\
        );

    \I__8918\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36959\
        );

    \I__8917\ : Span4Mux_v
    port map (
            O => \N__36966\,
            I => \N__36955\
        );

    \I__8916\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36952\
        );

    \I__8915\ : Span12Mux_s11_v
    port map (
            O => \N__36962\,
            I => \N__36949\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__36959\,
            I => \N__36946\
        );

    \I__8913\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36943\
        );

    \I__8912\ : Span4Mux_v
    port map (
            O => \N__36955\,
            I => \N__36939\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__36952\,
            I => \N__36936\
        );

    \I__8910\ : Span12Mux_h
    port map (
            O => \N__36949\,
            I => \N__36929\
        );

    \I__8909\ : Span12Mux_h
    port map (
            O => \N__36946\,
            I => \N__36929\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__36943\,
            I => \N__36929\
        );

    \I__8907\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36926\
        );

    \I__8906\ : Sp12to4
    port map (
            O => \N__36939\,
            I => \N__36921\
        );

    \I__8905\ : Span12Mux_v
    port map (
            O => \N__36936\,
            I => \N__36921\
        );

    \I__8904\ : Odrv12
    port map (
            O => \N__36929\,
            I => \debug_CH3_20A_c\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__36926\,
            I => \debug_CH3_20A_c\
        );

    \I__8902\ : Odrv12
    port map (
            O => \N__36921\,
            I => \debug_CH3_20A_c\
        );

    \I__8901\ : CascadeMux
    port map (
            O => \N__36914\,
            I => \N__36906\
        );

    \I__8900\ : CascadeMux
    port map (
            O => \N__36913\,
            I => \N__36903\
        );

    \I__8899\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36870\
        );

    \I__8898\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36867\
        );

    \I__8897\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36864\
        );

    \I__8896\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36851\
        );

    \I__8895\ : InMux
    port map (
            O => \N__36906\,
            I => \N__36851\
        );

    \I__8894\ : InMux
    port map (
            O => \N__36903\,
            I => \N__36851\
        );

    \I__8893\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36851\
        );

    \I__8892\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36851\
        );

    \I__8891\ : InMux
    port map (
            O => \N__36900\,
            I => \N__36851\
        );

    \I__8890\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36846\
        );

    \I__8889\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36846\
        );

    \I__8888\ : InMux
    port map (
            O => \N__36897\,
            I => \N__36843\
        );

    \I__8887\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36840\
        );

    \I__8886\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36837\
        );

    \I__8885\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36834\
        );

    \I__8884\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36831\
        );

    \I__8883\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36828\
        );

    \I__8882\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36825\
        );

    \I__8881\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36822\
        );

    \I__8880\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36817\
        );

    \I__8879\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36817\
        );

    \I__8878\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36814\
        );

    \I__8877\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36811\
        );

    \I__8876\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36808\
        );

    \I__8875\ : InMux
    port map (
            O => \N__36884\,
            I => \N__36805\
        );

    \I__8874\ : InMux
    port map (
            O => \N__36883\,
            I => \N__36802\
        );

    \I__8873\ : InMux
    port map (
            O => \N__36882\,
            I => \N__36799\
        );

    \I__8872\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36794\
        );

    \I__8871\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36794\
        );

    \I__8870\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36791\
        );

    \I__8869\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36788\
        );

    \I__8868\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36785\
        );

    \I__8867\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36782\
        );

    \I__8866\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36779\
        );

    \I__8865\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36774\
        );

    \I__8864\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36774\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__36870\,
            I => \N__36686\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__36867\,
            I => \N__36683\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__36864\,
            I => \N__36680\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__36851\,
            I => \N__36677\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__36846\,
            I => \N__36674\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__36843\,
            I => \N__36671\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36668\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__36837\,
            I => \N__36665\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__36834\,
            I => \N__36662\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__36831\,
            I => \N__36659\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36656\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__36825\,
            I => \N__36653\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__36822\,
            I => \N__36650\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__36817\,
            I => \N__36647\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36644\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__36811\,
            I => \N__36641\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__36808\,
            I => \N__36638\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__36805\,
            I => \N__36635\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__36802\,
            I => \N__36632\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__36799\,
            I => \N__36629\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__36794\,
            I => \N__36626\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36623\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36620\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36617\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__36782\,
            I => \N__36614\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__36779\,
            I => \N__36611\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__36774\,
            I => \N__36608\
        );

    \I__8836\ : SRMux
    port map (
            O => \N__36773\,
            I => \N__36383\
        );

    \I__8835\ : SRMux
    port map (
            O => \N__36772\,
            I => \N__36383\
        );

    \I__8834\ : SRMux
    port map (
            O => \N__36771\,
            I => \N__36383\
        );

    \I__8833\ : SRMux
    port map (
            O => \N__36770\,
            I => \N__36383\
        );

    \I__8832\ : SRMux
    port map (
            O => \N__36769\,
            I => \N__36383\
        );

    \I__8831\ : SRMux
    port map (
            O => \N__36768\,
            I => \N__36383\
        );

    \I__8830\ : SRMux
    port map (
            O => \N__36767\,
            I => \N__36383\
        );

    \I__8829\ : SRMux
    port map (
            O => \N__36766\,
            I => \N__36383\
        );

    \I__8828\ : SRMux
    port map (
            O => \N__36765\,
            I => \N__36383\
        );

    \I__8827\ : SRMux
    port map (
            O => \N__36764\,
            I => \N__36383\
        );

    \I__8826\ : SRMux
    port map (
            O => \N__36763\,
            I => \N__36383\
        );

    \I__8825\ : SRMux
    port map (
            O => \N__36762\,
            I => \N__36383\
        );

    \I__8824\ : SRMux
    port map (
            O => \N__36761\,
            I => \N__36383\
        );

    \I__8823\ : SRMux
    port map (
            O => \N__36760\,
            I => \N__36383\
        );

    \I__8822\ : SRMux
    port map (
            O => \N__36759\,
            I => \N__36383\
        );

    \I__8821\ : SRMux
    port map (
            O => \N__36758\,
            I => \N__36383\
        );

    \I__8820\ : SRMux
    port map (
            O => \N__36757\,
            I => \N__36383\
        );

    \I__8819\ : SRMux
    port map (
            O => \N__36756\,
            I => \N__36383\
        );

    \I__8818\ : SRMux
    port map (
            O => \N__36755\,
            I => \N__36383\
        );

    \I__8817\ : SRMux
    port map (
            O => \N__36754\,
            I => \N__36383\
        );

    \I__8816\ : SRMux
    port map (
            O => \N__36753\,
            I => \N__36383\
        );

    \I__8815\ : SRMux
    port map (
            O => \N__36752\,
            I => \N__36383\
        );

    \I__8814\ : SRMux
    port map (
            O => \N__36751\,
            I => \N__36383\
        );

    \I__8813\ : SRMux
    port map (
            O => \N__36750\,
            I => \N__36383\
        );

    \I__8812\ : SRMux
    port map (
            O => \N__36749\,
            I => \N__36383\
        );

    \I__8811\ : SRMux
    port map (
            O => \N__36748\,
            I => \N__36383\
        );

    \I__8810\ : SRMux
    port map (
            O => \N__36747\,
            I => \N__36383\
        );

    \I__8809\ : SRMux
    port map (
            O => \N__36746\,
            I => \N__36383\
        );

    \I__8808\ : SRMux
    port map (
            O => \N__36745\,
            I => \N__36383\
        );

    \I__8807\ : SRMux
    port map (
            O => \N__36744\,
            I => \N__36383\
        );

    \I__8806\ : SRMux
    port map (
            O => \N__36743\,
            I => \N__36383\
        );

    \I__8805\ : SRMux
    port map (
            O => \N__36742\,
            I => \N__36383\
        );

    \I__8804\ : SRMux
    port map (
            O => \N__36741\,
            I => \N__36383\
        );

    \I__8803\ : SRMux
    port map (
            O => \N__36740\,
            I => \N__36383\
        );

    \I__8802\ : SRMux
    port map (
            O => \N__36739\,
            I => \N__36383\
        );

    \I__8801\ : SRMux
    port map (
            O => \N__36738\,
            I => \N__36383\
        );

    \I__8800\ : SRMux
    port map (
            O => \N__36737\,
            I => \N__36383\
        );

    \I__8799\ : SRMux
    port map (
            O => \N__36736\,
            I => \N__36383\
        );

    \I__8798\ : SRMux
    port map (
            O => \N__36735\,
            I => \N__36383\
        );

    \I__8797\ : SRMux
    port map (
            O => \N__36734\,
            I => \N__36383\
        );

    \I__8796\ : SRMux
    port map (
            O => \N__36733\,
            I => \N__36383\
        );

    \I__8795\ : SRMux
    port map (
            O => \N__36732\,
            I => \N__36383\
        );

    \I__8794\ : SRMux
    port map (
            O => \N__36731\,
            I => \N__36383\
        );

    \I__8793\ : SRMux
    port map (
            O => \N__36730\,
            I => \N__36383\
        );

    \I__8792\ : SRMux
    port map (
            O => \N__36729\,
            I => \N__36383\
        );

    \I__8791\ : SRMux
    port map (
            O => \N__36728\,
            I => \N__36383\
        );

    \I__8790\ : SRMux
    port map (
            O => \N__36727\,
            I => \N__36383\
        );

    \I__8789\ : SRMux
    port map (
            O => \N__36726\,
            I => \N__36383\
        );

    \I__8788\ : SRMux
    port map (
            O => \N__36725\,
            I => \N__36383\
        );

    \I__8787\ : SRMux
    port map (
            O => \N__36724\,
            I => \N__36383\
        );

    \I__8786\ : SRMux
    port map (
            O => \N__36723\,
            I => \N__36383\
        );

    \I__8785\ : SRMux
    port map (
            O => \N__36722\,
            I => \N__36383\
        );

    \I__8784\ : SRMux
    port map (
            O => \N__36721\,
            I => \N__36383\
        );

    \I__8783\ : SRMux
    port map (
            O => \N__36720\,
            I => \N__36383\
        );

    \I__8782\ : SRMux
    port map (
            O => \N__36719\,
            I => \N__36383\
        );

    \I__8781\ : SRMux
    port map (
            O => \N__36718\,
            I => \N__36383\
        );

    \I__8780\ : SRMux
    port map (
            O => \N__36717\,
            I => \N__36383\
        );

    \I__8779\ : SRMux
    port map (
            O => \N__36716\,
            I => \N__36383\
        );

    \I__8778\ : SRMux
    port map (
            O => \N__36715\,
            I => \N__36383\
        );

    \I__8777\ : SRMux
    port map (
            O => \N__36714\,
            I => \N__36383\
        );

    \I__8776\ : SRMux
    port map (
            O => \N__36713\,
            I => \N__36383\
        );

    \I__8775\ : SRMux
    port map (
            O => \N__36712\,
            I => \N__36383\
        );

    \I__8774\ : SRMux
    port map (
            O => \N__36711\,
            I => \N__36383\
        );

    \I__8773\ : SRMux
    port map (
            O => \N__36710\,
            I => \N__36383\
        );

    \I__8772\ : SRMux
    port map (
            O => \N__36709\,
            I => \N__36383\
        );

    \I__8771\ : SRMux
    port map (
            O => \N__36708\,
            I => \N__36383\
        );

    \I__8770\ : SRMux
    port map (
            O => \N__36707\,
            I => \N__36383\
        );

    \I__8769\ : SRMux
    port map (
            O => \N__36706\,
            I => \N__36383\
        );

    \I__8768\ : SRMux
    port map (
            O => \N__36705\,
            I => \N__36383\
        );

    \I__8767\ : SRMux
    port map (
            O => \N__36704\,
            I => \N__36383\
        );

    \I__8766\ : SRMux
    port map (
            O => \N__36703\,
            I => \N__36383\
        );

    \I__8765\ : SRMux
    port map (
            O => \N__36702\,
            I => \N__36383\
        );

    \I__8764\ : SRMux
    port map (
            O => \N__36701\,
            I => \N__36383\
        );

    \I__8763\ : SRMux
    port map (
            O => \N__36700\,
            I => \N__36383\
        );

    \I__8762\ : SRMux
    port map (
            O => \N__36699\,
            I => \N__36383\
        );

    \I__8761\ : SRMux
    port map (
            O => \N__36698\,
            I => \N__36383\
        );

    \I__8760\ : SRMux
    port map (
            O => \N__36697\,
            I => \N__36383\
        );

    \I__8759\ : SRMux
    port map (
            O => \N__36696\,
            I => \N__36383\
        );

    \I__8758\ : SRMux
    port map (
            O => \N__36695\,
            I => \N__36383\
        );

    \I__8757\ : SRMux
    port map (
            O => \N__36694\,
            I => \N__36383\
        );

    \I__8756\ : SRMux
    port map (
            O => \N__36693\,
            I => \N__36383\
        );

    \I__8755\ : SRMux
    port map (
            O => \N__36692\,
            I => \N__36383\
        );

    \I__8754\ : SRMux
    port map (
            O => \N__36691\,
            I => \N__36383\
        );

    \I__8753\ : SRMux
    port map (
            O => \N__36690\,
            I => \N__36383\
        );

    \I__8752\ : SRMux
    port map (
            O => \N__36689\,
            I => \N__36383\
        );

    \I__8751\ : Glb2LocalMux
    port map (
            O => \N__36686\,
            I => \N__36383\
        );

    \I__8750\ : Glb2LocalMux
    port map (
            O => \N__36683\,
            I => \N__36383\
        );

    \I__8749\ : Glb2LocalMux
    port map (
            O => \N__36680\,
            I => \N__36383\
        );

    \I__8748\ : Glb2LocalMux
    port map (
            O => \N__36677\,
            I => \N__36383\
        );

    \I__8747\ : Glb2LocalMux
    port map (
            O => \N__36674\,
            I => \N__36383\
        );

    \I__8746\ : Glb2LocalMux
    port map (
            O => \N__36671\,
            I => \N__36383\
        );

    \I__8745\ : Glb2LocalMux
    port map (
            O => \N__36668\,
            I => \N__36383\
        );

    \I__8744\ : Glb2LocalMux
    port map (
            O => \N__36665\,
            I => \N__36383\
        );

    \I__8743\ : Glb2LocalMux
    port map (
            O => \N__36662\,
            I => \N__36383\
        );

    \I__8742\ : Glb2LocalMux
    port map (
            O => \N__36659\,
            I => \N__36383\
        );

    \I__8741\ : Glb2LocalMux
    port map (
            O => \N__36656\,
            I => \N__36383\
        );

    \I__8740\ : Glb2LocalMux
    port map (
            O => \N__36653\,
            I => \N__36383\
        );

    \I__8739\ : Glb2LocalMux
    port map (
            O => \N__36650\,
            I => \N__36383\
        );

    \I__8738\ : Glb2LocalMux
    port map (
            O => \N__36647\,
            I => \N__36383\
        );

    \I__8737\ : Glb2LocalMux
    port map (
            O => \N__36644\,
            I => \N__36383\
        );

    \I__8736\ : Glb2LocalMux
    port map (
            O => \N__36641\,
            I => \N__36383\
        );

    \I__8735\ : Glb2LocalMux
    port map (
            O => \N__36638\,
            I => \N__36383\
        );

    \I__8734\ : Glb2LocalMux
    port map (
            O => \N__36635\,
            I => \N__36383\
        );

    \I__8733\ : Glb2LocalMux
    port map (
            O => \N__36632\,
            I => \N__36383\
        );

    \I__8732\ : Glb2LocalMux
    port map (
            O => \N__36629\,
            I => \N__36383\
        );

    \I__8731\ : Glb2LocalMux
    port map (
            O => \N__36626\,
            I => \N__36383\
        );

    \I__8730\ : Glb2LocalMux
    port map (
            O => \N__36623\,
            I => \N__36383\
        );

    \I__8729\ : Glb2LocalMux
    port map (
            O => \N__36620\,
            I => \N__36383\
        );

    \I__8728\ : Glb2LocalMux
    port map (
            O => \N__36617\,
            I => \N__36383\
        );

    \I__8727\ : Glb2LocalMux
    port map (
            O => \N__36614\,
            I => \N__36383\
        );

    \I__8726\ : Glb2LocalMux
    port map (
            O => \N__36611\,
            I => \N__36383\
        );

    \I__8725\ : Glb2LocalMux
    port map (
            O => \N__36608\,
            I => \N__36383\
        );

    \I__8724\ : GlobalMux
    port map (
            O => \N__36383\,
            I => \N__36380\
        );

    \I__8723\ : gio2CtrlBuf
    port map (
            O => \N__36380\,
            I => reset_system_g
        );

    \I__8722\ : IoInMux
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__8720\ : Odrv12
    port map (
            O => \N__36371\,
            I => \debug_CH3_20A_c_0\
        );

    \I__8719\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36365\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36362\
        );

    \I__8717\ : Span4Mux_h
    port map (
            O => \N__36362\,
            I => \N__36359\
        );

    \I__8716\ : Odrv4
    port map (
            O => \N__36359\,
            I => \uart_pc.data_Auxce_0_0_0\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__8714\ : InMux
    port map (
            O => \N__36353\,
            I => \N__36346\
        );

    \I__8713\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__8712\ : InMux
    port map (
            O => \N__36351\,
            I => \N__36340\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__36346\,
            I => \N__36335\
        );

    \I__8710\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36332\
        );

    \I__8709\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36329\
        );

    \I__8708\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36321\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36318\
        );

    \I__8706\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36315\
        );

    \I__8705\ : IoInMux
    port map (
            O => \N__36338\,
            I => \N__36311\
        );

    \I__8704\ : Span4Mux_h
    port map (
            O => \N__36335\,
            I => \N__36308\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__36332\,
            I => \N__36303\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36303\
        );

    \I__8701\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36294\
        );

    \I__8700\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36294\
        );

    \I__8699\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36294\
        );

    \I__8698\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36294\
        );

    \I__8697\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36291\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__36321\,
            I => \N__36284\
        );

    \I__8695\ : Span4Mux_v
    port map (
            O => \N__36318\,
            I => \N__36284\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36284\
        );

    \I__8693\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36281\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__36311\,
            I => \N__36278\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__36308\,
            I => \N__36275\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__36303\,
            I => \N__36270\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36270\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__36291\,
            I => \N__36263\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__36284\,
            I => \N__36263\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__36281\,
            I => \N__36263\
        );

    \I__8685\ : Span4Mux_s1_v
    port map (
            O => \N__36278\,
            I => \N__36260\
        );

    \I__8684\ : Sp12to4
    port map (
            O => \N__36275\,
            I => \N__36255\
        );

    \I__8683\ : Sp12to4
    port map (
            O => \N__36270\,
            I => \N__36255\
        );

    \I__8682\ : Sp12to4
    port map (
            O => \N__36263\,
            I => \N__36252\
        );

    \I__8681\ : Span4Mux_h
    port map (
            O => \N__36260\,
            I => \N__36249\
        );

    \I__8680\ : Span12Mux_v
    port map (
            O => \N__36255\,
            I => \N__36246\
        );

    \I__8679\ : Span12Mux_v
    port map (
            O => \N__36252\,
            I => \N__36243\
        );

    \I__8678\ : Odrv4
    port map (
            O => \N__36249\,
            I => \debug_CH2_18A_c\
        );

    \I__8677\ : Odrv12
    port map (
            O => \N__36246\,
            I => \debug_CH2_18A_c\
        );

    \I__8676\ : Odrv12
    port map (
            O => \N__36243\,
            I => \debug_CH2_18A_c\
        );

    \I__8675\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36231\
        );

    \I__8674\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36225\
        );

    \I__8673\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36225\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36222\
        );

    \I__8671\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36219\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36213\
        );

    \I__8669\ : Span4Mux_h
    port map (
            O => \N__36222\,
            I => \N__36208\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36208\
        );

    \I__8667\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36201\
        );

    \I__8666\ : InMux
    port map (
            O => \N__36217\,
            I => \N__36201\
        );

    \I__8665\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36201\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__36213\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8663\ : Odrv4
    port map (
            O => \N__36208\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__36201\,
            I => \uart_pc.un1_state_2_0\
        );

    \I__8661\ : CascadeMux
    port map (
            O => \N__36194\,
            I => \N__36191\
        );

    \I__8660\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36188\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36185\
        );

    \I__8658\ : Span4Mux_h
    port map (
            O => \N__36185\,
            I => \N__36181\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__8656\ : Span4Mux_h
    port map (
            O => \N__36181\,
            I => \N__36175\
        );

    \I__8655\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36172\
        );

    \I__8654\ : Odrv4
    port map (
            O => \N__36175\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__36172\,
            I => \uart_pc.data_AuxZ1Z_0\
        );

    \I__8652\ : ClkMux
    port map (
            O => \N__36167\,
            I => \N__35690\
        );

    \I__8651\ : ClkMux
    port map (
            O => \N__36166\,
            I => \N__35690\
        );

    \I__8650\ : ClkMux
    port map (
            O => \N__36165\,
            I => \N__35690\
        );

    \I__8649\ : ClkMux
    port map (
            O => \N__36164\,
            I => \N__35690\
        );

    \I__8648\ : ClkMux
    port map (
            O => \N__36163\,
            I => \N__35690\
        );

    \I__8647\ : ClkMux
    port map (
            O => \N__36162\,
            I => \N__35690\
        );

    \I__8646\ : ClkMux
    port map (
            O => \N__36161\,
            I => \N__35690\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__36160\,
            I => \N__35690\
        );

    \I__8644\ : ClkMux
    port map (
            O => \N__36159\,
            I => \N__35690\
        );

    \I__8643\ : ClkMux
    port map (
            O => \N__36158\,
            I => \N__35690\
        );

    \I__8642\ : ClkMux
    port map (
            O => \N__36157\,
            I => \N__35690\
        );

    \I__8641\ : ClkMux
    port map (
            O => \N__36156\,
            I => \N__35690\
        );

    \I__8640\ : ClkMux
    port map (
            O => \N__36155\,
            I => \N__35690\
        );

    \I__8639\ : ClkMux
    port map (
            O => \N__36154\,
            I => \N__35690\
        );

    \I__8638\ : ClkMux
    port map (
            O => \N__36153\,
            I => \N__35690\
        );

    \I__8637\ : ClkMux
    port map (
            O => \N__36152\,
            I => \N__35690\
        );

    \I__8636\ : ClkMux
    port map (
            O => \N__36151\,
            I => \N__35690\
        );

    \I__8635\ : ClkMux
    port map (
            O => \N__36150\,
            I => \N__35690\
        );

    \I__8634\ : ClkMux
    port map (
            O => \N__36149\,
            I => \N__35690\
        );

    \I__8633\ : ClkMux
    port map (
            O => \N__36148\,
            I => \N__35690\
        );

    \I__8632\ : ClkMux
    port map (
            O => \N__36147\,
            I => \N__35690\
        );

    \I__8631\ : ClkMux
    port map (
            O => \N__36146\,
            I => \N__35690\
        );

    \I__8630\ : ClkMux
    port map (
            O => \N__36145\,
            I => \N__35690\
        );

    \I__8629\ : ClkMux
    port map (
            O => \N__36144\,
            I => \N__35690\
        );

    \I__8628\ : ClkMux
    port map (
            O => \N__36143\,
            I => \N__35690\
        );

    \I__8627\ : ClkMux
    port map (
            O => \N__36142\,
            I => \N__35690\
        );

    \I__8626\ : ClkMux
    port map (
            O => \N__36141\,
            I => \N__35690\
        );

    \I__8625\ : ClkMux
    port map (
            O => \N__36140\,
            I => \N__35690\
        );

    \I__8624\ : ClkMux
    port map (
            O => \N__36139\,
            I => \N__35690\
        );

    \I__8623\ : ClkMux
    port map (
            O => \N__36138\,
            I => \N__35690\
        );

    \I__8622\ : ClkMux
    port map (
            O => \N__36137\,
            I => \N__35690\
        );

    \I__8621\ : ClkMux
    port map (
            O => \N__36136\,
            I => \N__35690\
        );

    \I__8620\ : ClkMux
    port map (
            O => \N__36135\,
            I => \N__35690\
        );

    \I__8619\ : ClkMux
    port map (
            O => \N__36134\,
            I => \N__35690\
        );

    \I__8618\ : ClkMux
    port map (
            O => \N__36133\,
            I => \N__35690\
        );

    \I__8617\ : ClkMux
    port map (
            O => \N__36132\,
            I => \N__35690\
        );

    \I__8616\ : ClkMux
    port map (
            O => \N__36131\,
            I => \N__35690\
        );

    \I__8615\ : ClkMux
    port map (
            O => \N__36130\,
            I => \N__35690\
        );

    \I__8614\ : ClkMux
    port map (
            O => \N__36129\,
            I => \N__35690\
        );

    \I__8613\ : ClkMux
    port map (
            O => \N__36128\,
            I => \N__35690\
        );

    \I__8612\ : ClkMux
    port map (
            O => \N__36127\,
            I => \N__35690\
        );

    \I__8611\ : ClkMux
    port map (
            O => \N__36126\,
            I => \N__35690\
        );

    \I__8610\ : ClkMux
    port map (
            O => \N__36125\,
            I => \N__35690\
        );

    \I__8609\ : ClkMux
    port map (
            O => \N__36124\,
            I => \N__35690\
        );

    \I__8608\ : ClkMux
    port map (
            O => \N__36123\,
            I => \N__35690\
        );

    \I__8607\ : ClkMux
    port map (
            O => \N__36122\,
            I => \N__35690\
        );

    \I__8606\ : ClkMux
    port map (
            O => \N__36121\,
            I => \N__35690\
        );

    \I__8605\ : ClkMux
    port map (
            O => \N__36120\,
            I => \N__35690\
        );

    \I__8604\ : ClkMux
    port map (
            O => \N__36119\,
            I => \N__35690\
        );

    \I__8603\ : ClkMux
    port map (
            O => \N__36118\,
            I => \N__35690\
        );

    \I__8602\ : ClkMux
    port map (
            O => \N__36117\,
            I => \N__35690\
        );

    \I__8601\ : ClkMux
    port map (
            O => \N__36116\,
            I => \N__35690\
        );

    \I__8600\ : ClkMux
    port map (
            O => \N__36115\,
            I => \N__35690\
        );

    \I__8599\ : ClkMux
    port map (
            O => \N__36114\,
            I => \N__35690\
        );

    \I__8598\ : ClkMux
    port map (
            O => \N__36113\,
            I => \N__35690\
        );

    \I__8597\ : ClkMux
    port map (
            O => \N__36112\,
            I => \N__35690\
        );

    \I__8596\ : ClkMux
    port map (
            O => \N__36111\,
            I => \N__35690\
        );

    \I__8595\ : ClkMux
    port map (
            O => \N__36110\,
            I => \N__35690\
        );

    \I__8594\ : ClkMux
    port map (
            O => \N__36109\,
            I => \N__35690\
        );

    \I__8593\ : ClkMux
    port map (
            O => \N__36108\,
            I => \N__35690\
        );

    \I__8592\ : ClkMux
    port map (
            O => \N__36107\,
            I => \N__35690\
        );

    \I__8591\ : ClkMux
    port map (
            O => \N__36106\,
            I => \N__35690\
        );

    \I__8590\ : ClkMux
    port map (
            O => \N__36105\,
            I => \N__35690\
        );

    \I__8589\ : ClkMux
    port map (
            O => \N__36104\,
            I => \N__35690\
        );

    \I__8588\ : ClkMux
    port map (
            O => \N__36103\,
            I => \N__35690\
        );

    \I__8587\ : ClkMux
    port map (
            O => \N__36102\,
            I => \N__35690\
        );

    \I__8586\ : ClkMux
    port map (
            O => \N__36101\,
            I => \N__35690\
        );

    \I__8585\ : ClkMux
    port map (
            O => \N__36100\,
            I => \N__35690\
        );

    \I__8584\ : ClkMux
    port map (
            O => \N__36099\,
            I => \N__35690\
        );

    \I__8583\ : ClkMux
    port map (
            O => \N__36098\,
            I => \N__35690\
        );

    \I__8582\ : ClkMux
    port map (
            O => \N__36097\,
            I => \N__35690\
        );

    \I__8581\ : ClkMux
    port map (
            O => \N__36096\,
            I => \N__35690\
        );

    \I__8580\ : ClkMux
    port map (
            O => \N__36095\,
            I => \N__35690\
        );

    \I__8579\ : ClkMux
    port map (
            O => \N__36094\,
            I => \N__35690\
        );

    \I__8578\ : ClkMux
    port map (
            O => \N__36093\,
            I => \N__35690\
        );

    \I__8577\ : ClkMux
    port map (
            O => \N__36092\,
            I => \N__35690\
        );

    \I__8576\ : ClkMux
    port map (
            O => \N__36091\,
            I => \N__35690\
        );

    \I__8575\ : ClkMux
    port map (
            O => \N__36090\,
            I => \N__35690\
        );

    \I__8574\ : ClkMux
    port map (
            O => \N__36089\,
            I => \N__35690\
        );

    \I__8573\ : ClkMux
    port map (
            O => \N__36088\,
            I => \N__35690\
        );

    \I__8572\ : ClkMux
    port map (
            O => \N__36087\,
            I => \N__35690\
        );

    \I__8571\ : ClkMux
    port map (
            O => \N__36086\,
            I => \N__35690\
        );

    \I__8570\ : ClkMux
    port map (
            O => \N__36085\,
            I => \N__35690\
        );

    \I__8569\ : ClkMux
    port map (
            O => \N__36084\,
            I => \N__35690\
        );

    \I__8568\ : ClkMux
    port map (
            O => \N__36083\,
            I => \N__35690\
        );

    \I__8567\ : ClkMux
    port map (
            O => \N__36082\,
            I => \N__35690\
        );

    \I__8566\ : ClkMux
    port map (
            O => \N__36081\,
            I => \N__35690\
        );

    \I__8565\ : ClkMux
    port map (
            O => \N__36080\,
            I => \N__35690\
        );

    \I__8564\ : ClkMux
    port map (
            O => \N__36079\,
            I => \N__35690\
        );

    \I__8563\ : ClkMux
    port map (
            O => \N__36078\,
            I => \N__35690\
        );

    \I__8562\ : ClkMux
    port map (
            O => \N__36077\,
            I => \N__35690\
        );

    \I__8561\ : ClkMux
    port map (
            O => \N__36076\,
            I => \N__35690\
        );

    \I__8560\ : ClkMux
    port map (
            O => \N__36075\,
            I => \N__35690\
        );

    \I__8559\ : ClkMux
    port map (
            O => \N__36074\,
            I => \N__35690\
        );

    \I__8558\ : ClkMux
    port map (
            O => \N__36073\,
            I => \N__35690\
        );

    \I__8557\ : ClkMux
    port map (
            O => \N__36072\,
            I => \N__35690\
        );

    \I__8556\ : ClkMux
    port map (
            O => \N__36071\,
            I => \N__35690\
        );

    \I__8555\ : ClkMux
    port map (
            O => \N__36070\,
            I => \N__35690\
        );

    \I__8554\ : ClkMux
    port map (
            O => \N__36069\,
            I => \N__35690\
        );

    \I__8553\ : ClkMux
    port map (
            O => \N__36068\,
            I => \N__35690\
        );

    \I__8552\ : ClkMux
    port map (
            O => \N__36067\,
            I => \N__35690\
        );

    \I__8551\ : ClkMux
    port map (
            O => \N__36066\,
            I => \N__35690\
        );

    \I__8550\ : ClkMux
    port map (
            O => \N__36065\,
            I => \N__35690\
        );

    \I__8549\ : ClkMux
    port map (
            O => \N__36064\,
            I => \N__35690\
        );

    \I__8548\ : ClkMux
    port map (
            O => \N__36063\,
            I => \N__35690\
        );

    \I__8547\ : ClkMux
    port map (
            O => \N__36062\,
            I => \N__35690\
        );

    \I__8546\ : ClkMux
    port map (
            O => \N__36061\,
            I => \N__35690\
        );

    \I__8545\ : ClkMux
    port map (
            O => \N__36060\,
            I => \N__35690\
        );

    \I__8544\ : ClkMux
    port map (
            O => \N__36059\,
            I => \N__35690\
        );

    \I__8543\ : ClkMux
    port map (
            O => \N__36058\,
            I => \N__35690\
        );

    \I__8542\ : ClkMux
    port map (
            O => \N__36057\,
            I => \N__35690\
        );

    \I__8541\ : ClkMux
    port map (
            O => \N__36056\,
            I => \N__35690\
        );

    \I__8540\ : ClkMux
    port map (
            O => \N__36055\,
            I => \N__35690\
        );

    \I__8539\ : ClkMux
    port map (
            O => \N__36054\,
            I => \N__35690\
        );

    \I__8538\ : ClkMux
    port map (
            O => \N__36053\,
            I => \N__35690\
        );

    \I__8537\ : ClkMux
    port map (
            O => \N__36052\,
            I => \N__35690\
        );

    \I__8536\ : ClkMux
    port map (
            O => \N__36051\,
            I => \N__35690\
        );

    \I__8535\ : ClkMux
    port map (
            O => \N__36050\,
            I => \N__35690\
        );

    \I__8534\ : ClkMux
    port map (
            O => \N__36049\,
            I => \N__35690\
        );

    \I__8533\ : ClkMux
    port map (
            O => \N__36048\,
            I => \N__35690\
        );

    \I__8532\ : ClkMux
    port map (
            O => \N__36047\,
            I => \N__35690\
        );

    \I__8531\ : ClkMux
    port map (
            O => \N__36046\,
            I => \N__35690\
        );

    \I__8530\ : ClkMux
    port map (
            O => \N__36045\,
            I => \N__35690\
        );

    \I__8529\ : ClkMux
    port map (
            O => \N__36044\,
            I => \N__35690\
        );

    \I__8528\ : ClkMux
    port map (
            O => \N__36043\,
            I => \N__35690\
        );

    \I__8527\ : ClkMux
    port map (
            O => \N__36042\,
            I => \N__35690\
        );

    \I__8526\ : ClkMux
    port map (
            O => \N__36041\,
            I => \N__35690\
        );

    \I__8525\ : ClkMux
    port map (
            O => \N__36040\,
            I => \N__35690\
        );

    \I__8524\ : ClkMux
    port map (
            O => \N__36039\,
            I => \N__35690\
        );

    \I__8523\ : ClkMux
    port map (
            O => \N__36038\,
            I => \N__35690\
        );

    \I__8522\ : ClkMux
    port map (
            O => \N__36037\,
            I => \N__35690\
        );

    \I__8521\ : ClkMux
    port map (
            O => \N__36036\,
            I => \N__35690\
        );

    \I__8520\ : ClkMux
    port map (
            O => \N__36035\,
            I => \N__35690\
        );

    \I__8519\ : ClkMux
    port map (
            O => \N__36034\,
            I => \N__35690\
        );

    \I__8518\ : ClkMux
    port map (
            O => \N__36033\,
            I => \N__35690\
        );

    \I__8517\ : ClkMux
    port map (
            O => \N__36032\,
            I => \N__35690\
        );

    \I__8516\ : ClkMux
    port map (
            O => \N__36031\,
            I => \N__35690\
        );

    \I__8515\ : ClkMux
    port map (
            O => \N__36030\,
            I => \N__35690\
        );

    \I__8514\ : ClkMux
    port map (
            O => \N__36029\,
            I => \N__35690\
        );

    \I__8513\ : ClkMux
    port map (
            O => \N__36028\,
            I => \N__35690\
        );

    \I__8512\ : ClkMux
    port map (
            O => \N__36027\,
            I => \N__35690\
        );

    \I__8511\ : ClkMux
    port map (
            O => \N__36026\,
            I => \N__35690\
        );

    \I__8510\ : ClkMux
    port map (
            O => \N__36025\,
            I => \N__35690\
        );

    \I__8509\ : ClkMux
    port map (
            O => \N__36024\,
            I => \N__35690\
        );

    \I__8508\ : ClkMux
    port map (
            O => \N__36023\,
            I => \N__35690\
        );

    \I__8507\ : ClkMux
    port map (
            O => \N__36022\,
            I => \N__35690\
        );

    \I__8506\ : ClkMux
    port map (
            O => \N__36021\,
            I => \N__35690\
        );

    \I__8505\ : ClkMux
    port map (
            O => \N__36020\,
            I => \N__35690\
        );

    \I__8504\ : ClkMux
    port map (
            O => \N__36019\,
            I => \N__35690\
        );

    \I__8503\ : ClkMux
    port map (
            O => \N__36018\,
            I => \N__35690\
        );

    \I__8502\ : ClkMux
    port map (
            O => \N__36017\,
            I => \N__35690\
        );

    \I__8501\ : ClkMux
    port map (
            O => \N__36016\,
            I => \N__35690\
        );

    \I__8500\ : ClkMux
    port map (
            O => \N__36015\,
            I => \N__35690\
        );

    \I__8499\ : ClkMux
    port map (
            O => \N__36014\,
            I => \N__35690\
        );

    \I__8498\ : ClkMux
    port map (
            O => \N__36013\,
            I => \N__35690\
        );

    \I__8497\ : ClkMux
    port map (
            O => \N__36012\,
            I => \N__35690\
        );

    \I__8496\ : ClkMux
    port map (
            O => \N__36011\,
            I => \N__35690\
        );

    \I__8495\ : ClkMux
    port map (
            O => \N__36010\,
            I => \N__35690\
        );

    \I__8494\ : ClkMux
    port map (
            O => \N__36009\,
            I => \N__35690\
        );

    \I__8493\ : GlobalMux
    port map (
            O => \N__35690\,
            I => \N__35687\
        );

    \I__8492\ : gio2CtrlBuf
    port map (
            O => \N__35687\,
            I => clk_system_c_g
        );

    \I__8491\ : SRMux
    port map (
            O => \N__35684\,
            I => \N__35680\
        );

    \I__8490\ : SRMux
    port map (
            O => \N__35683\,
            I => \N__35676\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__35680\,
            I => \N__35672\
        );

    \I__8488\ : SRMux
    port map (
            O => \N__35679\,
            I => \N__35669\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__35676\,
            I => \N__35666\
        );

    \I__8486\ : SRMux
    port map (
            O => \N__35675\,
            I => \N__35663\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__35672\,
            I => \N__35660\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__35669\,
            I => \N__35657\
        );

    \I__8483\ : Span4Mux_v
    port map (
            O => \N__35666\,
            I => \N__35652\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__35663\,
            I => \N__35652\
        );

    \I__8481\ : Odrv4
    port map (
            O => \N__35660\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8480\ : Odrv12
    port map (
            O => \N__35657\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8479\ : Odrv4
    port map (
            O => \N__35652\,
            I => \uart_pc.state_RNIEAGSZ0Z_4\
        );

    \I__8478\ : InMux
    port map (
            O => \N__35645\,
            I => \N__35641\
        );

    \I__8477\ : InMux
    port map (
            O => \N__35644\,
            I => \N__35638\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35635\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__35638\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__35635\,
            I => \reset_module_System.countZ0Z_18\
        );

    \I__8473\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35626\
        );

    \I__8472\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35623\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__35626\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__35623\,
            I => \reset_module_System.countZ0Z_16\
        );

    \I__8469\ : CascadeMux
    port map (
            O => \N__35618\,
            I => \reset_module_System.reset6_3_cascade_\
        );

    \I__8468\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__35612\,
            I => \reset_module_System.reset6_13\
        );

    \I__8466\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35606\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__35606\,
            I => \N__35602\
        );

    \I__8464\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35599\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__35602\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__35599\,
            I => \reset_module_System.countZ0Z_12\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__35594\,
            I => \reset_module_System.reset6_17_cascade_\
        );

    \I__8460\ : CascadeMux
    port map (
            O => \N__35591\,
            I => \reset_module_System.reset6_19_cascade_\
        );

    \I__8459\ : CascadeMux
    port map (
            O => \N__35588\,
            I => \N__35582\
        );

    \I__8458\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35575\
        );

    \I__8457\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35575\
        );

    \I__8456\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35575\
        );

    \I__8455\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35572\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__35575\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__35572\,
            I => \reset_module_System.countZ0Z_0\
        );

    \I__8452\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35560\
        );

    \I__8451\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35560\
        );

    \I__8450\ : InMux
    port map (
            O => \N__35565\,
            I => \N__35557\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__35560\,
            I => \reset_module_System.reset6_15\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__35557\,
            I => \reset_module_System.reset6_15\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__35552\,
            I => \reset_module_System.count_1_1_cascade_\
        );

    \I__8446\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35544\
        );

    \I__8445\ : InMux
    port map (
            O => \N__35548\,
            I => \N__35539\
        );

    \I__8444\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35539\
        );

    \I__8443\ : LocalMux
    port map (
            O => \N__35544\,
            I => \reset_module_System.reset6_19\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__35539\,
            I => \reset_module_System.reset6_19\
        );

    \I__8441\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35529\
        );

    \I__8440\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35524\
        );

    \I__8439\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35524\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__35529\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__35524\,
            I => \reset_module_System.countZ0Z_1\
        );

    \I__8436\ : InMux
    port map (
            O => \N__35519\,
            I => \N__35515\
        );

    \I__8435\ : InMux
    port map (
            O => \N__35518\,
            I => \N__35512\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__35515\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__35512\,
            I => \reset_module_System.countZ0Z_14\
        );

    \I__8432\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35503\
        );

    \I__8431\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35500\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__35503\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__35500\,
            I => \reset_module_System.countZ0Z_11\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__35495\,
            I => \N__35492\
        );

    \I__8427\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35488\
        );

    \I__8426\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35485\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__35488\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__35485\,
            I => \reset_module_System.countZ0Z_17\
        );

    \I__8423\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35476\
        );

    \I__8422\ : InMux
    port map (
            O => \N__35479\,
            I => \N__35473\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__35476\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__35473\,
            I => \reset_module_System.countZ0Z_10\
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__8418\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35457\
        );

    \I__8417\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35457\
        );

    \I__8416\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35454\
        );

    \I__8415\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35451\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__35457\,
            I => \N__35448\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__35454\,
            I => \reset_module_System.reset6_14\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__35451\,
            I => \reset_module_System.reset6_14\
        );

    \I__8411\ : Odrv4
    port map (
            O => \N__35448\,
            I => \reset_module_System.reset6_14\
        );

    \I__8410\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35437\
        );

    \I__8409\ : InMux
    port map (
            O => \N__35440\,
            I => \N__35434\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__35437\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__35434\,
            I => \reset_module_System.countZ0Z_19\
        );

    \I__8406\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35425\
        );

    \I__8405\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35422\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__35425\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__35422\,
            I => \reset_module_System.countZ0Z_15\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__35417\,
            I => \N__35413\
        );

    \I__8401\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35410\
        );

    \I__8400\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35407\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__35410\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__35407\,
            I => \reset_module_System.countZ0Z_21\
        );

    \I__8397\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35398\
        );

    \I__8396\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35395\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__35398\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__35395\,
            I => \reset_module_System.countZ0Z_13\
        );

    \I__8393\ : InMux
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__35387\,
            I => \reset_module_System.reset6_11\
        );

    \I__8391\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35381\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__35381\,
            I => \N__35378\
        );

    \I__8389\ : Span4Mux_h
    port map (
            O => \N__35378\,
            I => \N__35375\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__35375\,
            I => \uart_pc.data_Auxce_0_3\
        );

    \I__8387\ : CascadeMux
    port map (
            O => \N__35372\,
            I => \N__35369\
        );

    \I__8386\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35362\
        );

    \I__8384\ : CascadeMux
    port map (
            O => \N__35365\,
            I => \N__35359\
        );

    \I__8383\ : Span4Mux_h
    port map (
            O => \N__35362\,
            I => \N__35356\
        );

    \I__8382\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35353\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__35356\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__35353\,
            I => \uart_pc.data_AuxZ0Z_3\
        );

    \I__8379\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__35345\,
            I => \N__35341\
        );

    \I__8377\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35338\
        );

    \I__8376\ : Span4Mux_h
    port map (
            O => \N__35341\,
            I => \N__35332\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__35338\,
            I => \N__35332\
        );

    \I__8374\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35329\
        );

    \I__8373\ : Sp12to4
    port map (
            O => \N__35332\,
            I => \N__35319\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__35329\,
            I => \N__35319\
        );

    \I__8371\ : InMux
    port map (
            O => \N__35328\,
            I => \N__35314\
        );

    \I__8370\ : InMux
    port map (
            O => \N__35327\,
            I => \N__35314\
        );

    \I__8369\ : InMux
    port map (
            O => \N__35326\,
            I => \N__35309\
        );

    \I__8368\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35309\
        );

    \I__8367\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35306\
        );

    \I__8366\ : Odrv12
    port map (
            O => \N__35319\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__35314\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__35309\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__35306\,
            I => \uart_pc.timer_CountZ1Z_3\
        );

    \I__8362\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35294\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__35294\,
            I => \N__35289\
        );

    \I__8360\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35284\
        );

    \I__8359\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35284\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__35289\,
            I => \N__35279\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__35284\,
            I => \N__35279\
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__35279\,
            I => \uart_pc.N_126_li\
        );

    \I__8355\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35273\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__35273\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_4\
        );

    \I__8353\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35265\
        );

    \I__8352\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35260\
        );

    \I__8351\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35257\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__35265\,
            I => \N__35253\
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__35264\,
            I => \N__35250\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__35263\,
            I => \N__35247\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__35260\,
            I => \N__35241\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__35257\,
            I => \N__35241\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__35256\,
            I => \N__35237\
        );

    \I__8344\ : Span4Mux_h
    port map (
            O => \N__35253\,
            I => \N__35233\
        );

    \I__8343\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35228\
        );

    \I__8342\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35228\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__35246\,
            I => \N__35225\
        );

    \I__8340\ : Span4Mux_h
    port map (
            O => \N__35241\,
            I => \N__35222\
        );

    \I__8339\ : InMux
    port map (
            O => \N__35240\,
            I => \N__35217\
        );

    \I__8338\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35217\
        );

    \I__8337\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35214\
        );

    \I__8336\ : Span4Mux_v
    port map (
            O => \N__35233\,
            I => \N__35209\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35209\
        );

    \I__8334\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35206\
        );

    \I__8333\ : Odrv4
    port map (
            O => \N__35222\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__35217\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__35214\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__8330\ : Odrv4
    port map (
            O => \N__35209\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__35206\,
            I => \uart_pc.timer_CountZ0Z_4\
        );

    \I__8328\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35192\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__35192\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_2\
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__8325\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__8324\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35179\
        );

    \I__8323\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35176\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__35179\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__35176\,
            I => \uart_pc.timer_CountZ1Z_2\
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__35171\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\
        );

    \I__8319\ : InMux
    port map (
            O => \N__35168\,
            I => \N__35164\
        );

    \I__8318\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35161\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__35164\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__35161\,
            I => \uart_pc.timer_CountZ1Z_1\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__35156\,
            I => \N__35149\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__35155\,
            I => \N__35146\
        );

    \I__8313\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35140\
        );

    \I__8312\ : InMux
    port map (
            O => \N__35153\,
            I => \N__35140\
        );

    \I__8311\ : InMux
    port map (
            O => \N__35152\,
            I => \N__35135\
        );

    \I__8310\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35135\
        );

    \I__8309\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35130\
        );

    \I__8308\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35130\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35127\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__35135\,
            I => \uart_pc.N_143\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__35130\,
            I => \uart_pc.N_143\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__35127\,
            I => \uart_pc.N_143\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__35120\,
            I => \N__35116\
        );

    \I__8302\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35109\
        );

    \I__8301\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35109\
        );

    \I__8300\ : CascadeMux
    port map (
            O => \N__35115\,
            I => \N__35105\
        );

    \I__8299\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35102\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__35109\,
            I => \N__35099\
        );

    \I__8297\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35094\
        );

    \I__8296\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35094\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__35102\,
            I => \N__35091\
        );

    \I__8294\ : Span4Mux_v
    port map (
            O => \N__35099\,
            I => \N__35084\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__35094\,
            I => \N__35084\
        );

    \I__8292\ : Span4Mux_h
    port map (
            O => \N__35091\,
            I => \N__35084\
        );

    \I__8291\ : Odrv4
    port map (
            O => \N__35084\,
            I => \uart_pc.timer_Count_0_sqmuxa\
        );

    \I__8290\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35072\
        );

    \I__8289\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35069\
        );

    \I__8288\ : IoInMux
    port map (
            O => \N__35079\,
            I => \N__35066\
        );

    \I__8287\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35060\
        );

    \I__8286\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35051\
        );

    \I__8285\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35048\
        );

    \I__8284\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35045\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__35072\,
            I => \N__35042\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__35069\,
            I => \N__35039\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35036\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__35065\,
            I => \N__35029\
        );

    \I__8279\ : CascadeMux
    port map (
            O => \N__35064\,
            I => \N__35026\
        );

    \I__8278\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35017\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__35060\,
            I => \N__35014\
        );

    \I__8276\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35011\
        );

    \I__8275\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35008\
        );

    \I__8274\ : InMux
    port map (
            O => \N__35057\,
            I => \N__34999\
        );

    \I__8273\ : InMux
    port map (
            O => \N__35056\,
            I => \N__34999\
        );

    \I__8272\ : InMux
    port map (
            O => \N__35055\,
            I => \N__34999\
        );

    \I__8271\ : InMux
    port map (
            O => \N__35054\,
            I => \N__34999\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__35051\,
            I => \N__34994\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__34994\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__35045\,
            I => \N__34991\
        );

    \I__8267\ : Span4Mux_v
    port map (
            O => \N__35042\,
            I => \N__34986\
        );

    \I__8266\ : Span4Mux_h
    port map (
            O => \N__35039\,
            I => \N__34986\
        );

    \I__8265\ : IoSpan4Mux
    port map (
            O => \N__35036\,
            I => \N__34983\
        );

    \I__8264\ : InMux
    port map (
            O => \N__35035\,
            I => \N__34980\
        );

    \I__8263\ : InMux
    port map (
            O => \N__35034\,
            I => \N__34975\
        );

    \I__8262\ : InMux
    port map (
            O => \N__35033\,
            I => \N__34975\
        );

    \I__8261\ : InMux
    port map (
            O => \N__35032\,
            I => \N__34972\
        );

    \I__8260\ : InMux
    port map (
            O => \N__35029\,
            I => \N__34969\
        );

    \I__8259\ : InMux
    port map (
            O => \N__35026\,
            I => \N__34966\
        );

    \I__8258\ : InMux
    port map (
            O => \N__35025\,
            I => \N__34963\
        );

    \I__8257\ : InMux
    port map (
            O => \N__35024\,
            I => \N__34960\
        );

    \I__8256\ : InMux
    port map (
            O => \N__35023\,
            I => \N__34955\
        );

    \I__8255\ : InMux
    port map (
            O => \N__35022\,
            I => \N__34955\
        );

    \I__8254\ : InMux
    port map (
            O => \N__35021\,
            I => \N__34952\
        );

    \I__8253\ : InMux
    port map (
            O => \N__35020\,
            I => \N__34949\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__34944\
        );

    \I__8251\ : Span4Mux_v
    port map (
            O => \N__35014\,
            I => \N__34944\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__34941\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__34938\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34931\
        );

    \I__8247\ : Span4Mux_v
    port map (
            O => \N__34994\,
            I => \N__34931\
        );

    \I__8246\ : Span4Mux_v
    port map (
            O => \N__34991\,
            I => \N__34931\
        );

    \I__8245\ : Span4Mux_h
    port map (
            O => \N__34986\,
            I => \N__34928\
        );

    \I__8244\ : Span4Mux_s3_v
    port map (
            O => \N__34983\,
            I => \N__34925\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__34980\,
            I => \N__34922\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__34975\,
            I => \N__34919\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34916\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34913\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34902\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__34963\,
            I => \N__34902\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__34960\,
            I => \N__34902\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__34955\,
            I => \N__34902\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__34952\,
            I => \N__34902\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34899\
        );

    \I__8233\ : Sp12to4
    port map (
            O => \N__34944\,
            I => \N__34894\
        );

    \I__8232\ : Span12Mux_s6_v
    port map (
            O => \N__34941\,
            I => \N__34894\
        );

    \I__8231\ : Span4Mux_v
    port map (
            O => \N__34938\,
            I => \N__34887\
        );

    \I__8230\ : Span4Mux_h
    port map (
            O => \N__34931\,
            I => \N__34887\
        );

    \I__8229\ : Span4Mux_h
    port map (
            O => \N__34928\,
            I => \N__34887\
        );

    \I__8228\ : Span4Mux_v
    port map (
            O => \N__34925\,
            I => \N__34884\
        );

    \I__8227\ : Span4Mux_v
    port map (
            O => \N__34922\,
            I => \N__34879\
        );

    \I__8226\ : Span4Mux_v
    port map (
            O => \N__34919\,
            I => \N__34879\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__34916\,
            I => \N__34874\
        );

    \I__8224\ : Span4Mux_h
    port map (
            O => \N__34913\,
            I => \N__34874\
        );

    \I__8223\ : Span4Mux_v
    port map (
            O => \N__34902\,
            I => \N__34869\
        );

    \I__8222\ : Span4Mux_h
    port map (
            O => \N__34899\,
            I => \N__34869\
        );

    \I__8221\ : Span12Mux_v
    port map (
            O => \N__34894\,
            I => \N__34866\
        );

    \I__8220\ : Span4Mux_v
    port map (
            O => \N__34887\,
            I => \N__34861\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__34884\,
            I => \N__34861\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__34879\,
            I => reset_system
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__34874\,
            I => reset_system
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__34869\,
            I => reset_system
        );

    \I__8215\ : Odrv12
    port map (
            O => \N__34866\,
            I => reset_system
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__34861\,
            I => reset_system
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34844\
        );

    \I__8212\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34841\
        );

    \I__8211\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34838\
        );

    \I__8210\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34833\
        );

    \I__8209\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34833\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__34841\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__34838\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__34833\,
            I => \uart_pc.timer_CountZ0Z_0\
        );

    \I__8205\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34822\
        );

    \I__8204\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34819\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__34822\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__34819\,
            I => \reset_module_System.countZ0Z_8\
        );

    \I__8201\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34810\
        );

    \I__8200\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34807\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__34810\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__34807\,
            I => \reset_module_System.countZ0Z_7\
        );

    \I__8197\ : CascadeMux
    port map (
            O => \N__34802\,
            I => \N__34799\
        );

    \I__8196\ : InMux
    port map (
            O => \N__34799\,
            I => \N__34795\
        );

    \I__8195\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34792\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34789\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__34792\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__34789\,
            I => \reset_module_System.countZ0Z_5\
        );

    \I__8191\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34780\
        );

    \I__8190\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34777\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__34780\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__34777\,
            I => \reset_module_System.countZ0Z_9\
        );

    \I__8187\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34768\
        );

    \I__8186\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34765\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__34768\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__34765\,
            I => \reset_module_System.countZ0Z_4\
        );

    \I__8183\ : InMux
    port map (
            O => \N__34760\,
            I => \reset_module_System.count_1_cry_20\
        );

    \I__8182\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34753\
        );

    \I__8181\ : CascadeMux
    port map (
            O => \N__34756\,
            I => \N__34748\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__34753\,
            I => \N__34743\
        );

    \I__8179\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34738\
        );

    \I__8178\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34738\
        );

    \I__8177\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34733\
        );

    \I__8176\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34733\
        );

    \I__8175\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34730\
        );

    \I__8174\ : Odrv4
    port map (
            O => \N__34743\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__34738\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__34733\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__34730\,
            I => \uart_pc.stateZ0Z_4\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__34721\,
            I => \uart_pc.state_srsts_0_0_0_cascade_\
        );

    \I__8169\ : CascadeMux
    port map (
            O => \N__34718\,
            I => \N__34715\
        );

    \I__8168\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__34709\,
            I => \N__34705\
        );

    \I__8165\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34702\
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__34705\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__34702\,
            I => \uart_pc.stateZ0Z_0\
        );

    \I__8162\ : CascadeMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__8161\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__8159\ : Span4Mux_h
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__34685\,
            I => \uart_pc.un1_state_2_0_a3_0\
        );

    \I__8157\ : InMux
    port map (
            O => \N__34682\,
            I => \uart_pc.un4_timer_Count_1_cry_1\
        );

    \I__8156\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__34676\,
            I => \uart_pc.timer_Count_RNO_0Z0Z_3\
        );

    \I__8154\ : InMux
    port map (
            O => \N__34673\,
            I => \uart_pc.un4_timer_Count_1_cry_2\
        );

    \I__8153\ : InMux
    port map (
            O => \N__34670\,
            I => \uart_pc.un4_timer_Count_1_cry_3\
        );

    \I__8152\ : InMux
    port map (
            O => \N__34667\,
            I => \reset_module_System.count_1_cry_11\
        );

    \I__8151\ : InMux
    port map (
            O => \N__34664\,
            I => \reset_module_System.count_1_cry_12\
        );

    \I__8150\ : InMux
    port map (
            O => \N__34661\,
            I => \reset_module_System.count_1_cry_13\
        );

    \I__8149\ : InMux
    port map (
            O => \N__34658\,
            I => \reset_module_System.count_1_cry_14\
        );

    \I__8148\ : InMux
    port map (
            O => \N__34655\,
            I => \reset_module_System.count_1_cry_15\
        );

    \I__8147\ : InMux
    port map (
            O => \N__34652\,
            I => \bfn_12_15_0_\
        );

    \I__8146\ : InMux
    port map (
            O => \N__34649\,
            I => \reset_module_System.count_1_cry_17\
        );

    \I__8145\ : InMux
    port map (
            O => \N__34646\,
            I => \reset_module_System.count_1_cry_18\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__34643\,
            I => \N__34640\
        );

    \I__8143\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34636\
        );

    \I__8142\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34633\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34630\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__34633\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__8139\ : Odrv4
    port map (
            O => \N__34630\,
            I => \reset_module_System.countZ0Z_20\
        );

    \I__8138\ : InMux
    port map (
            O => \N__34625\,
            I => \reset_module_System.count_1_cry_19\
        );

    \I__8137\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34618\
        );

    \I__8136\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34615\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__34618\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__34615\,
            I => \reset_module_System.countZ0Z_3\
        );

    \I__8133\ : InMux
    port map (
            O => \N__34610\,
            I => \reset_module_System.count_1_cry_2\
        );

    \I__8132\ : InMux
    port map (
            O => \N__34607\,
            I => \reset_module_System.count_1_cry_3\
        );

    \I__8131\ : InMux
    port map (
            O => \N__34604\,
            I => \reset_module_System.count_1_cry_4\
        );

    \I__8130\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34597\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34594\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__34597\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__34594\,
            I => \reset_module_System.countZ0Z_6\
        );

    \I__8126\ : InMux
    port map (
            O => \N__34589\,
            I => \reset_module_System.count_1_cry_5\
        );

    \I__8125\ : InMux
    port map (
            O => \N__34586\,
            I => \reset_module_System.count_1_cry_6\
        );

    \I__8124\ : InMux
    port map (
            O => \N__34583\,
            I => \reset_module_System.count_1_cry_7\
        );

    \I__8123\ : InMux
    port map (
            O => \N__34580\,
            I => \bfn_12_14_0_\
        );

    \I__8122\ : InMux
    port map (
            O => \N__34577\,
            I => \reset_module_System.count_1_cry_9\
        );

    \I__8121\ : InMux
    port map (
            O => \N__34574\,
            I => \reset_module_System.count_1_cry_10\
        );

    \I__8120\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34567\
        );

    \I__8119\ : CascadeMux
    port map (
            O => \N__34570\,
            I => \N__34562\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__34567\,
            I => \N__34555\
        );

    \I__8117\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34552\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34549\
        );

    \I__8115\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34543\
        );

    \I__8114\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34540\
        );

    \I__8113\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34533\
        );

    \I__8112\ : InMux
    port map (
            O => \N__34559\,
            I => \N__34533\
        );

    \I__8111\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34533\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__34555\,
            I => \N__34530\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__34552\,
            I => \N__34525\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__34549\,
            I => \N__34525\
        );

    \I__8107\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34518\
        );

    \I__8106\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34518\
        );

    \I__8105\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34518\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__34543\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__34540\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__34533\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__34530\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8100\ : Odrv12
    port map (
            O => \N__34525\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__34518\,
            I => \uart_pc.bit_CountZ0Z_0\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__34505\,
            I => \N__34501\
        );

    \I__8097\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34494\
        );

    \I__8096\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34494\
        );

    \I__8095\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34491\
        );

    \I__8094\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34488\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__34494\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__34491\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__34488\,
            I => \uart_pc.un1_state_4_0\
        );

    \I__8090\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34475\
        );

    \I__8089\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34475\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__34475\,
            I => \uart_pc.un1_state_7_0\
        );

    \I__8087\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34468\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__34471\,
            I => \N__34463\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__34468\,
            I => \N__34459\
        );

    \I__8084\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34456\
        );

    \I__8083\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34453\
        );

    \I__8082\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34443\
        );

    \I__8081\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34443\
        );

    \I__8080\ : Span4Mux_h
    port map (
            O => \N__34459\,
            I => \N__34440\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__34456\,
            I => \N__34435\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__34453\,
            I => \N__34435\
        );

    \I__8077\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34430\
        );

    \I__8076\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34430\
        );

    \I__8075\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34427\
        );

    \I__8074\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34422\
        );

    \I__8073\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34422\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__34443\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__34440\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8070\ : Odrv12
    port map (
            O => \N__34435\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__34430\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__34427\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__34422\,
            I => \uart_pc.bit_CountZ0Z_1\
        );

    \I__8066\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34406\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__34406\,
            I => \N__34402\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__34405\,
            I => \N__34399\
        );

    \I__8063\ : Span4Mux_h
    port map (
            O => \N__34402\,
            I => \N__34396\
        );

    \I__8062\ : InMux
    port map (
            O => \N__34399\,
            I => \N__34393\
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__34396\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__34393\,
            I => \uart_drone.data_AuxZ0Z_7\
        );

    \I__8059\ : IoInMux
    port map (
            O => \N__34388\,
            I => \N__34385\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34382\
        );

    \I__8057\ : IoSpan4Mux
    port map (
            O => \N__34382\,
            I => \N__34374\
        );

    \I__8056\ : CascadeMux
    port map (
            O => \N__34381\,
            I => \N__34371\
        );

    \I__8055\ : CascadeMux
    port map (
            O => \N__34380\,
            I => \N__34368\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34365\
        );

    \I__8053\ : InMux
    port map (
            O => \N__34378\,
            I => \N__34359\
        );

    \I__8052\ : InMux
    port map (
            O => \N__34377\,
            I => \N__34356\
        );

    \I__8051\ : Span4Mux_s0_v
    port map (
            O => \N__34374\,
            I => \N__34353\
        );

    \I__8050\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34339\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34339\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34339\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34339\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34339\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34339\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__34359\,
            I => \N__34336\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__34356\,
            I => \N__34332\
        );

    \I__8042\ : Sp12to4
    port map (
            O => \N__34353\,
            I => \N__34328\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__34352\,
            I => \N__34325\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__34339\,
            I => \N__34318\
        );

    \I__8039\ : Span4Mux_h
    port map (
            O => \N__34336\,
            I => \N__34318\
        );

    \I__8038\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34315\
        );

    \I__8037\ : Span4Mux_h
    port map (
            O => \N__34332\,
            I => \N__34312\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34309\
        );

    \I__8035\ : Span12Mux_v
    port map (
            O => \N__34328\,
            I => \N__34306\
        );

    \I__8034\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34303\
        );

    \I__8033\ : InMux
    port map (
            O => \N__34324\,
            I => \N__34300\
        );

    \I__8032\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34297\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__34318\,
            I => \N__34294\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34315\,
            I => \N__34287\
        );

    \I__8029\ : Sp12to4
    port map (
            O => \N__34312\,
            I => \N__34287\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__34309\,
            I => \N__34287\
        );

    \I__8027\ : Odrv12
    port map (
            O => \N__34306\,
            I => \debug_CH0_16A_c\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__34303\,
            I => \debug_CH0_16A_c\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__34300\,
            I => \debug_CH0_16A_c\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__34297\,
            I => \debug_CH0_16A_c\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__34294\,
            I => \debug_CH0_16A_c\
        );

    \I__8022\ : Odrv12
    port map (
            O => \N__34287\,
            I => \debug_CH0_16A_c\
        );

    \I__8021\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34271\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__34271\,
            I => \N__34261\
        );

    \I__8019\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34258\
        );

    \I__8018\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34245\
        );

    \I__8017\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34245\
        );

    \I__8016\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34245\
        );

    \I__8015\ : InMux
    port map (
            O => \N__34266\,
            I => \N__34245\
        );

    \I__8014\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34245\
        );

    \I__8013\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34245\
        );

    \I__8012\ : Span4Mux_v
    port map (
            O => \N__34261\,
            I => \N__34240\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34258\,
            I => \N__34240\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__34245\,
            I => \N__34237\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__34240\,
            I => \N__34234\
        );

    \I__8008\ : Span4Mux_v
    port map (
            O => \N__34237\,
            I => \N__34231\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__34234\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__34231\,
            I => \uart_drone.un1_state_2_0\
        );

    \I__8005\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34223\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34220\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__34220\,
            I => \N__34216\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__34219\,
            I => \N__34213\
        );

    \I__8001\ : Span4Mux_v
    port map (
            O => \N__34216\,
            I => \N__34210\
        );

    \I__8000\ : InMux
    port map (
            O => \N__34213\,
            I => \N__34207\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__34210\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__34207\,
            I => \uart_drone.data_AuxZ0Z_4\
        );

    \I__7997\ : SRMux
    port map (
            O => \N__34202\,
            I => \N__34198\
        );

    \I__7996\ : SRMux
    port map (
            O => \N__34201\,
            I => \N__34195\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34192\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34189\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__34192\,
            I => \N__34186\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__34189\,
            I => \N__34183\
        );

    \I__7991\ : Span4Mux_h
    port map (
            O => \N__34186\,
            I => \N__34179\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__34183\,
            I => \N__34176\
        );

    \I__7989\ : SRMux
    port map (
            O => \N__34182\,
            I => \N__34173\
        );

    \I__7988\ : Odrv4
    port map (
            O => \N__34179\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__34176\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__34173\,
            I => \uart_drone.state_RNIOU0NZ0Z_4\
        );

    \I__7985\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34155\
        );

    \I__7984\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34144\
        );

    \I__7983\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34144\
        );

    \I__7982\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34144\
        );

    \I__7981\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34144\
        );

    \I__7980\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34144\
        );

    \I__7979\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34137\
        );

    \I__7978\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34137\
        );

    \I__7977\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34137\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__34155\,
            I => \N__34134\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__34144\,
            I => \N__34124\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34124\
        );

    \I__7973\ : Span4Mux_h
    port map (
            O => \N__34134\,
            I => \N__34121\
        );

    \I__7972\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34114\
        );

    \I__7971\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34114\
        );

    \I__7970\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34114\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__34130\,
            I => \N__34111\
        );

    \I__7968\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34108\
        );

    \I__7967\ : Span4Mux_v
    port map (
            O => \N__34124\,
            I => \N__34105\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__34121\,
            I => \N__34102\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__34114\,
            I => \N__34099\
        );

    \I__7964\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34096\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__34108\,
            I => \N__34091\
        );

    \I__7962\ : Span4Mux_v
    port map (
            O => \N__34105\,
            I => \N__34091\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__34102\,
            I => \N__34088\
        );

    \I__7960\ : Sp12to4
    port map (
            O => \N__34099\,
            I => \N__34083\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__34096\,
            I => \N__34083\
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__34091\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__34088\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7956\ : Odrv12
    port map (
            O => \N__34083\,
            I => \pid_alt.stateZ0Z_0\
        );

    \I__7955\ : IoInMux
    port map (
            O => \N__34076\,
            I => \N__34073\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__34073\,
            I => \N__34070\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__34070\,
            I => \pid_alt.state_0_0\
        );

    \I__7952\ : CascadeMux
    port map (
            O => \N__34067\,
            I => \reset_module_System.reset6_15_cascade_\
        );

    \I__7951\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34060\
        );

    \I__7950\ : InMux
    port map (
            O => \N__34063\,
            I => \N__34057\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__34060\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__34057\,
            I => \reset_module_System.countZ0Z_2\
        );

    \I__7947\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34049\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__34049\,
            I => \reset_module_System.count_1_2\
        );

    \I__7945\ : InMux
    port map (
            O => \N__34046\,
            I => \reset_module_System.count_1_cry_1\
        );

    \I__7944\ : InMux
    port map (
            O => \N__34043\,
            I => \N__34037\
        );

    \I__7943\ : InMux
    port map (
            O => \N__34042\,
            I => \N__34032\
        );

    \I__7942\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34032\
        );

    \I__7941\ : InMux
    port map (
            O => \N__34040\,
            I => \N__34029\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__34037\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__34032\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__34029\,
            I => \Commands_frame_decoder.WDTZ0Z_14\
        );

    \I__7937\ : InMux
    port map (
            O => \N__34022\,
            I => \Commands_frame_decoder.un1_WDT_cry_13\
        );

    \I__7936\ : InMux
    port map (
            O => \N__34019\,
            I => \Commands_frame_decoder.un1_WDT_cry_14\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__34012\
        );

    \I__7934\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34007\
        );

    \I__7933\ : InMux
    port map (
            O => \N__34012\,
            I => \N__34000\
        );

    \I__7932\ : InMux
    port map (
            O => \N__34011\,
            I => \N__34000\
        );

    \I__7931\ : InMux
    port map (
            O => \N__34010\,
            I => \N__34000\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__34007\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__34000\,
            I => \Commands_frame_decoder.WDTZ0Z_15\
        );

    \I__7928\ : SRMux
    port map (
            O => \N__33995\,
            I => \N__33992\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__33992\,
            I => \N__33988\
        );

    \I__7926\ : SRMux
    port map (
            O => \N__33991\,
            I => \N__33985\
        );

    \I__7925\ : Span4Mux_v
    port map (
            O => \N__33988\,
            I => \N__33980\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33980\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__33980\,
            I => \N__33977\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__33977\,
            I => \N__33974\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__33974\,
            I => \Commands_frame_decoder.un1_state51_iZ0\
        );

    \I__7920\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33967\
        );

    \I__7919\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33964\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33961\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__33964\,
            I => \uart_pc.N_144_1\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__33961\,
            I => \uart_pc.N_144_1\
        );

    \I__7915\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33950\
        );

    \I__7914\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33947\
        );

    \I__7913\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33944\
        );

    \I__7912\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33941\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__33950\,
            I => \N__33938\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__33947\,
            I => \N__33935\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__33944\,
            I => \N__33932\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__33941\,
            I => \N__33929\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__33938\,
            I => \N__33926\
        );

    \I__7906\ : Span4Mux_h
    port map (
            O => \N__33935\,
            I => \N__33923\
        );

    \I__7905\ : Span4Mux_h
    port map (
            O => \N__33932\,
            I => \N__33918\
        );

    \I__7904\ : Span4Mux_h
    port map (
            O => \N__33929\,
            I => \N__33918\
        );

    \I__7903\ : Odrv4
    port map (
            O => \N__33926\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__33923\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__7901\ : Odrv4
    port map (
            O => \N__33918\,
            I => \uart_pc.data_rdyc_1\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33908\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__33908\,
            I => \N__33898\
        );

    \I__7898\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33893\
        );

    \I__7897\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33893\
        );

    \I__7896\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33888\
        );

    \I__7895\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33888\
        );

    \I__7894\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33885\
        );

    \I__7893\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33882\
        );

    \I__7892\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33879\
        );

    \I__7891\ : Span4Mux_v
    port map (
            O => \N__33898\,
            I => \N__33874\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__33893\,
            I => \N__33874\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33871\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__33885\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__33882\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__33879\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__7885\ : Odrv4
    port map (
            O => \N__33874\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__33871\,
            I => \uart_pc.stateZ0Z_3\
        );

    \I__7883\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33854\
        );

    \I__7882\ : InMux
    port map (
            O => \N__33859\,
            I => \N__33851\
        );

    \I__7881\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33848\
        );

    \I__7880\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33845\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__33854\,
            I => \uart_pc.N_152\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__33851\,
            I => \uart_pc.N_152\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__33848\,
            I => \uart_pc.N_152\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__33845\,
            I => \uart_pc.N_152\
        );

    \I__7875\ : InMux
    port map (
            O => \N__33836\,
            I => \N__33833\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__33833\,
            I => \uart_pc.CO0\
        );

    \I__7873\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33821\
        );

    \I__7871\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33818\
        );

    \I__7870\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33815\
        );

    \I__7869\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33807\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__33821\,
            I => \N__33804\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33799\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__33815\,
            I => \N__33799\
        );

    \I__7865\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33792\
        );

    \I__7864\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33792\
        );

    \I__7863\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33792\
        );

    \I__7862\ : InMux
    port map (
            O => \N__33811\,
            I => \N__33787\
        );

    \I__7861\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33787\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__33807\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__33804\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__7858\ : Odrv12
    port map (
            O => \N__33799\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__33792\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__33787\,
            I => \uart_pc.bit_CountZ0Z_2\
        );

    \I__7855\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33772\
        );

    \I__7854\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33769\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__33772\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__33769\,
            I => \Commands_frame_decoder.WDTZ0Z_6\
        );

    \I__7851\ : InMux
    port map (
            O => \N__33764\,
            I => \Commands_frame_decoder.un1_WDT_cry_5\
        );

    \I__7850\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33757\
        );

    \I__7849\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33754\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__33757\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__33754\,
            I => \Commands_frame_decoder.WDTZ0Z_7\
        );

    \I__7846\ : InMux
    port map (
            O => \N__33749\,
            I => \Commands_frame_decoder.un1_WDT_cry_6\
        );

    \I__7845\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33742\
        );

    \I__7844\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33739\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__33742\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__33739\,
            I => \Commands_frame_decoder.WDTZ0Z_8\
        );

    \I__7841\ : InMux
    port map (
            O => \N__33734\,
            I => \bfn_11_16_0_\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \N__33727\
        );

    \I__7839\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33724\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33721\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__33724\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__33721\,
            I => \Commands_frame_decoder.WDTZ0Z_9\
        );

    \I__7835\ : InMux
    port map (
            O => \N__33716\,
            I => \Commands_frame_decoder.un1_WDT_cry_8\
        );

    \I__7834\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33709\
        );

    \I__7833\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33706\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__33709\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__33706\,
            I => \Commands_frame_decoder.WDTZ0Z_10\
        );

    \I__7830\ : InMux
    port map (
            O => \N__33701\,
            I => \Commands_frame_decoder.un1_WDT_cry_9\
        );

    \I__7829\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33693\
        );

    \I__7828\ : InMux
    port map (
            O => \N__33697\,
            I => \N__33688\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33688\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__33693\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__33688\,
            I => \Commands_frame_decoder.WDTZ0Z_11\
        );

    \I__7824\ : InMux
    port map (
            O => \N__33683\,
            I => \Commands_frame_decoder.un1_WDT_cry_10\
        );

    \I__7823\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33675\
        );

    \I__7822\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33670\
        );

    \I__7821\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33670\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__33675\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__33670\,
            I => \Commands_frame_decoder.WDTZ0Z_12\
        );

    \I__7818\ : InMux
    port map (
            O => \N__33665\,
            I => \Commands_frame_decoder.un1_WDT_cry_11\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__33662\,
            I => \N__33658\
        );

    \I__7816\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33655\
        );

    \I__7815\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33652\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__33655\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33652\,
            I => \Commands_frame_decoder.WDTZ0Z_13\
        );

    \I__7812\ : InMux
    port map (
            O => \N__33647\,
            I => \Commands_frame_decoder.un1_WDT_cry_12\
        );

    \I__7811\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33637\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33643\,
            I => \N__33634\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__33642\,
            I => \N__33625\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__33641\,
            I => \N__33618\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__33640\,
            I => \N__33614\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__33637\,
            I => \N__33609\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__33634\,
            I => \N__33606\
        );

    \I__7804\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33603\
        );

    \I__7803\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33600\
        );

    \I__7802\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33597\
        );

    \I__7801\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33592\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33592\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33589\
        );

    \I__7798\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33580\
        );

    \I__7797\ : InMux
    port map (
            O => \N__33624\,
            I => \N__33580\
        );

    \I__7796\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33580\
        );

    \I__7795\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33580\
        );

    \I__7794\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33577\
        );

    \I__7793\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33570\
        );

    \I__7792\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33570\
        );

    \I__7791\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33570\
        );

    \I__7790\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33567\
        );

    \I__7789\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33564\
        );

    \I__7788\ : Span4Mux_h
    port map (
            O => \N__33609\,
            I => \N__33549\
        );

    \I__7787\ : Span4Mux_v
    port map (
            O => \N__33606\,
            I => \N__33549\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__33603\,
            I => \N__33549\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__33600\,
            I => \N__33549\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33549\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__33592\,
            I => \N__33546\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33543\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33538\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__33577\,
            I => \N__33538\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__33570\,
            I => \N__33535\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__33567\,
            I => \N__33530\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__33564\,
            I => \N__33530\
        );

    \I__7776\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33527\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33524\
        );

    \I__7774\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33519\
        );

    \I__7773\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33519\
        );

    \I__7772\ : Span4Mux_v
    port map (
            O => \N__33549\,
            I => \N__33514\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__33546\,
            I => \N__33514\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__33543\,
            I => \N__33507\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__33538\,
            I => \N__33507\
        );

    \I__7768\ : Span4Mux_h
    port map (
            O => \N__33535\,
            I => \N__33507\
        );

    \I__7767\ : Odrv4
    port map (
            O => \N__33530\,
            I => uart_pc_data_rdy
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__33527\,
            I => uart_pc_data_rdy
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33524\,
            I => uart_pc_data_rdy
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__33519\,
            I => uart_pc_data_rdy
        );

    \I__7763\ : Odrv4
    port map (
            O => \N__33514\,
            I => uart_pc_data_rdy
        );

    \I__7762\ : Odrv4
    port map (
            O => \N__33507\,
            I => uart_pc_data_rdy
        );

    \I__7761\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33485\
        );

    \I__7760\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33485\
        );

    \I__7759\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33482\
        );

    \I__7758\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33477\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33477\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33474\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__33482\,
            I => \N__33471\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__33477\,
            I => \N__33468\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__33474\,
            I => \N__33462\
        );

    \I__7752\ : Span4Mux_v
    port map (
            O => \N__33471\,
            I => \N__33462\
        );

    \I__7751\ : Span4Mux_h
    port map (
            O => \N__33468\,
            I => \N__33459\
        );

    \I__7750\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33456\
        );

    \I__7749\ : Odrv4
    port map (
            O => \N__33462\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__33459\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__33456\,
            I => \Commands_frame_decoder.stateZ0Z_11\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33440\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33448\,
            I => \N__33440\
        );

    \I__7744\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33440\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__33440\,
            I => \Commands_frame_decoder.count_RNIDLVE1Z0Z_2\
        );

    \I__7742\ : CascadeMux
    port map (
            O => \N__33437\,
            I => \N__33434\
        );

    \I__7741\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33428\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33428\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__33428\,
            I => \Commands_frame_decoder.countZ0Z_0\
        );

    \I__7738\ : CascadeMux
    port map (
            O => \N__33425\,
            I => \N__33421\
        );

    \I__7737\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33414\
        );

    \I__7736\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33414\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__33420\,
            I => \N__33411\
        );

    \I__7734\ : CascadeMux
    port map (
            O => \N__33419\,
            I => \N__33408\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__33414\,
            I => \N__33405\
        );

    \I__7732\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33402\
        );

    \I__7731\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33399\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__33405\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__33402\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__33399\,
            I => \uart_pc.stateZ0Z_2\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__33392\,
            I => \N__33388\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33385\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33382\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__33385\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__33382\,
            I => \Commands_frame_decoder.state_0_sqmuxa\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33374\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__33374\,
            I => \Commands_frame_decoder.WDTZ0Z_0\
        );

    \I__7720\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33368\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__33368\,
            I => \Commands_frame_decoder.WDTZ0Z_1\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33365\,
            I => \Commands_frame_decoder.un1_WDT_cry_0\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33359\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__33359\,
            I => \Commands_frame_decoder.WDTZ0Z_2\
        );

    \I__7715\ : InMux
    port map (
            O => \N__33356\,
            I => \Commands_frame_decoder.un1_WDT_cry_1\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33350\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33350\,
            I => \Commands_frame_decoder.WDTZ0Z_3\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33347\,
            I => \Commands_frame_decoder.un1_WDT_cry_2\
        );

    \I__7711\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33340\
        );

    \I__7710\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33337\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__33340\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__33337\,
            I => \Commands_frame_decoder.WDTZ0Z_4\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33332\,
            I => \Commands_frame_decoder.un1_WDT_cry_3\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33325\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33328\,
            I => \N__33322\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33325\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33322\,
            I => \Commands_frame_decoder.WDTZ0Z_5\
        );

    \I__7702\ : InMux
    port map (
            O => \N__33317\,
            I => \Commands_frame_decoder.un1_WDT_cry_4\
        );

    \I__7701\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33309\
        );

    \I__7700\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33304\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33304\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__33309\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__33304\,
            I => \dron_frame_decoder_1.WDTZ0Z_14\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33299\,
            I => \dron_frame_decoder_1.un1_WDT_cry_13\
        );

    \I__7695\ : InMux
    port map (
            O => \N__33296\,
            I => \dron_frame_decoder_1.un1_WDT_cry_14\
        );

    \I__7694\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33288\
        );

    \I__7693\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33283\
        );

    \I__7692\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33283\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__33288\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__33283\,
            I => \dron_frame_decoder_1.WDTZ0Z_15\
        );

    \I__7689\ : SRMux
    port map (
            O => \N__33278\,
            I => \N__33274\
        );

    \I__7688\ : SRMux
    port map (
            O => \N__33277\,
            I => \N__33271\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33268\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__33271\,
            I => \N__33265\
        );

    \I__7685\ : Span4Mux_v
    port map (
            O => \N__33268\,
            I => \N__33262\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__33265\,
            I => \N__33259\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__33262\,
            I => \N__33254\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__33259\,
            I => \N__33254\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__33254\,
            I => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__33251\,
            I => \N__33246\
        );

    \I__7679\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33243\
        );

    \I__7678\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33240\
        );

    \I__7677\ : InMux
    port map (
            O => \N__33246\,
            I => \N__33237\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33234\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__33240\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__33237\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__7673\ : Odrv12
    port map (
            O => \N__33234\,
            I => \uart_pc.stateZ0Z_1\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__33227\,
            I => \N__33221\
        );

    \I__7671\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33218\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33215\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33210\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33210\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__33218\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__33215\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33210\,
            I => \uart_drone.timer_CountZ0Z_0\
        );

    \I__7664\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33199\
        );

    \I__7663\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33196\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__33199\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33196\,
            I => \uart_drone.timer_CountZ1Z_1\
        );

    \I__7660\ : InMux
    port map (
            O => \N__33191\,
            I => \N__33188\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__33188\,
            I => \uart_drone.timer_Count_RNO_0_0_1\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__33185\,
            I => \Commands_frame_decoder.CO0_cascade_\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33179\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__33179\,
            I => \Commands_frame_decoder.CO0\
        );

    \I__7655\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33170\
        );

    \I__7654\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33170\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33170\,
            I => \Commands_frame_decoder.countZ0Z_1\
        );

    \I__7652\ : CascadeMux
    port map (
            O => \N__33167\,
            I => \N__33163\
        );

    \I__7651\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33160\
        );

    \I__7650\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33156\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33153\
        );

    \I__7648\ : CascadeMux
    port map (
            O => \N__33159\,
            I => \N__33150\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33144\
        );

    \I__7646\ : Span4Mux_v
    port map (
            O => \N__33153\,
            I => \N__33144\
        );

    \I__7645\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33139\
        );

    \I__7644\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33139\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__33144\,
            I => \Commands_frame_decoder.countZ0Z_2\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__33139\,
            I => \Commands_frame_decoder.countZ0Z_2\
        );

    \I__7641\ : InMux
    port map (
            O => \N__33134\,
            I => \dron_frame_decoder_1.un1_WDT_cry_4\
        );

    \I__7640\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33127\
        );

    \I__7639\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__33127\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__33124\,
            I => \dron_frame_decoder_1.WDTZ0Z_6\
        );

    \I__7636\ : InMux
    port map (
            O => \N__33119\,
            I => \dron_frame_decoder_1.un1_WDT_cry_5\
        );

    \I__7635\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33112\
        );

    \I__7634\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33109\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33112\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__33109\,
            I => \dron_frame_decoder_1.WDTZ0Z_7\
        );

    \I__7631\ : InMux
    port map (
            O => \N__33104\,
            I => \dron_frame_decoder_1.un1_WDT_cry_6\
        );

    \I__7630\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33097\
        );

    \I__7629\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33094\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__33097\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__33094\,
            I => \dron_frame_decoder_1.WDTZ0Z_8\
        );

    \I__7626\ : InMux
    port map (
            O => \N__33089\,
            I => \bfn_10_20_0_\
        );

    \I__7625\ : CascadeMux
    port map (
            O => \N__33086\,
            I => \N__33082\
        );

    \I__7624\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33079\
        );

    \I__7623\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33076\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__33079\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__33076\,
            I => \dron_frame_decoder_1.WDTZ0Z_9\
        );

    \I__7620\ : InMux
    port map (
            O => \N__33071\,
            I => \dron_frame_decoder_1.un1_WDT_cry_8\
        );

    \I__7619\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33064\
        );

    \I__7618\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33061\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__33064\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__33061\,
            I => \dron_frame_decoder_1.WDTZ0Z_10\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33056\,
            I => \dron_frame_decoder_1.un1_WDT_cry_9\
        );

    \I__7614\ : InMux
    port map (
            O => \N__33053\,
            I => \N__33048\
        );

    \I__7613\ : InMux
    port map (
            O => \N__33052\,
            I => \N__33045\
        );

    \I__7612\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33042\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__33048\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__33045\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__33042\,
            I => \dron_frame_decoder_1.WDTZ0Z_11\
        );

    \I__7608\ : InMux
    port map (
            O => \N__33035\,
            I => \dron_frame_decoder_1.un1_WDT_cry_10\
        );

    \I__7607\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33027\
        );

    \I__7606\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33024\
        );

    \I__7605\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33021\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__33027\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__33024\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__33021\,
            I => \dron_frame_decoder_1.WDTZ0Z_12\
        );

    \I__7601\ : InMux
    port map (
            O => \N__33014\,
            I => \dron_frame_decoder_1.un1_WDT_cry_11\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__33011\,
            I => \N__33007\
        );

    \I__7599\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33004\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33007\,
            I => \N__33001\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__33004\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__33001\,
            I => \dron_frame_decoder_1.WDTZ0Z_13\
        );

    \I__7595\ : InMux
    port map (
            O => \N__32996\,
            I => \dron_frame_decoder_1.un1_WDT_cry_12\
        );

    \I__7594\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32990\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__32990\,
            I => \N__32987\
        );

    \I__7592\ : Odrv4
    port map (
            O => \N__32987\,
            I => \uart_pc.data_Auxce_0_5\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__32984\,
            I => \N__32980\
        );

    \I__7590\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32977\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32980\,
            I => \N__32974\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__32977\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__32974\,
            I => \dron_frame_decoder_1.WDT10_0_i\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__32966\,
            I => \dron_frame_decoder_1.WDTZ0Z_0\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32960\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__32960\,
            I => \dron_frame_decoder_1.WDTZ0Z_1\
        );

    \I__7582\ : InMux
    port map (
            O => \N__32957\,
            I => \dron_frame_decoder_1.un1_WDT_cry_0\
        );

    \I__7581\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__32951\,
            I => \dron_frame_decoder_1.WDTZ0Z_2\
        );

    \I__7579\ : InMux
    port map (
            O => \N__32948\,
            I => \dron_frame_decoder_1.un1_WDT_cry_1\
        );

    \I__7578\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__32942\,
            I => \dron_frame_decoder_1.WDTZ0Z_3\
        );

    \I__7576\ : InMux
    port map (
            O => \N__32939\,
            I => \dron_frame_decoder_1.un1_WDT_cry_2\
        );

    \I__7575\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32932\
        );

    \I__7574\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32929\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__32932\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__32929\,
            I => \dron_frame_decoder_1.WDTZ0Z_4\
        );

    \I__7571\ : InMux
    port map (
            O => \N__32924\,
            I => \dron_frame_decoder_1.un1_WDT_cry_3\
        );

    \I__7570\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32917\
        );

    \I__7569\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32914\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__32917\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__32914\,
            I => \dron_frame_decoder_1.WDTZ0Z_5\
        );

    \I__7566\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32905\
        );

    \I__7565\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32902\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32897\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__32902\,
            I => \N__32897\
        );

    \I__7562\ : Span4Mux_h
    port map (
            O => \N__32897\,
            I => \N__32894\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__32894\,
            I => \Commands_frame_decoder.N_303_0\
        );

    \I__7560\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32885\
        );

    \I__7559\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32885\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__32885\,
            I => \Commands_frame_decoder.WDT8lt14_0\
        );

    \I__7557\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32876\
        );

    \I__7556\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32876\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32864\
        );

    \I__7554\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32857\
        );

    \I__7553\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32857\
        );

    \I__7552\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32857\
        );

    \I__7551\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32852\
        );

    \I__7550\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32852\
        );

    \I__7549\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32849\
        );

    \I__7548\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32842\
        );

    \I__7547\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32842\
        );

    \I__7546\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32842\
        );

    \I__7545\ : Sp12to4
    port map (
            O => \N__32864\,
            I => \N__32837\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32837\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__32852\,
            I => \N__32832\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32832\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__32842\,
            I => \N__32829\
        );

    \I__7540\ : Span12Mux_v
    port map (
            O => \N__32837\,
            I => \N__32826\
        );

    \I__7539\ : Span4Mux_v
    port map (
            O => \N__32832\,
            I => \N__32823\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__32829\,
            I => \N__32820\
        );

    \I__7537\ : Odrv12
    port map (
            O => \N__32826\,
            I => \Commands_frame_decoder.N_335\
        );

    \I__7536\ : Odrv4
    port map (
            O => \N__32823\,
            I => \Commands_frame_decoder.N_335\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__32820\,
            I => \Commands_frame_decoder.N_335\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__32813\,
            I => \N__32810\
        );

    \I__7533\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32807\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32802\
        );

    \I__7531\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32797\
        );

    \I__7530\ : InMux
    port map (
            O => \N__32805\,
            I => \N__32797\
        );

    \I__7529\ : Odrv12
    port map (
            O => \N__32802\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__32797\,
            I => \Commands_frame_decoder.preinitZ0\
        );

    \I__7527\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32789\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__32789\,
            I => \uart_pc.data_Auxce_0_6\
        );

    \I__7525\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32783\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__32783\,
            I => \N__32780\
        );

    \I__7523\ : Odrv4
    port map (
            O => \N__32780\,
            I => \uart_pc.data_Auxce_0_1\
        );

    \I__7522\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32774\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32774\,
            I => \N__32771\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__32771\,
            I => \uart_pc.data_Auxce_0_0_4\
        );

    \I__7519\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32765\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32762\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__32762\,
            I => \N__32759\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__32759\,
            I => \uart_drone.data_Auxce_0_1\
        );

    \I__7515\ : CascadeMux
    port map (
            O => \N__32756\,
            I => \uart_pc.un1_state_2_0_cascade_\
        );

    \I__7514\ : CascadeMux
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__7513\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32746\
        );

    \I__7512\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32743\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__32746\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__32743\,
            I => \uart_pc.data_AuxZ1Z_1\
        );

    \I__7509\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__32735\,
            I => \uart_pc.data_Auxce_0_0_2\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__7506\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32725\
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__32728\,
            I => \N__32722\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__32725\,
            I => \N__32719\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32716\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__32719\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__32716\,
            I => \uart_pc.data_AuxZ1Z_2\
        );

    \I__7500\ : CascadeMux
    port map (
            O => \N__32711\,
            I => \N__32707\
        );

    \I__7499\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32704\
        );

    \I__7498\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32701\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__32704\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__32701\,
            I => \uart_pc.data_AuxZ0Z_4\
        );

    \I__7495\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32692\
        );

    \I__7494\ : CascadeMux
    port map (
            O => \N__32695\,
            I => \N__32689\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__32692\,
            I => \N__32686\
        );

    \I__7492\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32683\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__32686\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__32683\,
            I => \uart_pc.data_AuxZ0Z_5\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \Commands_frame_decoder.WDT8lto13_1_cascade_\
        );

    \I__7488\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32672\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__32672\,
            I => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__32669\,
            I => \Commands_frame_decoder.WDT8lt14_0_cascade_\
        );

    \I__7485\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32663\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__32663\,
            I => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\
        );

    \I__7483\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32657\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__32657\,
            I => \uart_pc.state_srsts_i_0_2\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__32654\,
            I => \uart_pc.N_145_cascade_\
        );

    \I__7480\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32646\
        );

    \I__7479\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32637\
        );

    \I__7478\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32637\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__32646\,
            I => \N__32634\
        );

    \I__7476\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32629\
        );

    \I__7475\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32629\
        );

    \I__7474\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32624\
        );

    \I__7473\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32621\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__32637\,
            I => \N__32614\
        );

    \I__7471\ : Span4Mux_h
    port map (
            O => \N__32634\,
            I => \N__32614\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__32629\,
            I => \N__32614\
        );

    \I__7469\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32609\
        );

    \I__7468\ : InMux
    port map (
            O => \N__32627\,
            I => \N__32609\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__32624\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__32621\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__32614\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32609\,
            I => \uart_drone.timer_CountZ0Z_4\
        );

    \I__7463\ : InMux
    port map (
            O => \N__32600\,
            I => \N__32594\
        );

    \I__7462\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32591\
        );

    \I__7461\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32582\
        );

    \I__7460\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32582\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__32594\,
            I => \N__32579\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32576\
        );

    \I__7457\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32573\
        );

    \I__7456\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32568\
        );

    \I__7455\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32568\
        );

    \I__7454\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32565\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__32582\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7452\ : Odrv4
    port map (
            O => \N__32579\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__32576\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__32573\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__32568\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32565\,
            I => \uart_drone.timer_CountZ1Z_3\
        );

    \I__7447\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32549\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32546\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__32546\,
            I => \uart_drone.N_145\
        );

    \I__7444\ : CascadeMux
    port map (
            O => \N__32543\,
            I => \N__32539\
        );

    \I__7443\ : CascadeMux
    port map (
            O => \N__32542\,
            I => \N__32536\
        );

    \I__7442\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32531\
        );

    \I__7441\ : InMux
    port map (
            O => \N__32536\,
            I => \N__32528\
        );

    \I__7440\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32525\
        );

    \I__7439\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32522\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32517\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__32528\,
            I => \N__32517\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__32525\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__32522\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__32517\,
            I => \uart_drone.stateZ0Z_2\
        );

    \I__7433\ : CascadeMux
    port map (
            O => \N__32510\,
            I => \uart_drone.N_144_1_cascade_\
        );

    \I__7432\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__32504\,
            I => \uart_drone.N_144_1\
        );

    \I__7430\ : CascadeMux
    port map (
            O => \N__32501\,
            I => \N__32496\
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__32500\,
            I => \N__32493\
        );

    \I__7428\ : CascadeMux
    port map (
            O => \N__32499\,
            I => \N__32488\
        );

    \I__7427\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32479\
        );

    \I__7426\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32479\
        );

    \I__7425\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32479\
        );

    \I__7424\ : InMux
    port map (
            O => \N__32491\,
            I => \N__32479\
        );

    \I__7423\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32476\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__32479\,
            I => \uart_drone.N_143\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__32476\,
            I => \uart_drone.N_143\
        );

    \I__7420\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32468\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__32468\,
            I => \N__32461\
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__32467\,
            I => \N__32457\
        );

    \I__7417\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32454\
        );

    \I__7416\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32449\
        );

    \I__7415\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32449\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__32461\,
            I => \N__32446\
        );

    \I__7413\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32443\
        );

    \I__7412\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32440\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__32454\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__32449\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__32446\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__32443\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__32440\,
            I => \uart_drone.stateZ0Z_4\
        );

    \I__7406\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32426\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__32426\,
            I => \uart_drone.timer_Count_RNO_0_0_4\
        );

    \I__7404\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32418\
        );

    \I__7403\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32410\
        );

    \I__7402\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32407\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32403\
        );

    \I__7400\ : InMux
    port map (
            O => \N__32417\,
            I => \N__32400\
        );

    \I__7399\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32397\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32390\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32390\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32390\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32410\,
            I => \N__32384\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32384\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32381\
        );

    \I__7392\ : Span4Mux_v
    port map (
            O => \N__32403\,
            I => \N__32376\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32376\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32373\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__32390\,
            I => \N__32370\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32389\,
            I => \N__32367\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__32384\,
            I => \N__32364\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32357\
        );

    \I__7385\ : Span4Mux_v
    port map (
            O => \N__32376\,
            I => \N__32357\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__32373\,
            I => \N__32357\
        );

    \I__7383\ : Span4Mux_h
    port map (
            O => \N__32370\,
            I => \N__32353\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32350\
        );

    \I__7381\ : Span4Mux_h
    port map (
            O => \N__32364\,
            I => \N__32345\
        );

    \I__7380\ : Span4Mux_v
    port map (
            O => \N__32357\,
            I => \N__32345\
        );

    \I__7379\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32342\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__32353\,
            I => uart_drone_data_rdy
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__32350\,
            I => uart_drone_data_rdy
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__32345\,
            I => uart_drone_data_rdy
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32342\,
            I => uart_drone_data_rdy
        );

    \I__7374\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32330\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__32330\,
            I => \uart_drone.timer_Count_RNO_0_0_2\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32322\
        );

    \I__7371\ : InMux
    port map (
            O => \N__32326\,
            I => \N__32319\
        );

    \I__7370\ : InMux
    port map (
            O => \N__32325\,
            I => \N__32316\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32322\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__32319\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32316\,
            I => \uart_drone.timer_CountZ1Z_2\
        );

    \I__7366\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__32306\,
            I => \N__32303\
        );

    \I__7364\ : Odrv12
    port map (
            O => \N__32303\,
            I => \uart_drone.un1_state_2_0_a3_0\
        );

    \I__7363\ : CascadeMux
    port map (
            O => \N__32300\,
            I => \N__32297\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__32294\,
            I => \N__32291\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__32291\,
            I => \N__32287\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32284\
        );

    \I__7358\ : Odrv4
    port map (
            O => \N__32287\,
            I => \Commands_frame_decoder.state_ns_i_a3_1_0_0\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__32284\,
            I => \Commands_frame_decoder.state_ns_i_a3_1_0_0\
        );

    \I__7356\ : CascadeMux
    port map (
            O => \N__32279\,
            I => \N__32275\
        );

    \I__7355\ : InMux
    port map (
            O => \N__32278\,
            I => \N__32271\
        );

    \I__7354\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32266\
        );

    \I__7353\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32266\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__32271\,
            I => \uart_drone.N_126_li\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__32266\,
            I => \uart_drone.N_126_li\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__32261\,
            I => \N__32255\
        );

    \I__7349\ : CascadeMux
    port map (
            O => \N__32260\,
            I => \N__32252\
        );

    \I__7348\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32243\
        );

    \I__7347\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32243\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32243\
        );

    \I__7345\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32243\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__32243\,
            I => \N__32239\
        );

    \I__7343\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32236\
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__32239\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32236\,
            I => \uart_drone.timer_Count_0_sqmuxa\
        );

    \I__7340\ : CascadeMux
    port map (
            O => \N__32231\,
            I => \uart_drone.N_143_cascade_\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32222\
        );

    \I__7337\ : Odrv12
    port map (
            O => \N__32222\,
            I => \uart_drone.timer_Count_RNO_0_0_3\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32216\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__32216\,
            I => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\
        );

    \I__7334\ : CascadeMux
    port map (
            O => \N__32213\,
            I => \N__32210\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32207\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__32207\,
            I => \N__32203\
        );

    \I__7331\ : CascadeMux
    port map (
            O => \N__32206\,
            I => \N__32200\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__32203\,
            I => \N__32197\
        );

    \I__7329\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32194\
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__32197\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__32194\,
            I => \dron_frame_decoder_1.stateZ0Z_3\
        );

    \I__7326\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32179\
        );

    \I__7325\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32179\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32179\
        );

    \I__7323\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32175\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__32179\,
            I => \N__32171\
        );

    \I__7321\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32168\
        );

    \I__7320\ : LocalMux
    port map (
            O => \N__32175\,
            I => \N__32165\
        );

    \I__7319\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32162\
        );

    \I__7318\ : Span4Mux_h
    port map (
            O => \N__32171\,
            I => \N__32157\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32154\
        );

    \I__7316\ : Span4Mux_v
    port map (
            O => \N__32165\,
            I => \N__32149\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32162\,
            I => \N__32149\
        );

    \I__7314\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32146\
        );

    \I__7313\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32143\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__32157\,
            I => \N__32140\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__32154\,
            I => \N__32135\
        );

    \I__7310\ : Span4Mux_h
    port map (
            O => \N__32149\,
            I => \N__32135\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32146\,
            I => \N__32132\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__32143\,
            I => \N__32129\
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__32140\,
            I => \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\
        );

    \I__7306\ : Odrv4
    port map (
            O => \N__32135\,
            I => \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\
        );

    \I__7305\ : Odrv12
    port map (
            O => \N__32132\,
            I => \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\
        );

    \I__7304\ : Odrv4
    port map (
            O => \N__32129\,
            I => \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\
        );

    \I__7303\ : CascadeMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__7300\ : Span4Mux_h
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__32108\,
            I => \N__32104\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32107\,
            I => \N__32101\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__32104\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__32101\,
            I => \dron_frame_decoder_1.stateZ0Z_2\
        );

    \I__7295\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__32093\,
            I => \N__32087\
        );

    \I__7293\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32084\
        );

    \I__7292\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32081\
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__32090\,
            I => \N__32078\
        );

    \I__7290\ : Span4Mux_h
    port map (
            O => \N__32087\,
            I => \N__32071\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32084\,
            I => \N__32071\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__32081\,
            I => \N__32071\
        );

    \I__7287\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32068\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__32071\,
            I => \N__32063\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__32068\,
            I => \N__32063\
        );

    \I__7284\ : Odrv4
    port map (
            O => \N__32063\,
            I => \frame_decoder_OFF3data_0\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32060\,
            I => \N__32056\
        );

    \I__7282\ : InMux
    port map (
            O => \N__32059\,
            I => \N__32052\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__32049\
        );

    \I__7280\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32046\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__32052\,
            I => \N__32038\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__32049\,
            I => \N__32038\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__32046\,
            I => \N__32038\
        );

    \I__7276\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32035\
        );

    \I__7275\ : Span4Mux_v
    port map (
            O => \N__32038\,
            I => \N__32030\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32030\
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__32030\,
            I => \frame_decoder_CH3data_0\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32023\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__32026\,
            I => \N__32020\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__32023\,
            I => \N__32017\
        );

    \I__7269\ : InMux
    port map (
            O => \N__32020\,
            I => \N__32014\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__32017\,
            I => scaler_3_data_4
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__32014\,
            I => scaler_3_data_4
        );

    \I__7266\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32005\
        );

    \I__7265\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32002\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__32005\,
            I => \N__31999\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__32002\,
            I => \N__31996\
        );

    \I__7262\ : Span4Mux_v
    port map (
            O => \N__31999\,
            I => \N__31991\
        );

    \I__7261\ : Span4Mux_v
    port map (
            O => \N__31996\,
            I => \N__31991\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__31991\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa\
        );

    \I__7259\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31984\
        );

    \I__7258\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31981\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__31984\,
            I => \N__31978\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__31981\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__31978\,
            I => \Commands_frame_decoder.stateZ0Z_9\
        );

    \I__7254\ : InMux
    port map (
            O => \N__31973\,
            I => \uart_drone.un4_timer_Count_1_cry_1\
        );

    \I__7253\ : InMux
    port map (
            O => \N__31970\,
            I => \uart_drone.un4_timer_Count_1_cry_2\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31967\,
            I => \uart_drone.un4_timer_Count_1_cry_3\
        );

    \I__7251\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31960\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__31963\,
            I => \N__31957\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31954\
        );

    \I__7248\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31951\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__31954\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__31951\,
            I => \uart_pc.data_AuxZ0Z_6\
        );

    \I__7245\ : CascadeMux
    port map (
            O => \N__31946\,
            I => \N__31943\
        );

    \I__7244\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31940\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31936\
        );

    \I__7242\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31933\
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__31936\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31933\,
            I => \uart_pc.data_AuxZ0Z_7\
        );

    \I__7239\ : CEMux
    port map (
            O => \N__31928\,
            I => \N__31925\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__7237\ : Odrv4
    port map (
            O => \N__31922\,
            I => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\
        );

    \I__7236\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31916\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__31916\,
            I => \N__31913\
        );

    \I__7234\ : Odrv4
    port map (
            O => \N__31913\,
            I => \uart_drone.data_Auxce_0_0_0\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__31910\,
            I => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\
        );

    \I__7232\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31904\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__31904\,
            I => \dron_frame_decoder_1.WDT10lto13_1\
        );

    \I__7230\ : InMux
    port map (
            O => \N__31901\,
            I => \N__31898\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__31898\,
            I => \dron_frame_decoder_1.WDT10lt14_0\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \dron_frame_decoder_1.WDT10lt14_0_cascade_\
        );

    \I__7227\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31889\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__31889\,
            I => \N__31886\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__31883\,
            I => \Commands_frame_decoder.count_1_sqmuxa\
        );

    \I__7223\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31870\
        );

    \I__7222\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31870\
        );

    \I__7221\ : CascadeMux
    port map (
            O => \N__31878\,
            I => \N__31867\
        );

    \I__7220\ : InMux
    port map (
            O => \N__31877\,
            I => \N__31859\
        );

    \I__7219\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31859\
        );

    \I__7218\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31859\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31856\
        );

    \I__7216\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31851\
        );

    \I__7215\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31851\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31848\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__31856\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__31851\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__31848\,
            I => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\
        );

    \I__7210\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31836\
        );

    \I__7209\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31830\
        );

    \I__7208\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31830\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31824\
        );

    \I__7206\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31819\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31815\
        );

    \I__7204\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31812\
        );

    \I__7203\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31809\
        );

    \I__7202\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31806\
        );

    \I__7201\ : Span4Mux_h
    port map (
            O => \N__31824\,
            I => \N__31803\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31799\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31796\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__31819\,
            I => \N__31793\
        );

    \I__7197\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31790\
        );

    \I__7196\ : Span4Mux_h
    port map (
            O => \N__31815\,
            I => \N__31787\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__31812\,
            I => \N__31783\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__31809\,
            I => \N__31778\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__31806\,
            I => \N__31778\
        );

    \I__7192\ : Sp12to4
    port map (
            O => \N__31803\,
            I => \N__31775\
        );

    \I__7191\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31772\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__31799\,
            I => \N__31769\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__31796\,
            I => \N__31764\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__31793\,
            I => \N__31764\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__31790\,
            I => \N__31761\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__31787\,
            I => \N__31758\
        );

    \I__7185\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31755\
        );

    \I__7184\ : Span12Mux_s9_h
    port map (
            O => \N__31783\,
            I => \N__31752\
        );

    \I__7183\ : Span12Mux_v
    port map (
            O => \N__31778\,
            I => \N__31747\
        );

    \I__7182\ : Span12Mux_v
    port map (
            O => \N__31775\,
            I => \N__31747\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__31772\,
            I => \N__31736\
        );

    \I__7180\ : Span4Mux_v
    port map (
            O => \N__31769\,
            I => \N__31736\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__31764\,
            I => \N__31736\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__31761\,
            I => \N__31736\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__31758\,
            I => \N__31736\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__31755\,
            I => uart_pc_data_1
        );

    \I__7175\ : Odrv12
    port map (
            O => \N__31752\,
            I => uart_pc_data_1
        );

    \I__7174\ : Odrv12
    port map (
            O => \N__31747\,
            I => uart_pc_data_1
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__31736\,
            I => uart_pc_data_1
        );

    \I__7172\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31716\
        );

    \I__7171\ : InMux
    port map (
            O => \N__31726\,
            I => \N__31716\
        );

    \I__7170\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31711\
        );

    \I__7169\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31711\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31704\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31704\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31704\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__31716\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__31711\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__31704\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31692\
        );

    \I__7161\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31686\
        );

    \I__7160\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31683\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__31692\,
            I => \N__31680\
        );

    \I__7158\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31677\
        );

    \I__7157\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31674\
        );

    \I__7156\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31671\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31667\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__31683\,
            I => \N__31660\
        );

    \I__7153\ : Span4Mux_h
    port map (
            O => \N__31680\,
            I => \N__31660\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31660\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__31674\,
            I => \N__31655\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__31671\,
            I => \N__31655\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31648\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__31667\,
            I => \N__31643\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__31660\,
            I => \N__31643\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__31655\,
            I => \N__31640\
        );

    \I__7145\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31637\
        );

    \I__7144\ : CascadeMux
    port map (
            O => \N__31653\,
            I => \N__31633\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31652\,
            I => \N__31630\
        );

    \I__7142\ : InMux
    port map (
            O => \N__31651\,
            I => \N__31627\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31624\
        );

    \I__7140\ : Span4Mux_h
    port map (
            O => \N__31643\,
            I => \N__31619\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__31640\,
            I => \N__31619\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__31637\,
            I => \N__31616\
        );

    \I__7137\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31613\
        );

    \I__7136\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31610\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__31630\,
            I => \N__31607\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__31627\,
            I => \N__31602\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__31624\,
            I => \N__31602\
        );

    \I__7132\ : Sp12to4
    port map (
            O => \N__31619\,
            I => \N__31595\
        );

    \I__7131\ : Span12Mux_s9_h
    port map (
            O => \N__31616\,
            I => \N__31595\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__31613\,
            I => \N__31595\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__31610\,
            I => uart_pc_data_4
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__31607\,
            I => uart_pc_data_4
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__31602\,
            I => uart_pc_data_4
        );

    \I__7126\ : Odrv12
    port map (
            O => \N__31595\,
            I => uart_pc_data_4
        );

    \I__7125\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31583\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__31583\,
            I => \uart_drone.data_Auxce_0_0_2\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31577\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__31577\,
            I => \uart_drone.data_Auxce_0_6\
        );

    \I__7121\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31571\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__31571\,
            I => \uart_drone.data_Auxce_0_5\
        );

    \I__7119\ : InMux
    port map (
            O => \N__31568\,
            I => \N__31565\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__31565\,
            I => \uart_drone.data_Auxce_0_3\
        );

    \I__7117\ : SRMux
    port map (
            O => \N__31562\,
            I => \N__31559\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__31559\,
            I => \N__31556\
        );

    \I__7115\ : Span4Mux_h
    port map (
            O => \N__31556\,
            I => \N__31552\
        );

    \I__7114\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31549\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__31552\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__31549\,
            I => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__31541\,
            I => \N__31536\
        );

    \I__7109\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31533\
        );

    \I__7108\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31530\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__31536\,
            I => \N__31523\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__31533\,
            I => \N__31523\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31523\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__31523\,
            I => \uart_drone.data_rdyc_1\
        );

    \I__7103\ : CEMux
    port map (
            O => \N__31520\,
            I => \N__31517\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__31517\,
            I => \N__31514\
        );

    \I__7101\ : Odrv12
    port map (
            O => \N__31514\,
            I => \uart_drone.data_rdyc_1_0\
        );

    \I__7100\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31507\
        );

    \I__7099\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31504\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__31507\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__31504\,
            I => \uart_drone.stateZ0Z_0\
        );

    \I__7096\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31495\
        );

    \I__7095\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31487\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__31495\,
            I => \N__31484\
        );

    \I__7093\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31481\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31478\
        );

    \I__7091\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31471\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31468\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31465\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__31487\,
            I => \N__31462\
        );

    \I__7087\ : Span4Mux_h
    port map (
            O => \N__31484\,
            I => \N__31459\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__31481\,
            I => \N__31456\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31478\,
            I => \N__31453\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__31477\,
            I => \N__31450\
        );

    \I__7083\ : CascadeMux
    port map (
            O => \N__31476\,
            I => \N__31446\
        );

    \I__7082\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31442\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31474\,
            I => \N__31439\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__31471\,
            I => \N__31432\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31468\,
            I => \N__31432\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__31465\,
            I => \N__31432\
        );

    \I__7077\ : Span4Mux_h
    port map (
            O => \N__31462\,
            I => \N__31427\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__31459\,
            I => \N__31427\
        );

    \I__7075\ : Span4Mux_h
    port map (
            O => \N__31456\,
            I => \N__31422\
        );

    \I__7074\ : Span4Mux_h
    port map (
            O => \N__31453\,
            I => \N__31422\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31450\,
            I => \N__31419\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31449\,
            I => \N__31416\
        );

    \I__7071\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31410\
        );

    \I__7070\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31410\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__31442\,
            I => \N__31399\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31399\
        );

    \I__7067\ : Span4Mux_v
    port map (
            O => \N__31432\,
            I => \N__31399\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__31427\,
            I => \N__31399\
        );

    \I__7065\ : Span4Mux_v
    port map (
            O => \N__31422\,
            I => \N__31399\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__31419\,
            I => \N__31396\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__31416\,
            I => \N__31393\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31390\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31387\
        );

    \I__7060\ : Span4Mux_h
    port map (
            O => \N__31399\,
            I => \N__31380\
        );

    \I__7059\ : Span4Mux_v
    port map (
            O => \N__31396\,
            I => \N__31380\
        );

    \I__7058\ : Span4Mux_v
    port map (
            O => \N__31393\,
            I => \N__31380\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__31390\,
            I => uart_pc_data_0
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__31387\,
            I => uart_pc_data_0
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__31380\,
            I => uart_pc_data_0
        );

    \I__7054\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31370\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31366\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31363\
        );

    \I__7051\ : Span4Mux_h
    port map (
            O => \N__31366\,
            I => \N__31353\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__31363\,
            I => \N__31350\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31362\,
            I => \N__31347\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31344\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31340\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31337\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31334\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31331\
        );

    \I__7043\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31328\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__31353\,
            I => \N__31323\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__31350\,
            I => \N__31323\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31347\,
            I => \N__31318\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31344\,
            I => \N__31318\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31315\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__31340\,
            I => \N__31312\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31308\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__31334\,
            I => \N__31304\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31331\,
            I => \N__31299\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31299\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__31323\,
            I => \N__31296\
        );

    \I__7031\ : Span4Mux_v
    port map (
            O => \N__31318\,
            I => \N__31291\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__31315\,
            I => \N__31291\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__31312\,
            I => \N__31288\
        );

    \I__7028\ : InMux
    port map (
            O => \N__31311\,
            I => \N__31285\
        );

    \I__7027\ : Span12Mux_s9_h
    port map (
            O => \N__31308\,
            I => \N__31282\
        );

    \I__7026\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31279\
        );

    \I__7025\ : Span4Mux_h
    port map (
            O => \N__31304\,
            I => \N__31272\
        );

    \I__7024\ : Span4Mux_v
    port map (
            O => \N__31299\,
            I => \N__31272\
        );

    \I__7023\ : Span4Mux_h
    port map (
            O => \N__31296\,
            I => \N__31272\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__31291\,
            I => \N__31265\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__31288\,
            I => \N__31265\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__31285\,
            I => \N__31265\
        );

    \I__7019\ : Odrv12
    port map (
            O => \N__31282\,
            I => uart_pc_data_6
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__31279\,
            I => uart_pc_data_6
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__31272\,
            I => uart_pc_data_6
        );

    \I__7016\ : Odrv4
    port map (
            O => \N__31265\,
            I => uart_pc_data_6
        );

    \I__7015\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31251\
        );

    \I__7014\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31248\
        );

    \I__7013\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31243\
        );

    \I__7012\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31243\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__31248\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__31243\,
            I => \uart_drone.stateZ0Z_1\
        );

    \I__7009\ : CascadeMux
    port map (
            O => \N__31238\,
            I => \uart_drone.state_srsts_i_0_2_cascade_\
        );

    \I__7008\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31232\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__31232\,
            I => \N__31229\
        );

    \I__7006\ : Span4Mux_v
    port map (
            O => \N__31229\,
            I => \N__31226\
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__31226\,
            I => \uart_drone_sync.aux_3__0__0_0\
        );

    \I__7004\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31217\
        );

    \I__7003\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31214\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__31221\,
            I => \N__31211\
        );

    \I__7001\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31206\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__31217\,
            I => \N__31203\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__31214\,
            I => \N__31196\
        );

    \I__6998\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31191\
        );

    \I__6997\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31191\
        );

    \I__6996\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31188\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__31206\,
            I => \N__31185\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__31203\,
            I => \N__31182\
        );

    \I__6993\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31179\
        );

    \I__6992\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31176\
        );

    \I__6991\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31173\
        );

    \I__6990\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31170\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__31196\,
            I => \N__31165\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__31191\,
            I => \N__31165\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31162\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__31185\,
            I => \N__31159\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__31182\,
            I => \N__31149\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31149\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31149\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__31173\,
            I => \N__31149\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31144\
        );

    \I__6980\ : Span4Mux_v
    port map (
            O => \N__31165\,
            I => \N__31144\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__31162\,
            I => \N__31138\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__31159\,
            I => \N__31138\
        );

    \I__6977\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31135\
        );

    \I__6976\ : Span4Mux_v
    port map (
            O => \N__31149\,
            I => \N__31130\
        );

    \I__6975\ : Span4Mux_v
    port map (
            O => \N__31144\,
            I => \N__31130\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31143\,
            I => \N__31127\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__31138\,
            I => \N__31124\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__31135\,
            I => \N__31121\
        );

    \I__6971\ : Sp12to4
    port map (
            O => \N__31130\,
            I => \N__31118\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__31127\,
            I => uart_pc_data_3
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__31124\,
            I => uart_pc_data_3
        );

    \I__6968\ : Odrv12
    port map (
            O => \N__31121\,
            I => uart_pc_data_3
        );

    \I__6967\ : Odrv12
    port map (
            O => \N__31118\,
            I => uart_pc_data_3
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\
        );

    \I__6965\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__31103\,
            I => \N__31098\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31093\
        );

    \I__6962\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31093\
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__31098\,
            I => \Commands_frame_decoder.N_342\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__31093\,
            I => \Commands_frame_decoder.N_342\
        );

    \I__6959\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31085\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31080\
        );

    \I__6957\ : InMux
    port map (
            O => \N__31084\,
            I => \N__31073\
        );

    \I__6956\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31073\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__31080\,
            I => \N__31070\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31067\
        );

    \I__6953\ : InMux
    port map (
            O => \N__31078\,
            I => \N__31064\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__31073\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__6951\ : Odrv4
    port map (
            O => \N__31070\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__31067\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__31064\,
            I => \Commands_frame_decoder.stateZ0Z_1\
        );

    \I__6948\ : InMux
    port map (
            O => \N__31055\,
            I => \N__31052\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__6946\ : Odrv4
    port map (
            O => \N__31049\,
            I => \Commands_frame_decoder.N_308_2\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31042\
        );

    \I__6944\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31039\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__31042\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__31039\,
            I => \Commands_frame_decoder.stateZ0Z_0\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__31034\,
            I => \Commands_frame_decoder.N_308_2_cascade_\
        );

    \I__6940\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31028\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__31028\,
            I => \Commands_frame_decoder.state_ns_i_1_0\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__31025\,
            I => \uart_drone.state_srsts_0_0_0_cascade_\
        );

    \I__6937\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__31019\,
            I => \uart_pc_sync.aux_1__0_Z0Z_0\
        );

    \I__6935\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31013\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__31010\,
            I => uart_input_pc_c
        );

    \I__6932\ : InMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__31004\,
            I => \uart_pc_sync.aux_0__0_Z0Z_0\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__31001\,
            I => \Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__30995\,
            I => \Commands_frame_decoder.N_338\
        );

    \I__6927\ : CascadeMux
    port map (
            O => \N__30992\,
            I => \Commands_frame_decoder.N_309_cascade_\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30984\
        );

    \I__6925\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30978\
        );

    \I__6924\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30975\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30970\
        );

    \I__6922\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30966\
        );

    \I__6921\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30963\
        );

    \I__6920\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30960\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__30978\,
            I => \N__30954\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__30975\,
            I => \N__30951\
        );

    \I__6917\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30946\
        );

    \I__6916\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30946\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__30970\,
            I => \N__30942\
        );

    \I__6914\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30939\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30934\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__30963\,
            I => \N__30934\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__30960\,
            I => \N__30931\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30959\,
            I => \N__30928\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30925\
        );

    \I__6908\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30922\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__30954\,
            I => \N__30916\
        );

    \I__6906\ : Span4Mux_v
    port map (
            O => \N__30951\,
            I => \N__30916\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__30946\,
            I => \N__30913\
        );

    \I__6904\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30910\
        );

    \I__6903\ : Span4Mux_v
    port map (
            O => \N__30942\,
            I => \N__30905\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30905\
        );

    \I__6901\ : Span4Mux_v
    port map (
            O => \N__30934\,
            I => \N__30902\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__30931\,
            I => \N__30897\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__30928\,
            I => \N__30897\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__30925\,
            I => \N__30892\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30892\
        );

    \I__6896\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30889\
        );

    \I__6895\ : Span4Mux_h
    port map (
            O => \N__30916\,
            I => \N__30880\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__30913\,
            I => \N__30880\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__30910\,
            I => \N__30880\
        );

    \I__6892\ : Span4Mux_h
    port map (
            O => \N__30905\,
            I => \N__30880\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__30902\,
            I => uart_pc_data_7
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__30897\,
            I => uart_pc_data_7
        );

    \I__6889\ : Odrv12
    port map (
            O => \N__30892\,
            I => uart_pc_data_7
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__30889\,
            I => uart_pc_data_7
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__30880\,
            I => uart_pc_data_7
        );

    \I__6886\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30864\
        );

    \I__6885\ : InMux
    port map (
            O => \N__30868\,
            I => \N__30861\
        );

    \I__6884\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30858\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30847\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__30861\,
            I => \N__30847\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30841\
        );

    \I__6880\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30838\
        );

    \I__6879\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30835\
        );

    \I__6878\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30829\
        );

    \I__6877\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30829\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30825\
        );

    \I__6875\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30822\
        );

    \I__6874\ : Span4Mux_v
    port map (
            O => \N__30847\,
            I => \N__30818\
        );

    \I__6873\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30813\
        );

    \I__6872\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30813\
        );

    \I__6871\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30810\
        );

    \I__6870\ : Span4Mux_h
    port map (
            O => \N__30841\,
            I => \N__30805\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30805\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30802\
        );

    \I__6867\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30799\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__30829\,
            I => \N__30796\
        );

    \I__6865\ : InMux
    port map (
            O => \N__30828\,
            I => \N__30793\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N__30788\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__30822\,
            I => \N__30788\
        );

    \I__6862\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30785\
        );

    \I__6861\ : Sp12to4
    port map (
            O => \N__30818\,
            I => \N__30780\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30780\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__30810\,
            I => \N__30777\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__30805\,
            I => \N__30768\
        );

    \I__6857\ : Span4Mux_h
    port map (
            O => \N__30802\,
            I => \N__30768\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30768\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__30796\,
            I => \N__30768\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__30793\,
            I => \N__30759\
        );

    \I__6853\ : Sp12to4
    port map (
            O => \N__30788\,
            I => \N__30759\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__30785\,
            I => \N__30759\
        );

    \I__6851\ : Span12Mux_s8_h
    port map (
            O => \N__30780\,
            I => \N__30759\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__30777\,
            I => uart_pc_data_2
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__30768\,
            I => uart_pc_data_2
        );

    \I__6848\ : Odrv12
    port map (
            O => \N__30759\,
            I => uart_pc_data_2
        );

    \I__6847\ : CascadeMux
    port map (
            O => \N__30752\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30746\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30742\
        );

    \I__6844\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30739\
        );

    \I__6843\ : Span4Mux_v
    port map (
            O => \N__30742\,
            I => \N__30731\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__30739\,
            I => \N__30731\
        );

    \I__6841\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30725\
        );

    \I__6840\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30721\
        );

    \I__6839\ : InMux
    port map (
            O => \N__30736\,
            I => \N__30718\
        );

    \I__6838\ : Span4Mux_v
    port map (
            O => \N__30731\,
            I => \N__30712\
        );

    \I__6837\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30706\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30706\
        );

    \I__6835\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30703\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__30725\,
            I => \N__30700\
        );

    \I__6833\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30697\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30692\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30692\
        );

    \I__6830\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30689\
        );

    \I__6829\ : InMux
    port map (
            O => \N__30716\,
            I => \N__30686\
        );

    \I__6828\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30683\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__30712\,
            I => \N__30679\
        );

    \I__6826\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30676\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__30706\,
            I => \N__30673\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30703\,
            I => \N__30670\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__30700\,
            I => \N__30667\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__30697\,
            I => \N__30664\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__30692\,
            I => \N__30655\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__30689\,
            I => \N__30655\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30686\,
            I => \N__30655\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__30683\,
            I => \N__30655\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30682\,
            I => \N__30652\
        );

    \I__6816\ : Span4Mux_h
    port map (
            O => \N__30679\,
            I => \N__30649\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30642\
        );

    \I__6814\ : Span4Mux_h
    port map (
            O => \N__30673\,
            I => \N__30642\
        );

    \I__6813\ : Span4Mux_h
    port map (
            O => \N__30670\,
            I => \N__30642\
        );

    \I__6812\ : Odrv4
    port map (
            O => \N__30667\,
            I => uart_pc_data_5
        );

    \I__6811\ : Odrv12
    port map (
            O => \N__30664\,
            I => uart_pc_data_5
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__30655\,
            I => uart_pc_data_5
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__30652\,
            I => uart_pc_data_5
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__30649\,
            I => uart_pc_data_5
        );

    \I__6807\ : Odrv4
    port map (
            O => \N__30642\,
            I => uart_pc_data_5
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__30629\,
            I => \Commands_frame_decoder.state_ns_0_a3_3_1_cascade_\
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__30626\,
            I => \N__30622\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30619\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30615\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30619\,
            I => \N__30612\
        );

    \I__6801\ : CascadeMux
    port map (
            O => \N__30618\,
            I => \N__30609\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__30615\,
            I => \N__30602\
        );

    \I__6799\ : Span4Mux_h
    port map (
            O => \N__30612\,
            I => \N__30602\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30599\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30594\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30607\,
            I => \N__30594\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__30602\,
            I => \N__30591\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__30599\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__30594\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__30591\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__30584\,
            I => \N__30580\
        );

    \I__6790\ : CascadeMux
    port map (
            O => \N__30583\,
            I => \N__30576\
        );

    \I__6789\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30572\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__30579\,
            I => \N__30564\
        );

    \I__6787\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30559\
        );

    \I__6786\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30559\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30554\
        );

    \I__6784\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30551\
        );

    \I__6783\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30546\
        );

    \I__6782\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30546\
        );

    \I__6781\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30540\
        );

    \I__6780\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30540\
        );

    \I__6779\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30537\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30534\
        );

    \I__6777\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30526\
        );

    \I__6776\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30526\
        );

    \I__6775\ : Span4Mux_s2_v
    port map (
            O => \N__30554\,
            I => \N__30523\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__30551\,
            I => \N__30520\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__30546\,
            I => \N__30517\
        );

    \I__6772\ : InMux
    port map (
            O => \N__30545\,
            I => \N__30514\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30511\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__30537\,
            I => \N__30506\
        );

    \I__6769\ : Span4Mux_s2_h
    port map (
            O => \N__30534\,
            I => \N__30506\
        );

    \I__6768\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30501\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30501\
        );

    \I__6766\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30498\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30495\
        );

    \I__6764\ : Sp12to4
    port map (
            O => \N__30523\,
            I => \N__30490\
        );

    \I__6763\ : Span12Mux_v
    port map (
            O => \N__30520\,
            I => \N__30490\
        );

    \I__6762\ : Span4Mux_h
    port map (
            O => \N__30517\,
            I => \N__30487\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30514\,
            I => \N__30482\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__30511\,
            I => \N__30482\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__30506\,
            I => \N__30479\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__30501\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__30498\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6756\ : Odrv12
    port map (
            O => \N__30495\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6755\ : Odrv12
    port map (
            O => \N__30490\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__30487\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6753\ : Odrv4
    port map (
            O => \N__30482\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__30479\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_7\
        );

    \I__6751\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30461\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30461\,
            I => \N__30458\
        );

    \I__6749\ : Span4Mux_h
    port map (
            O => \N__30458\,
            I => \N__30455\
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__30455\,
            I => \ppm_encoder_1.N_320\
        );

    \I__6747\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30449\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__30449\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30443\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30440\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__30440\,
            I => \ppm_encoder_1.pulses2countZ0Z_14\
        );

    \I__6742\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30434\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30434\,
            I => \N__30430\
        );

    \I__6740\ : InMux
    port map (
            O => \N__30433\,
            I => \N__30426\
        );

    \I__6739\ : Span4Mux_h
    port map (
            O => \N__30430\,
            I => \N__30423\
        );

    \I__6738\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30420\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__30426\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__30423\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__30420\,
            I => \ppm_encoder_1.counterZ0Z_14\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__30413\,
            I => \N__30410\
        );

    \I__6733\ : InMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30404\
        );

    \I__6731\ : Odrv12
    port map (
            O => \N__30404\,
            I => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__30398\,
            I => \N__30395\
        );

    \I__6728\ : Span4Mux_h
    port map (
            O => \N__30395\,
            I => \N__30391\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30387\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__30391\,
            I => \N__30384\
        );

    \I__6725\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30381\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30378\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__30384\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__30381\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__30378\,
            I => \ppm_encoder_1.init_pulsesZ0Z_16\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30364\
        );

    \I__6718\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30361\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__30364\,
            I => \N__30358\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30361\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__30358\,
            I => \ppm_encoder_1.pulses2countZ0Z_16\
        );

    \I__6714\ : InMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__30344\,
            I => \N__30339\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30343\,
            I => \N__30334\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30342\,
            I => \N__30334\
        );

    \I__6708\ : Odrv4
    port map (
            O => \N__30339\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__30334\,
            I => \ppm_encoder_1.init_pulsesZ0Z_17\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__30329\,
            I => \N__30326\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30326\,
            I => \N__30323\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__30323\,
            I => \N__30319\
        );

    \I__6703\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__6702\ : Span4Mux_s3_v
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__30316\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__30313\,
            I => \ppm_encoder_1.pulses2countZ0Z_17\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30301\
        );

    \I__6697\ : InMux
    port map (
            O => \N__30304\,
            I => \N__30298\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__30301\,
            I => \N__30295\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__30298\,
            I => \N__30291\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__30295\,
            I => \N__30288\
        );

    \I__6693\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30285\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__30291\,
            I => \N__30282\
        );

    \I__6691\ : Odrv4
    port map (
            O => \N__30288\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__30285\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__30282\,
            I => \ppm_encoder_1.init_pulsesZ0Z_18\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__6687\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30266\
        );

    \I__6686\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30266\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__30266\,
            I => \ppm_encoder_1.pulses2countZ0Z_18\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30260\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30257\
        );

    \I__6682\ : Span4Mux_h
    port map (
            O => \N__30257\,
            I => \N__30254\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__30254\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\
        );

    \I__6680\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30246\
        );

    \I__6679\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30241\
        );

    \I__6678\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30241\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__30246\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__30241\,
            I => \ppm_encoder_1.counterZ0Z_15\
        );

    \I__6675\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30231\
        );

    \I__6674\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30228\
        );

    \I__6673\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30225\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__30231\,
            I => \N__30222\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__30228\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30225\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__30222\,
            I => \ppm_encoder_1.counterZ0Z_17\
        );

    \I__6668\ : CascadeMux
    port map (
            O => \N__30215\,
            I => \N__30210\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30207\
        );

    \I__6666\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30204\
        );

    \I__6665\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30201\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__30207\,
            I => \N__30198\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__30204\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__30201\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__30198\,
            I => \ppm_encoder_1.counterZ0Z_16\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30186\
        );

    \I__6659\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30181\
        );

    \I__6658\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30181\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__30186\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__30181\,
            I => \ppm_encoder_1.counterZ0Z_18\
        );

    \I__6655\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30170\
        );

    \I__6654\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30170\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__30170\,
            I => \N__30167\
        );

    \I__6652\ : Span4Mux_v
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__6651\ : Odrv4
    port map (
            O => \N__30164\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30158\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__30158\,
            I => \N__30155\
        );

    \I__6648\ : Span12Mux_h
    port map (
            O => \N__30155\,
            I => \N__30150\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30145\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30145\
        );

    \I__6645\ : Odrv12
    port map (
            O => \N__30150\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__30145\,
            I => \ppm_encoder_1.init_pulsesZ0Z_15\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__30139\,
            I => \N__30131\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__30138\,
            I => \N__30128\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30121\
        );

    \I__6639\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30121\
        );

    \I__6638\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30121\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30118\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30113\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30113\
        );

    \I__6634\ : Span12Mux_v
    port map (
            O => \N__30113\,
            I => \N__30109\
        );

    \I__6633\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30106\
        );

    \I__6632\ : Odrv12
    port map (
            O => \N__30109\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__30106\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__30101\,
            I => \N__30093\
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__30100\,
            I => \N__30080\
        );

    \I__6628\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30077\
        );

    \I__6627\ : CascadeMux
    port map (
            O => \N__30098\,
            I => \N__30073\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__30097\,
            I => \N__30069\
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__30096\,
            I => \N__30066\
        );

    \I__6624\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30056\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30092\,
            I => \N__30056\
        );

    \I__6622\ : InMux
    port map (
            O => \N__30091\,
            I => \N__30056\
        );

    \I__6621\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30056\
        );

    \I__6620\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \N__30053\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__30088\,
            I => \N__30032\
        );

    \I__6618\ : CascadeMux
    port map (
            O => \N__30087\,
            I => \N__30029\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30017\
        );

    \I__6616\ : InMux
    port map (
            O => \N__30085\,
            I => \N__30017\
        );

    \I__6615\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30017\
        );

    \I__6614\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30014\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30011\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30008\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30005\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30073\,
            I => \N__29994\
        );

    \I__6609\ : InMux
    port map (
            O => \N__30072\,
            I => \N__29994\
        );

    \I__6608\ : InMux
    port map (
            O => \N__30069\,
            I => \N__29994\
        );

    \I__6607\ : InMux
    port map (
            O => \N__30066\,
            I => \N__29994\
        );

    \I__6606\ : InMux
    port map (
            O => \N__30065\,
            I => \N__29994\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__30056\,
            I => \N__29991\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30053\,
            I => \N__29982\
        );

    \I__6603\ : InMux
    port map (
            O => \N__30052\,
            I => \N__29982\
        );

    \I__6602\ : InMux
    port map (
            O => \N__30051\,
            I => \N__29982\
        );

    \I__6601\ : InMux
    port map (
            O => \N__30050\,
            I => \N__29982\
        );

    \I__6600\ : InMux
    port map (
            O => \N__30049\,
            I => \N__29973\
        );

    \I__6599\ : InMux
    port map (
            O => \N__30048\,
            I => \N__29973\
        );

    \I__6598\ : InMux
    port map (
            O => \N__30047\,
            I => \N__29973\
        );

    \I__6597\ : InMux
    port map (
            O => \N__30046\,
            I => \N__29973\
        );

    \I__6596\ : InMux
    port map (
            O => \N__30045\,
            I => \N__29968\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30044\,
            I => \N__29968\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30043\,
            I => \N__29959\
        );

    \I__6593\ : InMux
    port map (
            O => \N__30042\,
            I => \N__29952\
        );

    \I__6592\ : InMux
    port map (
            O => \N__30041\,
            I => \N__29952\
        );

    \I__6591\ : InMux
    port map (
            O => \N__30040\,
            I => \N__29952\
        );

    \I__6590\ : InMux
    port map (
            O => \N__30039\,
            I => \N__29945\
        );

    \I__6589\ : InMux
    port map (
            O => \N__30038\,
            I => \N__29945\
        );

    \I__6588\ : InMux
    port map (
            O => \N__30037\,
            I => \N__29945\
        );

    \I__6587\ : InMux
    port map (
            O => \N__30036\,
            I => \N__29940\
        );

    \I__6586\ : InMux
    port map (
            O => \N__30035\,
            I => \N__29940\
        );

    \I__6585\ : InMux
    port map (
            O => \N__30032\,
            I => \N__29929\
        );

    \I__6584\ : InMux
    port map (
            O => \N__30029\,
            I => \N__29929\
        );

    \I__6583\ : InMux
    port map (
            O => \N__30028\,
            I => \N__29929\
        );

    \I__6582\ : InMux
    port map (
            O => \N__30027\,
            I => \N__29929\
        );

    \I__6581\ : InMux
    port map (
            O => \N__30026\,
            I => \N__29929\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__30025\,
            I => \N__29924\
        );

    \I__6579\ : InMux
    port map (
            O => \N__30024\,
            I => \N__29921\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__30017\,
            I => \N__29918\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__30014\,
            I => \N__29915\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__30011\,
            I => \N__29905\
        );

    \I__6575\ : Span4Mux_v
    port map (
            O => \N__30008\,
            I => \N__29902\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__30005\,
            I => \N__29889\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29889\
        );

    \I__6572\ : Span4Mux_s2_h
    port map (
            O => \N__29991\,
            I => \N__29889\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__29982\,
            I => \N__29889\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__29973\,
            I => \N__29889\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29889\
        );

    \I__6568\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29866\
        );

    \I__6567\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29866\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29866\
        );

    \I__6565\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29866\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29866\
        );

    \I__6563\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29866\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29855\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29855\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__29945\,
            I => \N__29855\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29855\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__29929\,
            I => \N__29855\
        );

    \I__6557\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29848\
        );

    \I__6556\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29848\
        );

    \I__6555\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29848\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__29921\,
            I => \N__29845\
        );

    \I__6553\ : Span4Mux_h
    port map (
            O => \N__29918\,
            I => \N__29842\
        );

    \I__6552\ : Span4Mux_h
    port map (
            O => \N__29915\,
            I => \N__29839\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29832\
        );

    \I__6550\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29832\
        );

    \I__6549\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29832\
        );

    \I__6548\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29823\
        );

    \I__6547\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29823\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29823\
        );

    \I__6545\ : InMux
    port map (
            O => \N__29908\,
            I => \N__29823\
        );

    \I__6544\ : Span4Mux_v
    port map (
            O => \N__29905\,
            I => \N__29816\
        );

    \I__6543\ : Span4Mux_v
    port map (
            O => \N__29902\,
            I => \N__29816\
        );

    \I__6542\ : Span4Mux_v
    port map (
            O => \N__29889\,
            I => \N__29816\
        );

    \I__6541\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29803\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29803\
        );

    \I__6539\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29803\
        );

    \I__6538\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29803\
        );

    \I__6537\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29803\
        );

    \I__6536\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29803\
        );

    \I__6535\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29794\
        );

    \I__6534\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29794\
        );

    \I__6533\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29794\
        );

    \I__6532\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29794\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29785\
        );

    \I__6530\ : Span4Mux_s3_v
    port map (
            O => \N__29855\,
            I => \N__29785\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__29848\,
            I => \N__29785\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__29845\,
            I => \N__29785\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__29842\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__29839\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__29832\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__29823\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__29816\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__29803\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__29794\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__29785\,
            I => \ppm_encoder_1.PPM_STATE_59_d\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__29768\,
            I => \N__29764\
        );

    \I__6518\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__6517\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29758\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__29761\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__29758\,
            I => \ppm_encoder_1.pulses2countZ0Z_15\
        );

    \I__6514\ : CascadeMux
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29744\
        );

    \I__6512\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29744\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__29741\,
            I => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\
        );

    \I__6509\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29734\
        );

    \I__6508\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29731\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__29734\,
            I => \N__29726\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29726\
        );

    \I__6505\ : Odrv12
    port map (
            O => \N__29726\,
            I => scaler_3_data_11
        );

    \I__6504\ : InMux
    port map (
            O => \N__29723\,
            I => \scaler_3.un2_source_data_0_cry_6\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__6502\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29711\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29716\,
            I => \N__29711\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__6499\ : Odrv12
    port map (
            O => \N__29708\,
            I => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\
        );

    \I__6498\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29701\
        );

    \I__6497\ : InMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29692\
        );

    \I__6494\ : Odrv12
    port map (
            O => \N__29695\,
            I => scaler_3_data_12
        );

    \I__6493\ : Odrv12
    port map (
            O => \N__29692\,
            I => scaler_3_data_12
        );

    \I__6492\ : InMux
    port map (
            O => \N__29687\,
            I => \scaler_3.un2_source_data_0_cry_7\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29677\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29674\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__29677\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__29674\,
            I => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\
        );

    \I__6486\ : CascadeMux
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__6485\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29663\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__29660\,
            I => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29653\
        );

    \I__6481\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29650\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__29653\,
            I => \N__29647\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__29650\,
            I => \N__29644\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__6477\ : Span4Mux_v
    port map (
            O => \N__29644\,
            I => \N__29638\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__29641\,
            I => scaler_3_data_13
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__29638\,
            I => scaler_3_data_13
        );

    \I__6474\ : InMux
    port map (
            O => \N__29633\,
            I => \bfn_8_23_0_\
        );

    \I__6473\ : InMux
    port map (
            O => \N__29630\,
            I => \scaler_3.un2_source_data_0_cry_9\
        );

    \I__6472\ : InMux
    port map (
            O => \N__29627\,
            I => \N__29624\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__6470\ : Odrv12
    port map (
            O => \N__29621\,
            I => scaler_3_data_14
        );

    \I__6469\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29614\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__29617\,
            I => \N__29611\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__29614\,
            I => \N__29606\
        );

    \I__6466\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29601\
        );

    \I__6465\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29601\
        );

    \I__6464\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29598\
        );

    \I__6463\ : Span4Mux_v
    port map (
            O => \N__29606\,
            I => \N__29593\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__29601\,
            I => \N__29593\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__29598\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__29593\,
            I => \scaler_3.un2_source_data_0\
        );

    \I__6459\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__6457\ : Span4Mux_v
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__6456\ : Span4Mux_h
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__29576\,
            I => scaler_3_data_5
        );

    \I__6454\ : CEMux
    port map (
            O => \N__29573\,
            I => \N__29552\
        );

    \I__6453\ : CEMux
    port map (
            O => \N__29572\,
            I => \N__29552\
        );

    \I__6452\ : CEMux
    port map (
            O => \N__29571\,
            I => \N__29552\
        );

    \I__6451\ : CEMux
    port map (
            O => \N__29570\,
            I => \N__29552\
        );

    \I__6450\ : CEMux
    port map (
            O => \N__29569\,
            I => \N__29552\
        );

    \I__6449\ : CEMux
    port map (
            O => \N__29568\,
            I => \N__29552\
        );

    \I__6448\ : CEMux
    port map (
            O => \N__29567\,
            I => \N__29552\
        );

    \I__6447\ : GlobalMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__6446\ : gio2CtrlBuf
    port map (
            O => \N__29549\,
            I => \debug_CH3_20A_c_0_g\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__6443\ : Span4Mux_v
    port map (
            O => \N__29540\,
            I => \N__29537\
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__29537\,
            I => \ppm_encoder_1.N_305\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__29534\,
            I => \N__29530\
        );

    \I__6440\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29527\
        );

    \I__6439\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29524\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__29527\,
            I => \N__29520\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29517\
        );

    \I__6436\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29514\
        );

    \I__6435\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29509\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__29517\,
            I => \N__29509\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29514\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__6432\ : Odrv4
    port map (
            O => \N__29509\,
            I => \ppm_encoder_1.aileronZ0Z_13\
        );

    \I__6431\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29501\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__29501\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\
        );

    \I__6429\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29495\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29491\
        );

    \I__6427\ : InMux
    port map (
            O => \N__29494\,
            I => \N__29486\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__29491\,
            I => \N__29477\
        );

    \I__6425\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29474\
        );

    \I__6424\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29471\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__29486\,
            I => \N__29468\
        );

    \I__6422\ : InMux
    port map (
            O => \N__29485\,
            I => \N__29463\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__29484\,
            I => \N__29457\
        );

    \I__6420\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29454\
        );

    \I__6419\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29449\
        );

    \I__6418\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29449\
        );

    \I__6417\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29446\
        );

    \I__6416\ : Span4Mux_h
    port map (
            O => \N__29477\,
            I => \N__29441\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__29474\,
            I => \N__29441\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29436\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__29468\,
            I => \N__29436\
        );

    \I__6412\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29431\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29431\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__29463\,
            I => \N__29428\
        );

    \I__6409\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29423\
        );

    \I__6408\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29420\
        );

    \I__6407\ : InMux
    port map (
            O => \N__29460\,
            I => \N__29415\
        );

    \I__6406\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29415\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29412\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29409\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__29446\,
            I => \N__29402\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__29441\,
            I => \N__29402\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__29436\,
            I => \N__29402\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__29431\,
            I => \N__29399\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__29428\,
            I => \N__29396\
        );

    \I__6398\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29393\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29426\,
            I => \N__29389\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29385\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29374\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29415\,
            I => \N__29374\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__29412\,
            I => \N__29374\
        );

    \I__6392\ : Span4Mux_v
    port map (
            O => \N__29409\,
            I => \N__29374\
        );

    \I__6391\ : Span4Mux_v
    port map (
            O => \N__29402\,
            I => \N__29374\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__29399\,
            I => \N__29367\
        );

    \I__6389\ : Span4Mux_v
    port map (
            O => \N__29396\,
            I => \N__29367\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29367\
        );

    \I__6387\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29364\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__29389\,
            I => \N__29361\
        );

    \I__6385\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29358\
        );

    \I__6384\ : Span12Mux_v
    port map (
            O => \N__29385\,
            I => \N__29355\
        );

    \I__6383\ : Span4Mux_v
    port map (
            O => \N__29374\,
            I => \N__29352\
        );

    \I__6382\ : Span4Mux_v
    port map (
            O => \N__29367\,
            I => \N__29349\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__29364\,
            I => \N__29344\
        );

    \I__6380\ : Span12Mux_v
    port map (
            O => \N__29361\,
            I => \N__29344\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__29358\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6378\ : Odrv12
    port map (
            O => \N__29355\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__29352\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__29349\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6375\ : Odrv12
    port map (
            O => \N__29344\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\
        );

    \I__6374\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__29330\,
            I => \N__29326\
        );

    \I__6372\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29322\
        );

    \I__6371\ : Span4Mux_h
    port map (
            O => \N__29326\,
            I => \N__29319\
        );

    \I__6370\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29316\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29313\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__29319\,
            I => \N__29308\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29308\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__29313\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__6365\ : Odrv4
    port map (
            O => \N__29308\,
            I => \ppm_encoder_1.throttleZ0Z_6\
        );

    \I__6364\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29298\
        );

    \I__6363\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29295\
        );

    \I__6362\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29292\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29289\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__29295\,
            I => \N__29286\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__29292\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__6358\ : Odrv4
    port map (
            O => \N__29289\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__29286\,
            I => \ppm_encoder_1.elevatorZ0Z_6\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__29279\,
            I => \N__29276\
        );

    \I__6355\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29269\
        );

    \I__6354\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29263\
        );

    \I__6353\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29263\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29254\
        );

    \I__6351\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29254\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29269\,
            I => \N__29249\
        );

    \I__6349\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29246\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29241\
        );

    \I__6347\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29238\
        );

    \I__6346\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29230\
        );

    \I__6345\ : InMux
    port map (
            O => \N__29260\,
            I => \N__29230\
        );

    \I__6344\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29230\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29227\
        );

    \I__6342\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29224\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__29252\,
            I => \N__29219\
        );

    \I__6340\ : Span4Mux_s2_v
    port map (
            O => \N__29249\,
            I => \N__29214\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29211\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29206\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29206\
        );

    \I__6336\ : Span4Mux_v
    port map (
            O => \N__29241\,
            I => \N__29203\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__29238\,
            I => \N__29200\
        );

    \I__6334\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29197\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29230\,
            I => \N__29188\
        );

    \I__6332\ : Span4Mux_s2_v
    port map (
            O => \N__29227\,
            I => \N__29188\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__29224\,
            I => \N__29188\
        );

    \I__6330\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29185\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__29222\,
            I => \N__29182\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29174\
        );

    \I__6327\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29174\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29174\
        );

    \I__6325\ : Span4Mux_v
    port map (
            O => \N__29214\,
            I => \N__29169\
        );

    \I__6324\ : Span4Mux_v
    port map (
            O => \N__29211\,
            I => \N__29169\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__29206\,
            I => \N__29166\
        );

    \I__6322\ : Span4Mux_v
    port map (
            O => \N__29203\,
            I => \N__29161\
        );

    \I__6321\ : Span4Mux_h
    port map (
            O => \N__29200\,
            I => \N__29161\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__29197\,
            I => \N__29158\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29196\,
            I => \N__29153\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29153\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__29188\,
            I => \N__29148\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29148\
        );

    \I__6315\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29143\
        );

    \I__6314\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29143\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__29174\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6312\ : Odrv4
    port map (
            O => \N__29169\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6311\ : Odrv12
    port map (
            O => \N__29166\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__29161\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__29158\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__29153\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__29148\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29143\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__29126\,
            I => \ppm_encoder_1.N_298_cascade_\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \N__29119\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29116\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29113\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29109\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__29113\,
            I => \N__29106\
        );

    \I__6299\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29103\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__29109\,
            I => \N__29098\
        );

    \I__6297\ : Span4Mux_s3_h
    port map (
            O => \N__29106\,
            I => \N__29098\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__29103\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__6295\ : Odrv4
    port map (
            O => \N__29098\,
            I => \ppm_encoder_1.aileronZ0Z_6\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__29090\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29083\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29086\,
            I => \N__29080\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29074\
        );

    \I__6288\ : Span4Mux_h
    port map (
            O => \N__29077\,
            I => \N__29071\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__29074\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__29071\,
            I => \frame_decoder_OFF3data_7\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29063\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29059\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29056\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__29059\,
            I => \N__29053\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__29050\,
            I => \frame_decoder_CH3data_7\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__29047\,
            I => \frame_decoder_CH3data_7\
        );

    \I__6277\ : InMux
    port map (
            O => \N__29042\,
            I => \N__29039\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__29039\,
            I => \scaler_3.N_893_i_l_ofxZ0\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29030\,
            I => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\
        );

    \I__6272\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__29024\,
            I => \N__29020\
        );

    \I__6270\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29017\
        );

    \I__6269\ : Span4Mux_h
    port map (
            O => \N__29020\,
            I => \N__29014\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__29011\
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__29014\,
            I => scaler_3_data_6
        );

    \I__6266\ : Odrv12
    port map (
            O => \N__29011\,
            I => scaler_3_data_6
        );

    \I__6265\ : InMux
    port map (
            O => \N__29006\,
            I => \scaler_3.un2_source_data_0_cry_1\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__6263\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28994\
        );

    \I__6262\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28994\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__28991\,
            I => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__6258\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28979\
        );

    \I__6256\ : Span4Mux_h
    port map (
            O => \N__28979\,
            I => \N__28975\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28972\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__28975\,
            I => \N__28969\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28966\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__28969\,
            I => scaler_3_data_7
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__28966\,
            I => scaler_3_data_7
        );

    \I__6250\ : InMux
    port map (
            O => \N__28961\,
            I => \scaler_3.un2_source_data_0_cry_2\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__28958\,
            I => \N__28955\
        );

    \I__6248\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28949\
        );

    \I__6247\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28949\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__28949\,
            I => \N__28946\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__28946\,
            I => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\
        );

    \I__6244\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28940\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__28940\,
            I => \N__28936\
        );

    \I__6242\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28933\
        );

    \I__6241\ : Span4Mux_v
    port map (
            O => \N__28936\,
            I => \N__28928\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28928\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__28928\,
            I => scaler_3_data_8
        );

    \I__6238\ : InMux
    port map (
            O => \N__28925\,
            I => \scaler_3.un2_source_data_0_cry_3\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__28922\,
            I => \N__28919\
        );

    \I__6236\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28913\
        );

    \I__6235\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28913\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__28910\,
            I => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\
        );

    \I__6232\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28904\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28900\
        );

    \I__6230\ : InMux
    port map (
            O => \N__28903\,
            I => \N__28897\
        );

    \I__6229\ : Span12Mux_s8_h
    port map (
            O => \N__28900\,
            I => \N__28894\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__28897\,
            I => \N__28891\
        );

    \I__6227\ : Odrv12
    port map (
            O => \N__28894\,
            I => scaler_3_data_9
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__28891\,
            I => scaler_3_data_9
        );

    \I__6225\ : InMux
    port map (
            O => \N__28886\,
            I => \scaler_3.un2_source_data_0_cry_4\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__28883\,
            I => \N__28880\
        );

    \I__6223\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28874\
        );

    \I__6222\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28874\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__6220\ : Odrv12
    port map (
            O => \N__28871\,
            I => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\
        );

    \I__6219\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__28865\,
            I => \N__28861\
        );

    \I__6217\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28858\
        );

    \I__6216\ : Span4Mux_v
    port map (
            O => \N__28861\,
            I => \N__28853\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28853\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__28853\,
            I => scaler_3_data_10
        );

    \I__6213\ : InMux
    port map (
            O => \N__28850\,
            I => \scaler_3.un2_source_data_0_cry_5\
        );

    \I__6212\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__28844\,
            I => \frame_decoder_CH3data_2\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28838\
        );

    \I__6209\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28835\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28832\
        );

    \I__6207\ : Odrv12
    port map (
            O => \N__28832\,
            I => \frame_decoder_OFF3data_2\
        );

    \I__6206\ : InMux
    port map (
            O => \N__28829\,
            I => \scaler_3.un3_source_data_0_cry_1\
        );

    \I__6205\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__6203\ : Odrv4
    port map (
            O => \N__28820\,
            I => \frame_decoder_OFF3data_3\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__6201\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28811\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__28811\,
            I => \frame_decoder_CH3data_3\
        );

    \I__6199\ : InMux
    port map (
            O => \N__28808\,
            I => \scaler_3.un3_source_data_0_cry_2\
        );

    \I__6198\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__28799\,
            I => \N__28796\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__28796\,
            I => \frame_decoder_CH3data_4\
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__28793\,
            I => \N__28790\
        );

    \I__6193\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28787\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__28787\,
            I => \N__28784\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__28784\,
            I => \frame_decoder_OFF3data_4\
        );

    \I__6190\ : InMux
    port map (
            O => \N__28781\,
            I => \scaler_3.un3_source_data_0_cry_3\
        );

    \I__6189\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28775\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__28775\,
            I => \frame_decoder_CH3data_5\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__28772\,
            I => \N__28769\
        );

    \I__6186\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__6184\ : Odrv12
    port map (
            O => \N__28763\,
            I => \frame_decoder_OFF3data_5\
        );

    \I__6183\ : InMux
    port map (
            O => \N__28760\,
            I => \scaler_3.un3_source_data_0_cry_4\
        );

    \I__6182\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28754\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__28754\,
            I => \frame_decoder_CH3data_6\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__6179\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28745\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__28745\,
            I => \N__28742\
        );

    \I__6177\ : Odrv4
    port map (
            O => \N__28742\,
            I => \frame_decoder_OFF3data_6\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28739\,
            I => \scaler_3.un3_source_data_0_cry_5\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28733\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28730\
        );

    \I__6173\ : Span4Mux_v
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__28724\,
            I => \scaler_3.un3_source_data_0_axb_7\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28721\,
            I => \scaler_3.un3_source_data_0_cry_6\
        );

    \I__6169\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28714\
        );

    \I__6168\ : InMux
    port map (
            O => \N__28717\,
            I => \N__28711\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__28714\,
            I => \N__28708\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__28711\,
            I => \N__28705\
        );

    \I__6165\ : Span4Mux_h
    port map (
            O => \N__28708\,
            I => \N__28694\
        );

    \I__6164\ : Span4Mux_v
    port map (
            O => \N__28705\,
            I => \N__28694\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28691\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__28703\,
            I => \N__28687\
        );

    \I__6161\ : CascadeMux
    port map (
            O => \N__28702\,
            I => \N__28682\
        );

    \I__6160\ : CascadeMux
    port map (
            O => \N__28701\,
            I => \N__28679\
        );

    \I__6159\ : CascadeMux
    port map (
            O => \N__28700\,
            I => \N__28675\
        );

    \I__6158\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28668\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__28694\,
            I => \N__28663\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__28691\,
            I => \N__28663\
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__28690\,
            I => \N__28660\
        );

    \I__6154\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28654\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28641\
        );

    \I__6152\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28641\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28641\
        );

    \I__6150\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28641\
        );

    \I__6149\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28641\
        );

    \I__6148\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28641\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__28674\,
            I => \N__28638\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__28673\,
            I => \N__28635\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__28672\,
            I => \N__28632\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__28671\,
            I => \N__28629\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28626\
        );

    \I__6142\ : Span4Mux_h
    port map (
            O => \N__28663\,
            I => \N__28623\
        );

    \I__6141\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28620\
        );

    \I__6140\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28617\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__28658\,
            I => \N__28614\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \N__28611\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__28654\,
            I => \N__28606\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__28641\,
            I => \N__28606\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28603\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28599\
        );

    \I__6133\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28596\
        );

    \I__6132\ : InMux
    port map (
            O => \N__28629\,
            I => \N__28593\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__28626\,
            I => \N__28584\
        );

    \I__6130\ : Span4Mux_v
    port map (
            O => \N__28623\,
            I => \N__28584\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__28620\,
            I => \N__28584\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28617\,
            I => \N__28584\
        );

    \I__6127\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28581\
        );

    \I__6126\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28578\
        );

    \I__6125\ : Span4Mux_v
    port map (
            O => \N__28606\,
            I => \N__28573\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28573\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__28602\,
            I => \N__28570\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28562\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__28596\,
            I => \N__28562\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28559\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__28584\,
            I => \N__28556\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__28581\,
            I => \N__28553\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28548\
        );

    \I__6116\ : Span4Mux_v
    port map (
            O => \N__28573\,
            I => \N__28548\
        );

    \I__6115\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28545\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__28569\,
            I => \N__28542\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__28568\,
            I => \N__28539\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__28567\,
            I => \N__28536\
        );

    \I__6111\ : Span4Mux_v
    port map (
            O => \N__28562\,
            I => \N__28532\
        );

    \I__6110\ : Span4Mux_v
    port map (
            O => \N__28559\,
            I => \N__28529\
        );

    \I__6109\ : Span4Mux_v
    port map (
            O => \N__28556\,
            I => \N__28526\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__28553\,
            I => \N__28523\
        );

    \I__6107\ : Span4Mux_h
    port map (
            O => \N__28548\,
            I => \N__28518\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28518\
        );

    \I__6105\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28515\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28510\
        );

    \I__6103\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28510\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__28535\,
            I => \N__28507\
        );

    \I__6101\ : Span4Mux_h
    port map (
            O => \N__28532\,
            I => \N__28504\
        );

    \I__6100\ : Span4Mux_h
    port map (
            O => \N__28529\,
            I => \N__28497\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__28526\,
            I => \N__28497\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__28523\,
            I => \N__28497\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__28518\,
            I => \N__28490\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__28515\,
            I => \N__28490\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__28510\,
            I => \N__28490\
        );

    \I__6094\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28487\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__28504\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__28497\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__28490\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28487\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6089\ : InMux
    port map (
            O => \N__28478\,
            I => \bfn_8_21_0_\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28475\,
            I => \scaler_3.un3_source_data_0_cry_8\
        );

    \I__6087\ : CEMux
    port map (
            O => \N__28472\,
            I => \N__28469\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28465\
        );

    \I__6085\ : CEMux
    port map (
            O => \N__28468\,
            I => \N__28461\
        );

    \I__6084\ : Span4Mux_h
    port map (
            O => \N__28465\,
            I => \N__28458\
        );

    \I__6083\ : CEMux
    port map (
            O => \N__28464\,
            I => \N__28455\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28461\,
            I => \N__28452\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__28458\,
            I => \N__28447\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__28455\,
            I => \N__28447\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__28452\,
            I => \N__28444\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__28447\,
            I => \N__28441\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__28444\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__28441\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\
        );

    \I__6075\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__28433\,
            I => \frame_decoder_CH3data_1\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28424\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28421\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__28421\,
            I => \frame_decoder_OFF3data_1\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28418\,
            I => \scaler_3.un3_source_data_0_cry_0\
        );

    \I__6068\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28411\
        );

    \I__6067\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28408\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__28411\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__28408\,
            I => \uart_drone.data_AuxZ0Z_3\
        );

    \I__6064\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28399\
        );

    \I__6063\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28396\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__28399\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__28396\,
            I => \uart_drone.data_AuxZ0Z_5\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__28391\,
            I => \N__28387\
        );

    \I__6059\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28384\
        );

    \I__6058\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28381\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__28384\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__28381\,
            I => \uart_drone.data_AuxZ0Z_6\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__28376\,
            I => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\
        );

    \I__6054\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28369\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28366\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28369\,
            I => \N__28363\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__28366\,
            I => \N__28360\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__28363\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__28360\,
            I => \frame_decoder_OFF4data_7\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28351\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__28348\,
            I => \N__28342\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__28345\,
            I => \N__28339\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__28342\,
            I => \frame_decoder_CH4data_7\
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__28339\,
            I => \frame_decoder_CH4data_7\
        );

    \I__6041\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28328\
        );

    \I__6039\ : Span4Mux_v
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__28325\,
            I => \scaler_4.un3_source_data_0_axb_7\
        );

    \I__6037\ : CascadeMux
    port map (
            O => \N__28322\,
            I => \N__28318\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28321\,
            I => \N__28315\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28312\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__28315\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__28312\,
            I => \uart_drone.data_AuxZ0Z_0\
        );

    \I__6032\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28303\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28300\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__28303\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28300\,
            I => \uart_drone.data_AuxZ0Z_1\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__6027\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28288\
        );

    \I__6026\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28285\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28282\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__28285\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__28282\,
            I => \uart_drone.data_AuxZ0Z_2\
        );

    \I__6022\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28271\
        );

    \I__6021\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28271\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__28271\,
            I => \Commands_frame_decoder.stateZ0Z_7\
        );

    \I__6019\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__28259\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__28256\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28249\
        );

    \I__6013\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__28249\,
            I => \Commands_frame_decoder.stateZ0Z_8\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__28246\,
            I => \Commands_frame_decoder.stateZ0Z_8\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28231\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28231\
        );

    \I__6008\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28231\
        );

    \I__6007\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28228\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__28228\,
            I => \N__28220\
        );

    \I__6004\ : Span4Mux_v
    port map (
            O => \N__28225\,
            I => \N__28220\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__28220\,
            I => \dron_frame_decoder_1.stateZ0Z_5\
        );

    \I__6002\ : InMux
    port map (
            O => \N__28217\,
            I => \N__28213\
        );

    \I__6001\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28210\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__28213\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__28210\,
            I => \Commands_frame_decoder.source_CH3data_1_sqmuxa\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28201\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28198\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__28201\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__28198\,
            I => \Commands_frame_decoder.stateZ0Z_5\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__28190\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__5991\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28181\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__28181\,
            I => \N__28178\
        );

    \I__5989\ : Span4Mux_v
    port map (
            O => \N__28178\,
            I => \N__28173\
        );

    \I__5988\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28170\
        );

    \I__5987\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28166\
        );

    \I__5986\ : Span4Mux_h
    port map (
            O => \N__28173\,
            I => \N__28161\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28161\
        );

    \I__5984\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28158\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__28166\,
            I => \N__28153\
        );

    \I__5982\ : Sp12to4
    port map (
            O => \N__28161\,
            I => \N__28153\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__28158\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__5980\ : Odrv12
    port map (
            O => \N__28153\,
            I => \Commands_frame_decoder.stateZ0Z_6\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28144\
        );

    \I__5978\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28141\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__28144\,
            I => \N__28138\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__28141\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__5975\ : Odrv12
    port map (
            O => \N__28138\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa\
        );

    \I__5974\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28129\
        );

    \I__5973\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__28129\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__28126\,
            I => \Commands_frame_decoder.stateZ0Z_4\
        );

    \I__5970\ : CEMux
    port map (
            O => \N__28121\,
            I => \N__28118\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28115\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__28115\,
            I => \N__28112\
        );

    \I__5967\ : Span4Mux_h
    port map (
            O => \N__28112\,
            I => \N__28108\
        );

    \I__5966\ : CEMux
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__28108\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__28105\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__28100\,
            I => \N__28096\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__28099\,
            I => \N__28093\
        );

    \I__5961\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28087\
        );

    \I__5960\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28087\
        );

    \I__5959\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28084\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__28087\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__28084\,
            I => \dron_frame_decoder_1.stateZ0Z_4\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28073\
        );

    \I__5955\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28073\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__28073\,
            I => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\
        );

    \I__5953\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__28067\,
            I => \N__28063\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28060\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__28063\,
            I => \N__28057\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28054\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__28057\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1_0\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__28054\,
            I => \Commands_frame_decoder.state_ns_i_a2_1_1_0\
        );

    \I__5946\ : CEMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28042\
        );

    \I__5944\ : CEMux
    port map (
            O => \N__28045\,
            I => \N__28038\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__28042\,
            I => \N__28035\
        );

    \I__5942\ : CEMux
    port map (
            O => \N__28041\,
            I => \N__28032\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__28038\,
            I => \N__28029\
        );

    \I__5940\ : Span4Mux_h
    port map (
            O => \N__28035\,
            I => \N__28024\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28024\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__28029\,
            I => \N__28021\
        );

    \I__5937\ : Span4Mux_v
    port map (
            O => \N__28024\,
            I => \N__28018\
        );

    \I__5936\ : Span4Mux_h
    port map (
            O => \N__28021\,
            I => \N__28015\
        );

    \I__5935\ : Span4Mux_v
    port map (
            O => \N__28018\,
            I => \N__28012\
        );

    \I__5934\ : Span4Mux_h
    port map (
            O => \N__28015\,
            I => \N__28009\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__28012\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__28009\,
            I => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\
        );

    \I__5931\ : InMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__28001\,
            I => \N__27997\
        );

    \I__5929\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27994\
        );

    \I__5928\ : Odrv4
    port map (
            O => \N__27997\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__27994\,
            I => \Commands_frame_decoder.source_offset4data_1_sqmuxa\
        );

    \I__5926\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27980\
        );

    \I__5925\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27980\
        );

    \I__5924\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27980\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__27980\,
            I => \Commands_frame_decoder.stateZ0Z_10\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27977\,
            I => \ppm_encoder_1.un1_counter_13_cry_17\
        );

    \I__5921\ : SRMux
    port map (
            O => \N__27974\,
            I => \N__27965\
        );

    \I__5920\ : SRMux
    port map (
            O => \N__27973\,
            I => \N__27965\
        );

    \I__5919\ : SRMux
    port map (
            O => \N__27972\,
            I => \N__27965\
        );

    \I__5918\ : GlobalMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__5917\ : gio2CtrlBuf
    port map (
            O => \N__27962\,
            I => \ppm_encoder_1.N_320_g\
        );

    \I__5916\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27950\
        );

    \I__5915\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27950\
        );

    \I__5914\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27942\
        );

    \I__5913\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27942\
        );

    \I__5912\ : InMux
    port map (
            O => \N__27955\,
            I => \N__27938\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27935\
        );

    \I__5910\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27930\
        );

    \I__5909\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27930\
        );

    \I__5908\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27927\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27919\
        );

    \I__5906\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27916\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__27938\,
            I => \N__27907\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__27935\,
            I => \N__27907\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__27930\,
            I => \N__27907\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__27927\,
            I => \N__27907\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27902\
        );

    \I__5900\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27902\
        );

    \I__5899\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27899\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__27923\,
            I => \N__27891\
        );

    \I__5897\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27888\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__27919\,
            I => \N__27885\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27882\
        );

    \I__5894\ : Span4Mux_v
    port map (
            O => \N__27907\,
            I => \N__27877\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__27902\,
            I => \N__27877\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27874\
        );

    \I__5891\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27867\
        );

    \I__5890\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27867\
        );

    \I__5889\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27867\
        );

    \I__5888\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27862\
        );

    \I__5887\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27862\
        );

    \I__5886\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27859\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__27888\,
            I => \N__27856\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__27885\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__27882\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__27877\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__27874\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__27867\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__27862\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__27859\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5877\ : Odrv4
    port map (
            O => \N__27856\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \N__27834\
        );

    \I__5875\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27831\
        );

    \I__5874\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27828\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27825\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27822\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27819\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27816\
        );

    \I__5869\ : Span4Mux_h
    port map (
            O => \N__27822\,
            I => \N__27813\
        );

    \I__5868\ : Span4Mux_h
    port map (
            O => \N__27819\,
            I => \N__27806\
        );

    \I__5867\ : Span4Mux_s1_v
    port map (
            O => \N__27816\,
            I => \N__27806\
        );

    \I__5866\ : Span4Mux_v
    port map (
            O => \N__27813\,
            I => \N__27806\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__27806\,
            I => \ppm_encoder_1.init_pulsesZ0Z_12\
        );

    \I__5864\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27796\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27793\
        );

    \I__5861\ : Span4Mux_v
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__5860\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27786\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__27790\,
            I => \N__27783\
        );

    \I__5858\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27780\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__27786\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__27783\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27780\,
            I => \ppm_encoder_1.rudderZ0Z_12\
        );

    \I__5854\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27770\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__27770\,
            I => \uart_pc_sync.aux_2__0_Z0Z_0\
        );

    \I__5852\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__27764\,
            I => \uart_pc_sync.aux_3__0_Z0Z_0\
        );

    \I__5850\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27758\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__5848\ : Odrv12
    port map (
            O => \N__27755\,
            I => uart_input_drone_c
        );

    \I__5847\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27749\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27746\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__27746\,
            I => \uart_drone_sync.aux_0__0__0_0\
        );

    \I__5844\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__27740\,
            I => \uart_drone_sync.aux_1__0__0_0\
        );

    \I__5842\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__27734\,
            I => \uart_drone_sync.aux_2__0__0_0\
        );

    \I__5840\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27727\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27724\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__27727\,
            I => \N__27720\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27717\
        );

    \I__5836\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27714\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__27720\,
            I => \N__27711\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__27717\,
            I => \N__27708\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27714\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__27711\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__27708\,
            I => \ppm_encoder_1.counterZ0Z_9\
        );

    \I__5830\ : InMux
    port map (
            O => \N__27701\,
            I => \ppm_encoder_1.un1_counter_13_cry_8\
        );

    \I__5829\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27695\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27690\
        );

    \I__5827\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27687\
        );

    \I__5826\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27684\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__27690\,
            I => \N__27681\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__27687\,
            I => \N__27678\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__27684\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__27681\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__27678\,
            I => \ppm_encoder_1.counterZ0Z_10\
        );

    \I__5820\ : InMux
    port map (
            O => \N__27671\,
            I => \ppm_encoder_1.un1_counter_13_cry_9\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__27668\,
            I => \N__27665\
        );

    \I__5818\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27657\
        );

    \I__5816\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27654\
        );

    \I__5815\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27651\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__27657\,
            I => \N__27648\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__27654\,
            I => \N__27645\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__27651\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__27648\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__27645\,
            I => \ppm_encoder_1.counterZ0Z_11\
        );

    \I__5809\ : InMux
    port map (
            O => \N__27638\,
            I => \ppm_encoder_1.un1_counter_13_cry_10\
        );

    \I__5808\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27632\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__27632\,
            I => \N__27627\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27624\
        );

    \I__5805\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27621\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__27627\,
            I => \N__27618\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27615\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__27621\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__27618\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5800\ : Odrv12
    port map (
            O => \N__27615\,
            I => \ppm_encoder_1.counterZ0Z_12\
        );

    \I__5799\ : InMux
    port map (
            O => \N__27608\,
            I => \ppm_encoder_1.un1_counter_13_cry_11\
        );

    \I__5798\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__27602\,
            I => \N__27597\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27594\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27591\
        );

    \I__5794\ : Span4Mux_h
    port map (
            O => \N__27597\,
            I => \N__27588\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27585\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__27591\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__27588\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5790\ : Odrv4
    port map (
            O => \N__27585\,
            I => \ppm_encoder_1.counterZ0Z_13\
        );

    \I__5789\ : InMux
    port map (
            O => \N__27578\,
            I => \ppm_encoder_1.un1_counter_13_cry_12\
        );

    \I__5788\ : InMux
    port map (
            O => \N__27575\,
            I => \ppm_encoder_1.un1_counter_13_cry_13\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27572\,
            I => \ppm_encoder_1.un1_counter_13_cry_14\
        );

    \I__5786\ : InMux
    port map (
            O => \N__27569\,
            I => \bfn_7_28_0_\
        );

    \I__5785\ : InMux
    port map (
            O => \N__27566\,
            I => \ppm_encoder_1.un1_counter_13_cry_16\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__27563\,
            I => \N__27559\
        );

    \I__5783\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27554\
        );

    \I__5782\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27549\
        );

    \I__5781\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27549\
        );

    \I__5780\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27546\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__27554\,
            I => \N__27541\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__27549\,
            I => \N__27541\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__27546\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__27541\,
            I => \ppm_encoder_1.counterZ0Z_1\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27536\,
            I => \ppm_encoder_1.un1_counter_13_cry_0\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__27533\,
            I => \N__27528\
        );

    \I__5773\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27520\
        );

    \I__5772\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27520\
        );

    \I__5771\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27520\
        );

    \I__5770\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27517\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__27517\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__27514\,
            I => \ppm_encoder_1.counterZ0Z_2\
        );

    \I__5766\ : InMux
    port map (
            O => \N__27509\,
            I => \ppm_encoder_1.un1_counter_13_cry_1\
        );

    \I__5765\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27496\
        );

    \I__5764\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27496\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27496\
        );

    \I__5762\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27493\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__27496\,
            I => \N__27490\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__27493\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__27490\,
            I => \ppm_encoder_1.counterZ0Z_3\
        );

    \I__5758\ : InMux
    port map (
            O => \N__27485\,
            I => \ppm_encoder_1.un1_counter_13_cry_2\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27478\
        );

    \I__5756\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27474\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__27478\,
            I => \N__27471\
        );

    \I__5754\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27468\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27465\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__27471\,
            I => \N__27462\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27468\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__27465\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__27462\,
            I => \ppm_encoder_1.counterZ0Z_4\
        );

    \I__5748\ : InMux
    port map (
            O => \N__27455\,
            I => \ppm_encoder_1.un1_counter_13_cry_3\
        );

    \I__5747\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27448\
        );

    \I__5746\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27444\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27448\,
            I => \N__27441\
        );

    \I__5744\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27438\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27435\
        );

    \I__5742\ : Span4Mux_v
    port map (
            O => \N__27441\,
            I => \N__27432\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__27438\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__27435\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__27432\,
            I => \ppm_encoder_1.counterZ0Z_5\
        );

    \I__5738\ : InMux
    port map (
            O => \N__27425\,
            I => \ppm_encoder_1.un1_counter_13_cry_4\
        );

    \I__5737\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27418\
        );

    \I__5736\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27414\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27411\
        );

    \I__5734\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27408\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__27414\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__27411\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__27408\,
            I => \ppm_encoder_1.counterZ0Z_6\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27401\,
            I => \ppm_encoder_1.un1_counter_13_cry_5\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__5728\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27391\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27387\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__27391\,
            I => \N__27384\
        );

    \I__5725\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27381\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__27387\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__27384\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__27381\,
            I => \ppm_encoder_1.counterZ0Z_7\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27374\,
            I => \ppm_encoder_1.un1_counter_13_cry_6\
        );

    \I__5720\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27368\,
            I => \N__27364\
        );

    \I__5718\ : InMux
    port map (
            O => \N__27367\,
            I => \N__27361\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__27364\,
            I => \N__27357\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27361\,
            I => \N__27354\
        );

    \I__5715\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27351\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__27357\,
            I => \N__27348\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__27354\,
            I => \N__27345\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__27351\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__27348\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__27345\,
            I => \ppm_encoder_1.counterZ0Z_8\
        );

    \I__5709\ : InMux
    port map (
            O => \N__27338\,
            I => \bfn_7_27_0_\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27332\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__5706\ : Odrv4
    port map (
            O => \N__27329\,
            I => scaler_4_data_5
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__27326\,
            I => \N__27323\
        );

    \I__5704\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27320\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27316\
        );

    \I__5702\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27313\
        );

    \I__5701\ : Span12Mux_s7_h
    port map (
            O => \N__27316\,
            I => \N__27310\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27313\,
            I => \N__27307\
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__27310\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__5698\ : Odrv12
    port map (
            O => \N__27307\,
            I => \ppm_encoder_1.rudderZ0Z_5\
        );

    \I__5697\ : CEMux
    port map (
            O => \N__27302\,
            I => \N__27298\
        );

    \I__5696\ : CEMux
    port map (
            O => \N__27301\,
            I => \N__27295\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27290\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__27295\,
            I => \N__27287\
        );

    \I__5693\ : CEMux
    port map (
            O => \N__27294\,
            I => \N__27284\
        );

    \I__5692\ : CEMux
    port map (
            O => \N__27293\,
            I => \N__27280\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__27290\,
            I => \N__27277\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__27287\,
            I => \N__27274\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__27284\,
            I => \N__27271\
        );

    \I__5688\ : CEMux
    port map (
            O => \N__27283\,
            I => \N__27268\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__27280\,
            I => \N__27264\
        );

    \I__5686\ : Span4Mux_s2_h
    port map (
            O => \N__27277\,
            I => \N__27261\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__27274\,
            I => \N__27256\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__27271\,
            I => \N__27256\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__27268\,
            I => \N__27253\
        );

    \I__5682\ : CEMux
    port map (
            O => \N__27267\,
            I => \N__27250\
        );

    \I__5681\ : Odrv12
    port map (
            O => \N__27264\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__27261\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__27256\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5678\ : Odrv12
    port map (
            O => \N__27253\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__27250\,
            I => \ppm_encoder_1.pid_altitude_dv_0\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__5675\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27233\,
            I => \N__27230\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__27230\,
            I => \N__27227\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__27227\,
            I => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\
        );

    \I__5671\ : InMux
    port map (
            O => \N__27224\,
            I => \N__27221\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__27218\,
            I => \N__27215\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__27215\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\
        );

    \I__5667\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__27209\,
            I => \ppm_encoder_1.pulses2countZ0Z_6\
        );

    \I__5665\ : InMux
    port map (
            O => \N__27206\,
            I => \N__27203\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__27200\,
            I => \N__27197\
        );

    \I__5662\ : Span4Mux_h
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__27194\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27188\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__27188\,
            I => \N__27185\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__27185\,
            I => \N__27182\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__27182\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__27179\,
            I => \N__27176\
        );

    \I__5655\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27173\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__27173\,
            I => \ppm_encoder_1.pulses2countZ0Z_7\
        );

    \I__5653\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27167\,
            I => \N__27164\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__27161\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\
        );

    \I__5649\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__27155\,
            I => \ppm_encoder_1.pulses2countZ0Z_12\
        );

    \I__5647\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27149\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__27143\,
            I => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__27134\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27125\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__27125\,
            I => \ppm_encoder_1.pulses2countZ0Z_13\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__27122\,
            I => \N__27114\
        );

    \I__5636\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27098\
        );

    \I__5635\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27098\
        );

    \I__5634\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27098\
        );

    \I__5633\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27093\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27093\
        );

    \I__5631\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27080\
        );

    \I__5630\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27080\
        );

    \I__5629\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27080\
        );

    \I__5628\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27080\
        );

    \I__5627\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27080\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27080\
        );

    \I__5625\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27071\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27071\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27071\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27071\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27068\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__27093\,
            I => \N__27065\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__27080\,
            I => \N__27060\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__27071\,
            I => \N__27060\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__27068\,
            I => \N__27053\
        );

    \I__5616\ : Span4Mux_h
    port map (
            O => \N__27065\,
            I => \N__27053\
        );

    \I__5615\ : Span4Mux_v
    port map (
            O => \N__27060\,
            I => \N__27053\
        );

    \I__5614\ : Span4Mux_v
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__5613\ : Span4Mux_v
    port map (
            O => \N__27050\,
            I => \N__27047\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__27047\,
            I => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\
        );

    \I__5611\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__27041\,
            I => \N__27038\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__27035\,
            I => \N__27032\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__27029\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\
        );

    \I__5605\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27023\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__27020\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__27020\,
            I => \N__27017\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__27017\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\
        );

    \I__5601\ : CEMux
    port map (
            O => \N__27014\,
            I => \N__27010\
        );

    \I__5600\ : CEMux
    port map (
            O => \N__27013\,
            I => \N__27007\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__27010\,
            I => \N__27004\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__27007\,
            I => \N__27001\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__27004\,
            I => \N__26998\
        );

    \I__5596\ : Span4Mux_v
    port map (
            O => \N__27001\,
            I => \N__26994\
        );

    \I__5595\ : IoSpan4Mux
    port map (
            O => \N__26998\,
            I => \N__26991\
        );

    \I__5594\ : CEMux
    port map (
            O => \N__26997\,
            I => \N__26988\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__26994\,
            I => \N__26983\
        );

    \I__5592\ : Span4Mux_s2_v
    port map (
            O => \N__26991\,
            I => \N__26983\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26980\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__26983\,
            I => \N__26975\
        );

    \I__5589\ : Span4Mux_v
    port map (
            O => \N__26980\,
            I => \N__26975\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__26975\,
            I => \N__26972\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__26972\,
            I => \ppm_encoder_1.N_1014_0\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__26969\,
            I => \N__26965\
        );

    \I__5585\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26962\
        );

    \I__5584\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26959\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__26962\,
            I => \N__26954\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__26959\,
            I => \N__26954\
        );

    \I__5581\ : Span4Mux_v
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__26951\,
            I => \N__26948\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__26948\,
            I => \ppm_encoder_1.N_1014_i\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26945\,
            I => \N__26938\
        );

    \I__5577\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26938\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26935\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26932\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__26935\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__26932\,
            I => \ppm_encoder_1.counterZ0Z_0\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__5571\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26918\
        );

    \I__5570\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26918\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__26915\,
            I => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\
        );

    \I__5567\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__26909\,
            I => \N__26905\
        );

    \I__5565\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26902\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__26905\,
            I => \N__26899\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__26899\,
            I => \N__26893\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__26896\,
            I => scaler_4_data_11
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__26893\,
            I => scaler_4_data_11
        );

    \I__5559\ : InMux
    port map (
            O => \N__26888\,
            I => \scaler_4.un2_source_data_0_cry_6\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__5557\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26876\
        );

    \I__5556\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26876\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__5554\ : Odrv12
    port map (
            O => \N__26873\,
            I => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\
        );

    \I__5553\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26866\
        );

    \I__5552\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26863\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__26866\,
            I => \N__26860\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__26863\,
            I => \N__26857\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__26857\,
            I => \N__26849\
        );

    \I__5547\ : Span4Mux_v
    port map (
            O => \N__26854\,
            I => \N__26849\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__26849\,
            I => scaler_4_data_12
        );

    \I__5545\ : InMux
    port map (
            O => \N__26846\,
            I => \scaler_4.un2_source_data_0_cry_7\
        );

    \I__5544\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26840\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26836\
        );

    \I__5542\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26833\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__26836\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__26833\,
            I => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__5538\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__5536\ : Odrv4
    port map (
            O => \N__26819\,
            I => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__26816\,
            I => \N__26812\
        );

    \I__5534\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26809\
        );

    \I__5533\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26806\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__26809\,
            I => \N__26803\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__26806\,
            I => \N__26798\
        );

    \I__5530\ : Span4Mux_v
    port map (
            O => \N__26803\,
            I => \N__26798\
        );

    \I__5529\ : Span4Mux_v
    port map (
            O => \N__26798\,
            I => \N__26795\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__26795\,
            I => scaler_4_data_13
        );

    \I__5527\ : InMux
    port map (
            O => \N__26792\,
            I => \bfn_7_22_0_\
        );

    \I__5526\ : InMux
    port map (
            O => \N__26789\,
            I => \scaler_4.un2_source_data_0_cry_9\
        );

    \I__5525\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__26783\,
            I => \N__26780\
        );

    \I__5523\ : Span4Mux_v
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__26774\,
            I => scaler_4_data_14
        );

    \I__5520\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26767\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__26770\,
            I => \N__26764\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__26767\,
            I => \N__26759\
        );

    \I__5517\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26754\
        );

    \I__5516\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26754\
        );

    \I__5515\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26751\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__26759\,
            I => \N__26746\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26746\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__26751\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__26746\,
            I => \scaler_4.un2_source_data_0\
        );

    \I__5510\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26735\
        );

    \I__5509\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26732\
        );

    \I__5508\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26729\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__26738\,
            I => \N__26726\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26719\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26719\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26719\
        );

    \I__5503\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26716\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__26719\,
            I => \N__26711\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__26716\,
            I => \N__26711\
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__26711\,
            I => \frame_decoder_OFF4data_0\
        );

    \I__5499\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26703\
        );

    \I__5498\ : InMux
    port map (
            O => \N__26707\,
            I => \N__26700\
        );

    \I__5497\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26697\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__26703\,
            I => \N__26691\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__26700\,
            I => \N__26691\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__26697\,
            I => \N__26688\
        );

    \I__5493\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26685\
        );

    \I__5492\ : Odrv12
    port map (
            O => \N__26691\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__26688\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__26685\,
            I => \frame_decoder_CH4data_0\
        );

    \I__5489\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26674\
        );

    \I__5488\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26671\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__26674\,
            I => \N__26666\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__26671\,
            I => \N__26666\
        );

    \I__5485\ : Odrv12
    port map (
            O => \N__26666\,
            I => \ppm_encoder_1.elevatorZ0Z_4\
        );

    \I__5484\ : CascadeMux
    port map (
            O => \N__26663\,
            I => \N__26659\
        );

    \I__5483\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26656\
        );

    \I__5482\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__26656\,
            I => scaler_4_data_4
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__26653\,
            I => scaler_4_data_4
        );

    \I__5479\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26645\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__26645\,
            I => \N__26642\
        );

    \I__5477\ : Span4Mux_s3_v
    port map (
            O => \N__26642\,
            I => \N__26638\
        );

    \I__5476\ : InMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__26638\,
            I => \N__26632\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26629\
        );

    \I__5473\ : Odrv4
    port map (
            O => \N__26632\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__5472\ : Odrv12
    port map (
            O => \N__26629\,
            I => \ppm_encoder_1.rudderZ0Z_4\
        );

    \I__5471\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__26621\,
            I => \scaler_4.N_905_i_l_ofxZ0\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__26618\,
            I => \N__26615\
        );

    \I__5468\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__26612\,
            I => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\
        );

    \I__5466\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26605\
        );

    \I__5465\ : InMux
    port map (
            O => \N__26608\,
            I => \N__26602\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__26605\,
            I => \N__26599\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__26599\,
            I => \N__26593\
        );

    \I__5461\ : Span4Mux_v
    port map (
            O => \N__26596\,
            I => \N__26588\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__26593\,
            I => \N__26588\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__26588\,
            I => scaler_4_data_6
        );

    \I__5458\ : InMux
    port map (
            O => \N__26585\,
            I => \scaler_4.un2_source_data_0_cry_1\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__5456\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26573\
        );

    \I__5455\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26573\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__26573\,
            I => \N__26570\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__26570\,
            I => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\
        );

    \I__5452\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26563\
        );

    \I__5451\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26560\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__26563\,
            I => \N__26557\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__26560\,
            I => \N__26554\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__26557\,
            I => \N__26551\
        );

    \I__5447\ : Span4Mux_h
    port map (
            O => \N__26554\,
            I => \N__26546\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__26551\,
            I => \N__26546\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__26546\,
            I => scaler_4_data_7
        );

    \I__5444\ : InMux
    port map (
            O => \N__26543\,
            I => \scaler_4.un2_source_data_0_cry_2\
        );

    \I__5443\ : CascadeMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5442\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26531\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26531\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__26528\,
            I => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__26525\,
            I => \N__26521\
        );

    \I__5437\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__5436\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26515\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__26518\,
            I => \N__26512\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__26515\,
            I => \N__26509\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__26512\,
            I => \N__26506\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__26509\,
            I => \N__26503\
        );

    \I__5431\ : Span4Mux_v
    port map (
            O => \N__26506\,
            I => \N__26500\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__26503\,
            I => scaler_4_data_8
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__26500\,
            I => scaler_4_data_8
        );

    \I__5428\ : InMux
    port map (
            O => \N__26495\,
            I => \scaler_4.un2_source_data_0_cry_3\
        );

    \I__5427\ : CascadeMux
    port map (
            O => \N__26492\,
            I => \N__26489\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26483\
        );

    \I__5425\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26483\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__26480\,
            I => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\
        );

    \I__5422\ : InMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__26474\,
            I => \N__26470\
        );

    \I__5420\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26467\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__26470\,
            I => \N__26464\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__5417\ : Span4Mux_h
    port map (
            O => \N__26464\,
            I => \N__26456\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__26461\,
            I => \N__26456\
        );

    \I__5415\ : Span4Mux_v
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__26453\,
            I => scaler_4_data_9
        );

    \I__5413\ : InMux
    port map (
            O => \N__26450\,
            I => \scaler_4.un2_source_data_0_cry_4\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__26447\,
            I => \N__26444\
        );

    \I__5411\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26438\
        );

    \I__5410\ : InMux
    port map (
            O => \N__26443\,
            I => \N__26438\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__5408\ : Odrv12
    port map (
            O => \N__26435\,
            I => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\
        );

    \I__5407\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26428\
        );

    \I__5406\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26425\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__26428\,
            I => \N__26422\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26425\,
            I => \N__26417\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__26422\,
            I => \N__26417\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__26414\,
            I => scaler_4_data_10
        );

    \I__5400\ : InMux
    port map (
            O => \N__26411\,
            I => \scaler_4.un2_source_data_0_cry_5\
        );

    \I__5399\ : InMux
    port map (
            O => \N__26408\,
            I => \scaler_4.un3_source_data_0_cry_0\
        );

    \I__5398\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__5396\ : Odrv4
    port map (
            O => \N__26399\,
            I => \frame_decoder_OFF4data_2\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__5394\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__26390\,
            I => \frame_decoder_CH4data_2\
        );

    \I__5392\ : InMux
    port map (
            O => \N__26387\,
            I => \scaler_4.un3_source_data_0_cry_1\
        );

    \I__5391\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26381\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__26381\,
            I => \frame_decoder_CH4data_3\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__5386\ : Odrv12
    port map (
            O => \N__26369\,
            I => \frame_decoder_OFF4data_3\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26366\,
            I => \scaler_4.un3_source_data_0_cry_2\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__5382\ : Odrv12
    port map (
            O => \N__26357\,
            I => \frame_decoder_OFF4data_4\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__26348\,
            I => \frame_decoder_CH4data_4\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26345\,
            I => \scaler_4.un3_source_data_0_cry_3\
        );

    \I__5377\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26339\,
            I => \frame_decoder_CH4data_5\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5374\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__26330\,
            I => \N__26327\
        );

    \I__5372\ : Odrv12
    port map (
            O => \N__26327\,
            I => \frame_decoder_OFF4data_5\
        );

    \I__5371\ : InMux
    port map (
            O => \N__26324\,
            I => \scaler_4.un3_source_data_0_cry_4\
        );

    \I__5370\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__26318\,
            I => \frame_decoder_CH4data_6\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__5367\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__5365\ : Odrv12
    port map (
            O => \N__26306\,
            I => \frame_decoder_OFF4data_6\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26303\,
            I => \scaler_4.un3_source_data_0_cry_5\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26300\,
            I => \scaler_4.un3_source_data_0_cry_6\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26297\,
            I => \bfn_7_20_0_\
        );

    \I__5361\ : InMux
    port map (
            O => \N__26294\,
            I => \scaler_4.un3_source_data_0_cry_8\
        );

    \I__5360\ : CEMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__26282\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\
        );

    \I__5356\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__26276\,
            I => \frame_decoder_CH4data_1\
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__26264\,
            I => \frame_decoder_OFF4data_1\
        );

    \I__5350\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26256\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26253\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26250\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__26256\,
            I => \N__26245\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__26253\,
            I => \N__26245\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26242\
        );

    \I__5344\ : Span4Mux_h
    port map (
            O => \N__26245\,
            I => \N__26239\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26236\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__26239\,
            I => uart_drone_data_5
        );

    \I__5341\ : Odrv4
    port map (
            O => \N__26236\,
            I => uart_drone_data_5
        );

    \I__5340\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26226\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \N__26222\
        );

    \I__5338\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26219\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__26226\,
            I => \N__26216\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26213\
        );

    \I__5335\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26210\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26207\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__26216\,
            I => \N__26204\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26199\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N__26199\
        );

    \I__5330\ : Span12Mux_s7_h
    port map (
            O => \N__26207\,
            I => \N__26196\
        );

    \I__5329\ : Span4Mux_v
    port map (
            O => \N__26204\,
            I => \N__26193\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__26199\,
            I => \N__26190\
        );

    \I__5327\ : Odrv12
    port map (
            O => \N__26196\,
            I => uart_drone_data_6
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__26193\,
            I => uart_drone_data_6
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__26190\,
            I => uart_drone_data_6
        );

    \I__5324\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26175\
        );

    \I__5322\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26172\
        );

    \I__5321\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26169\
        );

    \I__5320\ : Span4Mux_h
    port map (
            O => \N__26175\,
            I => \N__26166\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26163\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__26169\,
            I => \N__26160\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26157\
        );

    \I__5316\ : Span12Mux_s7_h
    port map (
            O => \N__26163\,
            I => \N__26154\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__26160\,
            I => \N__26151\
        );

    \I__5314\ : Odrv4
    port map (
            O => \N__26157\,
            I => uart_drone_data_7
        );

    \I__5313\ : Odrv12
    port map (
            O => \N__26154\,
            I => uart_drone_data_7
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__26151\,
            I => uart_drone_data_7
        );

    \I__5311\ : CascadeMux
    port map (
            O => \N__26144\,
            I => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\
        );

    \I__5310\ : IoInMux
    port map (
            O => \N__26141\,
            I => \N__26138\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26135\
        );

    \I__5308\ : Span12Mux_s4_v
    port map (
            O => \N__26135\,
            I => \N__26132\
        );

    \I__5307\ : Span12Mux_v
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__5306\ : Odrv12
    port map (
            O => \N__26129\,
            I => \GB_BUFFER_reset_system_g_THRU_CO\
        );

    \I__5305\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26122\
        );

    \I__5304\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26119\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__26122\,
            I => \N__26115\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26119\,
            I => \N__26112\
        );

    \I__5301\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26109\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__26115\,
            I => \N__26106\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__26112\,
            I => \N__26101\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__26109\,
            I => \N__26101\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__26106\,
            I => \N__26098\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__26101\,
            I => \N__26095\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__26098\,
            I => uart_drone_data_0
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__26095\,
            I => uart_drone_data_0
        );

    \I__5293\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26086\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26083\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__26086\,
            I => \N__26076\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__26083\,
            I => \N__26076\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26073\
        );

    \I__5288\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26070\
        );

    \I__5287\ : Span4Mux_v
    port map (
            O => \N__26076\,
            I => \N__26067\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__26073\,
            I => \N__26062\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__26070\,
            I => \N__26062\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__26067\,
            I => \N__26059\
        );

    \I__5283\ : Span4Mux_h
    port map (
            O => \N__26062\,
            I => \N__26056\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__26059\,
            I => uart_drone_data_1
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__26056\,
            I => uart_drone_data_1
        );

    \I__5280\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26047\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__26050\,
            I => \N__26043\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26040\
        );

    \I__5277\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26037\
        );

    \I__5276\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26034\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__26040\,
            I => \N__26031\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__26037\,
            I => \N__26028\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__26034\,
            I => \N__26025\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__26031\,
            I => \N__26022\
        );

    \I__5271\ : Span4Mux_h
    port map (
            O => \N__26028\,
            I => \N__26019\
        );

    \I__5270\ : Span4Mux_h
    port map (
            O => \N__26025\,
            I => \N__26016\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__26022\,
            I => uart_drone_data_2
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__26019\,
            I => uart_drone_data_2
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__26016\,
            I => uart_drone_data_2
        );

    \I__5266\ : InMux
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__26006\,
            I => \N__26000\
        );

    \I__5264\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25997\
        );

    \I__5263\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25994\
        );

    \I__5262\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25991\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__26000\,
            I => \N__25988\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25985\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25980\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25980\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__25988\,
            I => \N__25977\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__25985\,
            I => \N__25974\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__25980\,
            I => \N__25971\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__25977\,
            I => uart_drone_data_3
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__25974\,
            I => uart_drone_data_3
        );

    \I__5252\ : Odrv4
    port map (
            O => \N__25971\,
            I => uart_drone_data_3
        );

    \I__5251\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25959\
        );

    \I__5250\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25955\
        );

    \I__5249\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25952\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25949\
        );

    \I__5247\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25946\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__25955\,
            I => \N__25943\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__25952\,
            I => \N__25940\
        );

    \I__5244\ : Span4Mux_v
    port map (
            O => \N__25949\,
            I => \N__25937\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__25946\,
            I => \N__25934\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__25943\,
            I => \N__25931\
        );

    \I__5241\ : Span4Mux_v
    port map (
            O => \N__25940\,
            I => \N__25928\
        );

    \I__5240\ : Span4Mux_v
    port map (
            O => \N__25937\,
            I => \N__25923\
        );

    \I__5239\ : Span4Mux_v
    port map (
            O => \N__25934\,
            I => \N__25923\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__25931\,
            I => uart_drone_data_4
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__25928\,
            I => uart_drone_data_4
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__25923\,
            I => uart_drone_data_4
        );

    \I__5235\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25907\
        );

    \I__5233\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25902\
        );

    \I__5232\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25902\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__25910\,
            I => \N__25898\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__25907\,
            I => \N__25892\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25892\
        );

    \I__5228\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25885\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25885\
        );

    \I__5226\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25885\
        );

    \I__5225\ : Span4Mux_v
    port map (
            O => \N__25892\,
            I => \N__25882\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__25885\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__25882\,
            I => \dron_frame_decoder_1.stateZ0Z_6\
        );

    \I__5222\ : CEMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__25874\,
            I => \N__25871\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__25868\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__25865\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\
        );

    \I__5217\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__25859\,
            I => \Commands_frame_decoder.state_ns_0_a3_0_3_2\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__5214\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25847\
        );

    \I__5213\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25847\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__25847\,
            I => \Commands_frame_decoder.stateZ0Z_2\
        );

    \I__5211\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25832\
        );

    \I__5210\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25832\
        );

    \I__5209\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25832\
        );

    \I__5208\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25832\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__25829\,
            I => \N__25825\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25822\
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__25825\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__25822\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__25817\,
            I => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\
        );

    \I__5201\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25810\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25807\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__25810\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__25807\,
            I => \Commands_frame_decoder.stateZ0Z_3\
        );

    \I__5197\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__25793\,
            I => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\
        );

    \I__5193\ : InMux
    port map (
            O => \N__25790\,
            I => \ppm_encoder_1.un1_rudder_cry_12\
        );

    \I__5192\ : InMux
    port map (
            O => \N__25787\,
            I => \bfn_5_30_0_\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__5190\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25774\
        );

    \I__5188\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__25774\,
            I => \N__25768\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__5184\ : Odrv12
    port map (
            O => \N__25765\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__25762\,
            I => \ppm_encoder_1.rudderZ0Z_14\
        );

    \I__5182\ : CEMux
    port map (
            O => \N__25757\,
            I => \N__25751\
        );

    \I__5181\ : CEMux
    port map (
            O => \N__25756\,
            I => \N__25748\
        );

    \I__5180\ : CEMux
    port map (
            O => \N__25755\,
            I => \N__25745\
        );

    \I__5179\ : CEMux
    port map (
            O => \N__25754\,
            I => \N__25742\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25739\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__25748\,
            I => \N__25736\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__25745\,
            I => \N__25733\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__25742\,
            I => \N__25730\
        );

    \I__5174\ : Span4Mux_v
    port map (
            O => \N__25739\,
            I => \N__25725\
        );

    \I__5173\ : Span4Mux_s3_h
    port map (
            O => \N__25736\,
            I => \N__25725\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__25733\,
            I => \N__25722\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__25730\,
            I => \N__25719\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__25725\,
            I => \N__25716\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__25722\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__25719\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__25716\,
            I => \Commands_frame_decoder.state_RNIF38SZ0Z_6\
        );

    \I__5166\ : CEMux
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__25706\,
            I => \N__25700\
        );

    \I__5164\ : CEMux
    port map (
            O => \N__25705\,
            I => \N__25697\
        );

    \I__5163\ : CEMux
    port map (
            O => \N__25704\,
            I => \N__25694\
        );

    \I__5162\ : CEMux
    port map (
            O => \N__25703\,
            I => \N__25691\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__25700\,
            I => \N__25686\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__25697\,
            I => \N__25686\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__25694\,
            I => \N__25683\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__25691\,
            I => \N__25680\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__25686\,
            I => \N__25677\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__25683\,
            I => \N__25674\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__25680\,
            I => \N__25671\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__25677\,
            I => \N__25668\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__25674\,
            I => \N__25665\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__25671\,
            I => \N__25660\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__25668\,
            I => \N__25660\
        );

    \I__5150\ : Odrv4
    port map (
            O => \N__25665\,
            I => \dron_frame_decoder_1.N_390_0\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__25660\,
            I => \dron_frame_decoder_1.N_390_0\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__25655\,
            I => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\
        );

    \I__5147\ : CEMux
    port map (
            O => \N__25652\,
            I => \N__25649\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25645\
        );

    \I__5145\ : CEMux
    port map (
            O => \N__25648\,
            I => \N__25642\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__25645\,
            I => \N__25637\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25637\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__25637\,
            I => \N__25633\
        );

    \I__5141\ : CEMux
    port map (
            O => \N__25636\,
            I => \N__25630\
        );

    \I__5140\ : Span4Mux_h
    port map (
            O => \N__25633\,
            I => \N__25627\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__25630\,
            I => \N__25624\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__25627\,
            I => \dron_frame_decoder_1.N_382_0\
        );

    \I__5137\ : Odrv12
    port map (
            O => \N__25624\,
            I => \dron_frame_decoder_1.N_382_0\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__25619\,
            I => \N__25614\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__25618\,
            I => \N__25611\
        );

    \I__5134\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25604\
        );

    \I__5133\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25604\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25611\,
            I => \N__25604\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__25604\,
            I => \dron_frame_decoder_1.stateZ0Z_7\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25598\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__25598\,
            I => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__25589\,
            I => \N__25586\
        );

    \I__5125\ : Span4Mux_v
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__5124\ : Odrv4
    port map (
            O => \N__25583\,
            I => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25580\,
            I => \ppm_encoder_1.un1_rudder_cry_6\
        );

    \I__5122\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25574\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__5120\ : Span4Mux_v
    port map (
            O => \N__25571\,
            I => \N__25568\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__25565\,
            I => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25562\,
            I => \ppm_encoder_1.un1_rudder_cry_7\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__5115\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__25547\,
            I => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25544\,
            I => \ppm_encoder_1.un1_rudder_cry_8\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25538\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__5108\ : Odrv12
    port map (
            O => \N__25535\,
            I => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25532\,
            I => \ppm_encoder_1.un1_rudder_cry_9\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__5105\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25523\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__5102\ : Span4Mux_v
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__25514\,
            I => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\
        );

    \I__5100\ : InMux
    port map (
            O => \N__25511\,
            I => \ppm_encoder_1.un1_rudder_cry_10\
        );

    \I__5099\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__5097\ : Span12Mux_v
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__5096\ : Odrv12
    port map (
            O => \N__25499\,
            I => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\
        );

    \I__5095\ : InMux
    port map (
            O => \N__25496\,
            I => \ppm_encoder_1.un1_rudder_cry_11\
        );

    \I__5094\ : InMux
    port map (
            O => \N__25493\,
            I => \ppm_encoder_1.counter24_0_N_2\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25482\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25477\
        );

    \I__5090\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25477\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25482\,
            I => \N__25474\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__25477\,
            I => \N__25471\
        );

    \I__5087\ : Span4Mux_h
    port map (
            O => \N__25474\,
            I => \N__25468\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__25471\,
            I => \N__25465\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__25468\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__25465\,
            I => \ppm_encoder_1.init_pulsesZ0Z_10\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25452\
        );

    \I__5081\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25449\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__25455\,
            I => \N__25446\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__25452\,
            I => \N__25443\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25440\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25437\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__25443\,
            I => \N__25434\
        );

    \I__5075\ : Span4Mux_h
    port map (
            O => \N__25440\,
            I => \N__25431\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__25437\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__25434\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__25431\,
            I => \ppm_encoder_1.rudderZ0Z_10\
        );

    \I__5071\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__25418\,
            I => \N__25415\
        );

    \I__5068\ : Odrv4
    port map (
            O => \N__25415\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25408\
        );

    \I__5066\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25405\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__25408\,
            I => \N__25402\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25405\,
            I => \ppm_encoder_1.N_238\
        );

    \I__5063\ : Odrv4
    port map (
            O => \N__25402\,
            I => \ppm_encoder_1.N_238\
        );

    \I__5062\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25392\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25389\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25386\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__25392\,
            I => \N__25383\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__25389\,
            I => \N__25377\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__25386\,
            I => \N__25377\
        );

    \I__5056\ : Span4Mux_s2_v
    port map (
            O => \N__25383\,
            I => \N__25374\
        );

    \I__5055\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25371\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__25377\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5053\ : Odrv4
    port map (
            O => \N__25374\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__25371\,
            I => \ppm_encoder_1.counter24_0_N_2_THRU_CO\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__25364\,
            I => \N__25359\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__25363\,
            I => \N__25354\
        );

    \I__5049\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25351\
        );

    \I__5048\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25348\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25341\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25341\
        );

    \I__5045\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25341\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25338\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__25348\,
            I => \N__25335\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__25341\,
            I => \N__25330\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__25338\,
            I => \N__25325\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__25335\,
            I => \N__25325\
        );

    \I__5039\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25320\
        );

    \I__5038\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25320\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__25330\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__25325\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__25320\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_0\
        );

    \I__5034\ : IoInMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__5032\ : Span4Mux_s2_v
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__5031\ : Sp12to4
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__5030\ : Odrv12
    port map (
            O => \N__25301\,
            I => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\
        );

    \I__5029\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25293\
        );

    \I__5028\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25289\
        );

    \I__5027\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25286\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__25293\,
            I => \N__25283\
        );

    \I__5025\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25280\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__25289\,
            I => \N__25274\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25274\
        );

    \I__5022\ : Span4Mux_s3_v
    port map (
            O => \N__25283\,
            I => \N__25271\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25268\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25279\,
            I => \N__25263\
        );

    \I__5019\ : Span4Mux_s3_v
    port map (
            O => \N__25274\,
            I => \N__25260\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__25271\,
            I => \N__25255\
        );

    \I__5017\ : Span4Mux_s3_v
    port map (
            O => \N__25268\,
            I => \N__25255\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25267\,
            I => \N__25252\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25249\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__25263\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__5013\ : Odrv4
    port map (
            O => \N__25260\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__25255\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__25252\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__25249\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\
        );

    \I__5009\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25233\
        );

    \I__5008\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25230\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__25236\,
            I => \N__25226\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25222\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25230\,
            I => \N__25219\
        );

    \I__5004\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25216\
        );

    \I__5003\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25210\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25210\
        );

    \I__5001\ : Span4Mux_s2_v
    port map (
            O => \N__25222\,
            I => \N__25207\
        );

    \I__5000\ : Span4Mux_s2_v
    port map (
            O => \N__25219\,
            I => \N__25202\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__25216\,
            I => \N__25202\
        );

    \I__4998\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25199\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25210\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__25207\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__25202\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__25199\,
            I => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\
        );

    \I__4993\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25181\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25176\
        );

    \I__4990\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25176\
        );

    \I__4989\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25173\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__25181\,
            I => \N__25168\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25168\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__25173\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__25168\,
            I => \ppm_encoder_1.init_pulsesZ0Z_3\
        );

    \I__4984\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25160\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__25160\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\
        );

    \I__4982\ : InMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__25154\,
            I => \ppm_encoder_1.pulses2countZ0Z_0\
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__25151\,
            I => \N__25148\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25145\,
            I => \ppm_encoder_1.pulses2countZ0Z_1\
        );

    \I__4977\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25136\
        );

    \I__4976\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25136\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__25136\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\
        );

    \I__4974\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__25130\,
            I => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__4971\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__25121\,
            I => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__25115\,
            I => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__25109\,
            I => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\
        );

    \I__4965\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__25103\,
            I => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\
        );

    \I__4963\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__4961\ : Odrv4
    port map (
            O => \N__25094\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__4959\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__4957\ : Span4Mux_v
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__25079\,
            I => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\
        );

    \I__4955\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__25070\,
            I => \N__25066\
        );

    \I__4952\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25063\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__25066\,
            I => throttle_command_1
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__25063\,
            I => throttle_command_1
        );

    \I__4949\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__25055\,
            I => \N__25050\
        );

    \I__4947\ : InMux
    port map (
            O => \N__25054\,
            I => \N__25047\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25044\
        );

    \I__4945\ : Span4Mux_h
    port map (
            O => \N__25050\,
            I => \N__25041\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__25047\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25044\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__25041\,
            I => \ppm_encoder_1.throttleZ0Z_1\
        );

    \I__4941\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__25025\,
            I => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\
        );

    \I__4937\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25018\
        );

    \I__4936\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25015\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__25018\,
            I => \N__25012\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__25012\,
            I => \N__25004\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__25009\,
            I => \N__25004\
        );

    \I__4931\ : Odrv4
    port map (
            O => \N__25004\,
            I => throttle_command_3
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__25001\,
            I => \N__24993\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__25000\,
            I => \N__24988\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__24999\,
            I => \N__24977\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__24998\,
            I => \N__24974\
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__24997\,
            I => \N__24967\
        );

    \I__4925\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24964\
        );

    \I__4924\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24957\
        );

    \I__4923\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24957\
        );

    \I__4922\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24957\
        );

    \I__4921\ : InMux
    port map (
            O => \N__24988\,
            I => \N__24948\
        );

    \I__4920\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24948\
        );

    \I__4919\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24948\
        );

    \I__4918\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24948\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__24984\,
            I => \N__24933\
        );

    \I__4916\ : CascadeMux
    port map (
            O => \N__24983\,
            I => \N__24930\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__24982\,
            I => \N__24925\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__24981\,
            I => \N__24922\
        );

    \I__4913\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24914\
        );

    \I__4912\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24914\
        );

    \I__4911\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24914\
        );

    \I__4910\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24909\
        );

    \I__4909\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24909\
        );

    \I__4908\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24902\
        );

    \I__4907\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24902\
        );

    \I__4906\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24902\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__24964\,
            I => \N__24897\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__24957\,
            I => \N__24897\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__24948\,
            I => \N__24894\
        );

    \I__4902\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24883\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24883\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24883\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24883\
        );

    \I__4898\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24883\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__24942\,
            I => \N__24880\
        );

    \I__4896\ : CascadeMux
    port map (
            O => \N__24941\,
            I => \N__24876\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__24940\,
            I => \N__24873\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__24939\,
            I => \N__24870\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__24938\,
            I => \N__24867\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__24937\,
            I => \N__24864\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__24936\,
            I => \N__24861\
        );

    \I__4890\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24855\
        );

    \I__4889\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24850\
        );

    \I__4888\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24850\
        );

    \I__4887\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24841\
        );

    \I__4886\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24841\
        );

    \I__4885\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24841\
        );

    \I__4884\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24841\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__24914\,
            I => \N__24836\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__24909\,
            I => \N__24836\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__24902\,
            I => \N__24831\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__24897\,
            I => \N__24831\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__24894\,
            I => \N__24826\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N__24826\
        );

    \I__4877\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24823\
        );

    \I__4876\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24816\
        );

    \I__4875\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24816\
        );

    \I__4874\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24816\
        );

    \I__4873\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24801\
        );

    \I__4872\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24801\
        );

    \I__4871\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24801\
        );

    \I__4870\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24801\
        );

    \I__4869\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24801\
        );

    \I__4868\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24801\
        );

    \I__4867\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24801\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__24855\,
            I => \N__24796\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24796\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24793\
        );

    \I__4863\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24786\
        );

    \I__4862\ : Span4Mux_v
    port map (
            O => \N__24831\,
            I => \N__24786\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__24826\,
            I => \N__24786\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__24823\,
            I => pid_altitude_dv
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__24816\,
            I => pid_altitude_dv
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__24801\,
            I => pid_altitude_dv
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__24796\,
            I => pid_altitude_dv
        );

    \I__4856\ : Odrv12
    port map (
            O => \N__24793\,
            I => pid_altitude_dv
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__24786\,
            I => pid_altitude_dv
        );

    \I__4854\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24765\
        );

    \I__4852\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24762\
        );

    \I__4851\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24759\
        );

    \I__4850\ : Span4Mux_s2_v
    port map (
            O => \N__24765\,
            I => \N__24756\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24753\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__24759\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__24756\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__4846\ : Odrv12
    port map (
            O => \N__24753\,
            I => \ppm_encoder_1.throttleZ0Z_3\
        );

    \I__4845\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24743\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\
        );

    \I__4843\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__4842\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24729\
        );

    \I__4841\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24729\
        );

    \I__4840\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24726\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__24734\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__24729\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24726\,
            I => \ppm_encoder_1.PPM_STATEZ0Z_1\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__24719\,
            I => \ppm_encoder_1.N_140_0_cascade_\
        );

    \I__4835\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__24713\,
            I => \ppm_encoder_1.N_145\
        );

    \I__4833\ : IoInMux
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__4831\ : Span4Mux_s0_v
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__4830\ : Sp12to4
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__4829\ : Span12Mux_h
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__4828\ : Span12Mux_v
    port map (
            O => \N__24695\,
            I => \N__24692\
        );

    \I__4827\ : Span12Mux_v
    port map (
            O => \N__24692\,
            I => \N__24688\
        );

    \I__4826\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24685\
        );

    \I__4825\ : Odrv12
    port map (
            O => \N__24688\,
            I => ppm_output_c
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__24685\,
            I => ppm_output_c
        );

    \I__4823\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24677\,
            I => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\
        );

    \I__4821\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24671\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__24668\,
            I => \ppm_encoder_1.pulses2countZ0Z_3\
        );

    \I__4818\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24662\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__24662\,
            I => \N__24659\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__24659\,
            I => \ppm_encoder_1.pulses2countZ0Z_2\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24649\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24646\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__24649\,
            I => \N__24643\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24640\
        );

    \I__4810\ : Sp12to4
    port map (
            O => \N__24643\,
            I => \N__24635\
        );

    \I__4809\ : Sp12to4
    port map (
            O => \N__24640\,
            I => \N__24635\
        );

    \I__4808\ : Odrv12
    port map (
            O => \N__24635\,
            I => scaler_2_data_6
        );

    \I__4807\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24629\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__4804\ : Span4Mux_v
    port map (
            O => \N__24623\,
            I => \N__24618\
        );

    \I__4803\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24613\
        );

    \I__4802\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24613\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__24618\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__24613\,
            I => \ppm_encoder_1.init_pulsesZ0Z_6\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__24608\,
            I => \N__24603\
        );

    \I__4798\ : InMux
    port map (
            O => \N__24607\,
            I => \N__24600\
        );

    \I__4797\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24595\
        );

    \I__4796\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24595\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__24600\,
            I => \N__24592\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__24595\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__24592\,
            I => \ppm_encoder_1.rudderZ0Z_6\
        );

    \I__4792\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__24581\,
            I => \N__24577\
        );

    \I__4789\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24574\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__24577\,
            I => \N__24568\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24568\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24565\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__24568\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__24565\,
            I => \ppm_encoder_1.init_pulsesZ0Z_13\
        );

    \I__4783\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24556\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__24559\,
            I => \N__24552\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__24556\,
            I => \N__24549\
        );

    \I__4780\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24544\
        );

    \I__4779\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24544\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__24549\,
            I => \N__24541\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24544\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__24541\,
            I => \ppm_encoder_1.rudderZ0Z_13\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__4773\ : Span4Mux_h
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__24527\,
            I => \N__24523\
        );

    \I__4771\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24520\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__24523\,
            I => throttle_command_0
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__24520\,
            I => throttle_command_0
        );

    \I__4768\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24509\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24509\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24504\
        );

    \I__4765\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24499\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24499\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__24504\,
            I => \N__24496\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__24499\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__24496\,
            I => \ppm_encoder_1.throttleZ0Z_0\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24488\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__24488\,
            I => \N__24485\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__4757\ : Span4Mux_v
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__24479\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__24473\,
            I => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\
        );

    \I__4753\ : InMux
    port map (
            O => \N__24470\,
            I => \ppm_encoder_1.un1_elevator_cry_7\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__4751\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__24458\,
            I => \N__24455\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__24455\,
            I => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\
        );

    \I__4747\ : InMux
    port map (
            O => \N__24452\,
            I => \ppm_encoder_1.un1_elevator_cry_8\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__24446\,
            I => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24443\,
            I => \ppm_encoder_1.un1_elevator_cry_9\
        );

    \I__4743\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24434\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__24434\,
            I => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\
        );

    \I__4740\ : InMux
    port map (
            O => \N__24431\,
            I => \ppm_encoder_1.un1_elevator_cry_10\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__24425\,
            I => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\
        );

    \I__4737\ : InMux
    port map (
            O => \N__24422\,
            I => \ppm_encoder_1.un1_elevator_cry_11\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__24416\,
            I => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\
        );

    \I__4734\ : InMux
    port map (
            O => \N__24413\,
            I => \ppm_encoder_1.un1_elevator_cry_12\
        );

    \I__4733\ : InMux
    port map (
            O => \N__24410\,
            I => \bfn_5_23_0_\
        );

    \I__4732\ : InMux
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__24404\,
            I => \N__24400\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24397\
        );

    \I__4729\ : Span4Mux_v
    port map (
            O => \N__24400\,
            I => \N__24392\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__24397\,
            I => \N__24392\
        );

    \I__4727\ : Span4Mux_h
    port map (
            O => \N__24392\,
            I => \N__24389\
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__24389\,
            I => \ppm_encoder_1.elevatorZ0Z_14\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__24386\,
            I => \N__24382\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24378\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24375\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24371\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24378\,
            I => \N__24368\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__24375\,
            I => \N__24365\
        );

    \I__4719\ : InMux
    port map (
            O => \N__24374\,
            I => \N__24362\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24359\
        );

    \I__4717\ : Span4Mux_h
    port map (
            O => \N__24368\,
            I => \N__24352\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__24365\,
            I => \N__24352\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24352\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__24359\,
            I => \N__24349\
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__24352\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__24349\,
            I => \ppm_encoder_1.init_pulsesZ0Z_0\
        );

    \I__4711\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__24338\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__24329\,
            I => \N__24324\
        );

    \I__4705\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24321\
        );

    \I__4704\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24318\
        );

    \I__4703\ : Span4Mux_s2_h
    port map (
            O => \N__24324\,
            I => \N__24315\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24321\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__24318\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__24315\,
            I => \ppm_encoder_1.elevatorZ0Z_13\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24297\
        );

    \I__4696\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24294\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24291\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__24297\,
            I => \N__24288\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24285\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24282\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__24288\,
            I => \N__24279\
        );

    \I__4690\ : Span4Mux_s2_v
    port map (
            O => \N__24285\,
            I => \N__24276\
        );

    \I__4689\ : Span12Mux_v
    port map (
            O => \N__24282\,
            I => \N__24273\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__24279\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__24276\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4686\ : Odrv12
    port map (
            O => \N__24273\,
            I => \ppm_encoder_1.init_pulsesZ0Z_14\
        );

    \I__4685\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__4683\ : Span4Mux_v
    port map (
            O => \N__24260\,
            I => \N__24255\
        );

    \I__4682\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24252\
        );

    \I__4681\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24249\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__24255\,
            I => \N__24244\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24244\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24249\,
            I => \N__24241\
        );

    \I__4677\ : Odrv4
    port map (
            O => \N__24244\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__24241\,
            I => \ppm_encoder_1.init_pulsesZ0Z_8\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \N__24233\
        );

    \I__4674\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24230\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24227\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__24227\,
            I => \N__24222\
        );

    \I__4671\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24217\
        );

    \I__4670\ : InMux
    port map (
            O => \N__24225\,
            I => \N__24217\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__24222\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__24217\,
            I => \ppm_encoder_1.rudderZ0Z_8\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__4665\ : Sp12to4
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__4664\ : Odrv12
    port map (
            O => \N__24203\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\
        );

    \I__4663\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24196\
        );

    \I__4662\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24193\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24190\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N__24187\
        );

    \I__4659\ : Span4Mux_v
    port map (
            O => \N__24190\,
            I => \N__24184\
        );

    \I__4658\ : Span12Mux_v
    port map (
            O => \N__24187\,
            I => \N__24181\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__24184\,
            I => scaler_2_data_10
        );

    \I__4656\ : Odrv12
    port map (
            O => \N__24181\,
            I => scaler_2_data_10
        );

    \I__4655\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24173\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24170\
        );

    \I__4653\ : Span4Mux_h
    port map (
            O => \N__24170\,
            I => \N__24167\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__24167\,
            I => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\
        );

    \I__4651\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__24161\,
            I => \N__24157\
        );

    \I__4649\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24154\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__24157\,
            I => \N__24148\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24148\
        );

    \I__4646\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24145\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__24148\,
            I => \N__24142\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__24145\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__4643\ : Odrv4
    port map (
            O => \N__24142\,
            I => \ppm_encoder_1.aileronZ0Z_10\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24134\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__24134\,
            I => \N__24130\
        );

    \I__4640\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24127\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__24130\,
            I => \N__24122\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24122\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__24122\,
            I => \N__24119\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__24119\,
            I => scaler_2_data_13
        );

    \I__4635\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__4633\ : Odrv12
    port map (
            O => \N__24110\,
            I => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__24104\,
            I => \N__24100\
        );

    \I__4630\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24097\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__24100\,
            I => \N__24091\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__24097\,
            I => \N__24091\
        );

    \I__4627\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24088\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__24091\,
            I => \N__24085\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__24088\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__24085\,
            I => \ppm_encoder_1.elevatorZ0Z_10\
        );

    \I__4623\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24077\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__24071\,
            I => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24068\,
            I => \ppm_encoder_1.un1_elevator_cry_6\
        );

    \I__4618\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24059\
        );

    \I__4617\ : InMux
    port map (
            O => \N__24064\,
            I => \N__24054\
        );

    \I__4616\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24054\
        );

    \I__4615\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24051\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__24059\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__24054\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__24051\,
            I => \dron_frame_decoder_1.stateZ0Z_0\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__24044\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\
        );

    \I__4610\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24035\
        );

    \I__4609\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24035\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__24035\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_1\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__24032\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__24029\,
            I => \N__24025\
        );

    \I__4605\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24021\
        );

    \I__4604\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24018\
        );

    \I__4603\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24015\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__24021\,
            I => \N__24012\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__24009\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__24015\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__24012\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__24009\,
            I => \dron_frame_decoder_1.stateZ0Z_1\
        );

    \I__4597\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__23999\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3\
        );

    \I__4595\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23992\
        );

    \I__4594\ : IoInMux
    port map (
            O => \N__23995\,
            I => \N__23989\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__23992\,
            I => \N__23986\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23982\
        );

    \I__4591\ : Span4Mux_v
    port map (
            O => \N__23986\,
            I => \N__23978\
        );

    \I__4590\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23975\
        );

    \I__4589\ : Span12Mux_s9_v
    port map (
            O => \N__23982\,
            I => \N__23972\
        );

    \I__4588\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23969\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__23978\,
            I => \N__23964\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__23975\,
            I => \N__23964\
        );

    \I__4585\ : Odrv12
    port map (
            O => \N__23972\,
            I => \debug_CH1_0A_c\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__23969\,
            I => \debug_CH1_0A_c\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__23964\,
            I => \debug_CH1_0A_c\
        );

    \I__4582\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23944\
        );

    \I__4581\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23941\
        );

    \I__4580\ : CascadeMux
    port map (
            O => \N__23955\,
            I => \N__23936\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__23954\,
            I => \N__23933\
        );

    \I__4578\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23917\
        );

    \I__4577\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23917\
        );

    \I__4576\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23917\
        );

    \I__4575\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23917\
        );

    \I__4574\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23917\
        );

    \I__4573\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23917\
        );

    \I__4572\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23917\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__23944\,
            I => \N__23914\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23909\
        );

    \I__4569\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23898\
        );

    \I__4568\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23898\
        );

    \I__4567\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23898\
        );

    \I__4566\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23898\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23898\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23895\
        );

    \I__4563\ : Span4Mux_v
    port map (
            O => \N__23914\,
            I => \N__23892\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23887\
        );

    \I__4561\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23887\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__23909\,
            I => \N__23882\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__23898\,
            I => \N__23879\
        );

    \I__4558\ : Span4Mux_v
    port map (
            O => \N__23895\,
            I => \N__23872\
        );

    \I__4557\ : Span4Mux_v
    port map (
            O => \N__23892\,
            I => \N__23872\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23872\
        );

    \I__4555\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23864\
        );

    \I__4554\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23861\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__23882\,
            I => \N__23858\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__23879\,
            I => \N__23853\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__23872\,
            I => \N__23853\
        );

    \I__4550\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23846\
        );

    \I__4549\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23846\
        );

    \I__4548\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23846\
        );

    \I__4547\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23843\
        );

    \I__4546\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23840\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__23864\,
            I => \pid_alt.N_60_i\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__23861\,
            I => \pid_alt.N_60_i\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__23858\,
            I => \pid_alt.N_60_i\
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__23853\,
            I => \pid_alt.N_60_i\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__23846\,
            I => \pid_alt.N_60_i\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__23843\,
            I => \pid_alt.N_60_i\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__23840\,
            I => \pid_alt.N_60_i\
        );

    \I__4538\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23822\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__23822\,
            I => \pid_alt.state_RNIFCSD1Z0Z_0\
        );

    \I__4536\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23814\
        );

    \I__4535\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23811\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__23817\,
            I => \N__23808\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__23814\,
            I => \N__23805\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__23811\,
            I => \N__23801\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23798\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__23805\,
            I => \N__23795\
        );

    \I__4529\ : InMux
    port map (
            O => \N__23804\,
            I => \N__23792\
        );

    \I__4528\ : Span12Mux_v
    port map (
            O => \N__23801\,
            I => \N__23787\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23787\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__23795\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__23792\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__4524\ : Odrv12
    port map (
            O => \N__23787\,
            I => \frame_decoder_OFF2data_0\
        );

    \I__4523\ : InMux
    port map (
            O => \N__23780\,
            I => \N__23776\
        );

    \I__4522\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23773\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__23776\,
            I => \N__23770\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__23773\,
            I => \N__23766\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__23770\,
            I => \N__23763\
        );

    \I__4518\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23759\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__23766\,
            I => \N__23754\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__23763\,
            I => \N__23754\
        );

    \I__4515\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23751\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23748\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__23754\,
            I => \frame_decoder_CH2data_0\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__23751\,
            I => \frame_decoder_CH2data_0\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__23748\,
            I => \frame_decoder_CH2data_0\
        );

    \I__4510\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23734\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__23737\,
            I => \N__23731\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__4506\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23725\
        );

    \I__4505\ : Odrv4
    port map (
            O => \N__23728\,
            I => scaler_2_data_4
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__23725\,
            I => scaler_2_data_4
        );

    \I__4503\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__23711\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\
        );

    \I__4499\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23701\
        );

    \I__4497\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__23701\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__23698\,
            I => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23685\
        );

    \I__4492\ : InMux
    port map (
            O => \N__23689\,
            I => \N__23682\
        );

    \I__4491\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23679\
        );

    \I__4490\ : Span4Mux_h
    port map (
            O => \N__23685\,
            I => \N__23676\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__23682\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__23679\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__23676\,
            I => \ppm_encoder_1.throttleZ0Z_13\
        );

    \I__4486\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__23663\,
            I => \frame_decoder_OFF2data_5\
        );

    \I__4483\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__23654\,
            I => \frame_decoder_OFF2data_6\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23645\
        );

    \I__4479\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23645\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__23645\,
            I => \frame_decoder_OFF2data_7\
        );

    \I__4477\ : CEMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4474\ : Span4Mux_h
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__23630\,
            I => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__23621\,
            I => \dron_frame_decoder_1.state_RNO_1Z0Z_0\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__23612\,
            I => \dron_frame_decoder_1.N_194_4\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__4465\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23603\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__23600\,
            I => \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\
        );

    \I__4462\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__23594\,
            I => \dron_frame_decoder_1.state_RNO_0Z0Z_0\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__23591\,
            I => \N__23588\
        );

    \I__4459\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__4457\ : Odrv12
    port map (
            O => \N__23582\,
            I => alt_command_5
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__23570\,
            I => alt_command_6
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__4451\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__23558\,
            I => alt_command_7
        );

    \I__4448\ : CEMux
    port map (
            O => \N__23555\,
            I => \N__23552\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__23552\,
            I => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__4445\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__4443\ : Odrv12
    port map (
            O => \N__23540\,
            I => \frame_decoder_OFF2data_1\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__4441\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__23528\,
            I => \frame_decoder_OFF2data_2\
        );

    \I__4438\ : CascadeMux
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23519\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__23516\,
            I => \frame_decoder_OFF2data_3\
        );

    \I__4434\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__23510\,
            I => \N__23507\
        );

    \I__4432\ : Span4Mux_s3_h
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__23504\,
            I => \frame_decoder_OFF2data_4\
        );

    \I__4430\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__23498\,
            I => \dron_frame_decoder_1.drone_altitude_4\
        );

    \I__4428\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__23489\,
            I => drone_altitude_i_4
        );

    \I__4425\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__23483\,
            I => \dron_frame_decoder_1.drone_altitude_5\
        );

    \I__4423\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__23477\,
            I => \N__23474\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__23474\,
            I => drone_altitude_i_5
        );

    \I__4420\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__23468\,
            I => \dron_frame_decoder_1.drone_altitude_6\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__23459\,
            I => drone_altitude_i_6
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__4414\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__4412\ : Span4Mux_s3_h
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__23444\,
            I => alt_command_4
        );

    \I__4410\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__4408\ : Span4Mux_v
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__23432\,
            I => \ppm_encoder_1.N_301\
        );

    \I__4406\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__4404\ : Span4Mux_h
    port map (
            O => \N__23423\,
            I => \N__23418\
        );

    \I__4403\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23413\
        );

    \I__4402\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23413\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__23418\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__23413\,
            I => \ppm_encoder_1.aileronZ0Z_9\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__23408\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\
        );

    \I__4398\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__4396\ : Span4Mux_s3_v
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__23396\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__23387\,
            I => \ppm_encoder_1.pulses2countZ0Z_9\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__4390\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__4388\ : Span4Mux_v
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__23372\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__23369\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\
        );

    \I__4385\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__23363\,
            I => \N__23358\
        );

    \I__4383\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23353\
        );

    \I__4382\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23353\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__23358\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__23353\,
            I => \ppm_encoder_1.init_pulsesZ0Z_1\
        );

    \I__4379\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__23342\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\
        );

    \I__4376\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23334\
        );

    \I__4375\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23331\
        );

    \I__4374\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23328\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__23334\,
            I => \N__23325\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__23331\,
            I => \N__23322\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__23328\,
            I => \N__23319\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__23325\,
            I => \N__23316\
        );

    \I__4369\ : Span4Mux_s1_v
    port map (
            O => \N__23322\,
            I => \N__23309\
        );

    \I__4368\ : Span4Mux_h
    port map (
            O => \N__23319\,
            I => \N__23309\
        );

    \I__4367\ : Span4Mux_v
    port map (
            O => \N__23316\,
            I => \N__23309\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__23309\,
            I => \ppm_encoder_1.init_pulsesZ0Z_11\
        );

    \I__4365\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__23300\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_11\
        );

    \I__4362\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23289\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__23296\,
            I => \N__23285\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23277\
        );

    \I__4359\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23277\
        );

    \I__4358\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23277\
        );

    \I__4357\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23274\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23271\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23264\
        );

    \I__4354\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23264\
        );

    \I__4353\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23264\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23261\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__23274\,
            I => \N__23254\
        );

    \I__4350\ : Span4Mux_h
    port map (
            O => \N__23271\,
            I => \N__23254\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__23264\,
            I => \N__23254\
        );

    \I__4348\ : Span4Mux_s3_v
    port map (
            O => \N__23261\,
            I => \N__23250\
        );

    \I__4347\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23247\
        );

    \I__4346\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23244\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__23250\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__23247\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__23244\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\
        );

    \I__4342\ : InMux
    port map (
            O => \N__23237\,
            I => \N__23224\
        );

    \I__4341\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23219\
        );

    \I__4340\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23219\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__23234\,
            I => \N__23216\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__23233\,
            I => \N__23213\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__23232\,
            I => \N__23208\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__23231\,
            I => \N__23205\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23202\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__23229\,
            I => \N__23198\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \N__23195\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23188\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23183\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23183\
        );

    \I__4329\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23178\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23178\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23173\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23173\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23168\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23168\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23164\
        );

    \I__4322\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23161\
        );

    \I__4321\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23156\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23156\
        );

    \I__4319\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23151\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23151\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__23192\,
            I => \N__23148\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__23191\,
            I => \N__23145\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23142\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__23183\,
            I => \N__23137\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__23178\,
            I => \N__23137\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23132\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23132\
        );

    \I__4310\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23129\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__23164\,
            I => \N__23122\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23122\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__23156\,
            I => \N__23122\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N__23119\
        );

    \I__4305\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23114\
        );

    \I__4304\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23114\
        );

    \I__4303\ : Span4Mux_s1_v
    port map (
            O => \N__23142\,
            I => \N__23105\
        );

    \I__4302\ : Span4Mux_s1_v
    port map (
            O => \N__23137\,
            I => \N__23105\
        );

    \I__4301\ : Span4Mux_s2_h
    port map (
            O => \N__23132\,
            I => \N__23105\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__23129\,
            I => \N__23105\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__23122\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__4298\ : Odrv4
    port map (
            O => \N__23119\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__23114\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__23105\,
            I => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\
        );

    \I__4295\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__23093\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\
        );

    \I__4293\ : CascadeMux
    port map (
            O => \N__23090\,
            I => \N__23077\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23072\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23069\
        );

    \I__4290\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23064\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23064\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__23085\,
            I => \N__23056\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__23084\,
            I => \N__23052\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \N__23048\
        );

    \I__4285\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23041\
        );

    \I__4284\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23036\
        );

    \I__4283\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23036\
        );

    \I__4282\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23031\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23031\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23026\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23023\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23018\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23018\
        );

    \I__4276\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23011\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23011\
        );

    \I__4274\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23011\
        );

    \I__4273\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23002\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23002\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23002\
        );

    \I__4270\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23002\
        );

    \I__4269\ : InMux
    port map (
            O => \N__23052\,
            I => \N__22997\
        );

    \I__4268\ : InMux
    port map (
            O => \N__23051\,
            I => \N__22997\
        );

    \I__4267\ : InMux
    port map (
            O => \N__23048\,
            I => \N__22994\
        );

    \I__4266\ : InMux
    port map (
            O => \N__23047\,
            I => \N__22989\
        );

    \I__4265\ : InMux
    port map (
            O => \N__23046\,
            I => \N__22989\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__23045\,
            I => \N__22986\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__23044\,
            I => \N__22979\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__23041\,
            I => \N__22971\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__22971\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__22971\
        );

    \I__4259\ : InMux
    port map (
            O => \N__23030\,
            I => \N__22966\
        );

    \I__4258\ : InMux
    port map (
            O => \N__23029\,
            I => \N__22966\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__23026\,
            I => \N__22963\
        );

    \I__4256\ : Span4Mux_v
    port map (
            O => \N__23023\,
            I => \N__22960\
        );

    \I__4255\ : Span4Mux_h
    port map (
            O => \N__23018\,
            I => \N__22951\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__23011\,
            I => \N__22951\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__23002\,
            I => \N__22951\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22951\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__22994\,
            I => \N__22937\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__22989\,
            I => \N__22937\
        );

    \I__4249\ : InMux
    port map (
            O => \N__22986\,
            I => \N__22928\
        );

    \I__4248\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22928\
        );

    \I__4247\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22928\
        );

    \I__4246\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22928\
        );

    \I__4245\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22921\
        );

    \I__4244\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22921\
        );

    \I__4243\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22921\
        );

    \I__4242\ : Span4Mux_s2_v
    port map (
            O => \N__22971\,
            I => \N__22916\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22916\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__22963\,
            I => \N__22909\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__22960\,
            I => \N__22909\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__22951\,
            I => \N__22909\
        );

    \I__4237\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22902\
        );

    \I__4236\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22902\
        );

    \I__4235\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22902\
        );

    \I__4234\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22893\
        );

    \I__4233\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22893\
        );

    \I__4232\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22893\
        );

    \I__4231\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22893\
        );

    \I__4230\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22888\
        );

    \I__4229\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22888\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__22937\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__22928\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__22921\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__22916\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__22909\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__22902\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__22893\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__22888\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\
        );

    \I__4220\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22865\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__22865\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_16\
        );

    \I__4217\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__4215\ : Odrv12
    port map (
            O => \N__22856\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\
        );

    \I__4214\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__22850\,
            I => \ppm_encoder_1.pulses2countZ0Z_10\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22844\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__4210\ : Span4Mux_v
    port map (
            O => \N__22841\,
            I => \N__22838\
        );

    \I__4209\ : Span4Mux_h
    port map (
            O => \N__22838\,
            I => \N__22835\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__22832\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\
        );

    \I__4206\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22826\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__22820\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__4201\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__22811\,
            I => \ppm_encoder_1.pulses2countZ0Z_11\
        );

    \I__4199\ : InMux
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__22799\,
            I => \ppm_encoder_1.N_300\
        );

    \I__4195\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__22793\,
            I => \N__22788\
        );

    \I__4193\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22783\
        );

    \I__4192\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22783\
        );

    \I__4191\ : Odrv12
    port map (
            O => \N__22788\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__22783\,
            I => \ppm_encoder_1.aileronZ0Z_8\
        );

    \I__4189\ : CascadeMux
    port map (
            O => \N__22778\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\
        );

    \I__4188\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__22772\,
            I => \N__22768\
        );

    \I__4186\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22765\
        );

    \I__4185\ : Span4Mux_v
    port map (
            O => \N__22768\,
            I => \N__22759\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22759\
        );

    \I__4183\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22756\
        );

    \I__4182\ : Span4Mux_v
    port map (
            O => \N__22759\,
            I => \N__22753\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__22756\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__22753\,
            I => \ppm_encoder_1.throttleZ0Z_2\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__22748\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__4178\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__22736\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\
        );

    \I__4174\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__22730\,
            I => \ppm_encoder_1.pulses2countZ0Z_8\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__22727\,
            I => \ppm_encoder_1.N_145_17_cascade_\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__22724\,
            I => \N__22721\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__22718\,
            I => \ppm_encoder_1.N_145_17\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__22715\,
            I => \ppm_encoder_1.N_238_cascade_\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22709\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__4164\ : Odrv4
    port map (
            O => \N__22703\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\
        );

    \I__4163\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22697\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\
        );

    \I__4161\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__22691\,
            I => \ppm_encoder_1.pulses2countZ0Z_4\
        );

    \I__4159\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22682\
        );

    \I__4157\ : Odrv12
    port map (
            O => \N__22682\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\
        );

    \I__4156\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__22670\,
            I => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__22661\,
            I => \ppm_encoder_1.pulses2countZ0Z_5\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__22658\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__22655\,
            I => \N__22652\
        );

    \I__4147\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22649\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__22643\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\
        );

    \I__4143\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22636\
        );

    \I__4142\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22633\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__22636\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__22633\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22624\
        );

    \I__4138\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22621\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22618\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22615\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__22618\,
            I => \N__22610\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__22615\,
            I => \N__22610\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__22610\,
            I => \ppm_encoder_1.un1_init_pulses_0_11\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22603\
        );

    \I__4131\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22600\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__22603\,
            I => \N__22596\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22593\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22590\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__22596\,
            I => \N__22585\
        );

    \I__4126\ : Span4Mux_v
    port map (
            O => \N__22593\,
            I => \N__22585\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__22590\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__22585\,
            I => \ppm_encoder_1.throttleZ0Z_10\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__22580\,
            I => \ppm_encoder_1.N_302_cascade_\
        );

    \I__4122\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22571\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22568\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22565\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22562\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22571\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__22568\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__22565\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__22562\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__22550\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__22547\,
            I => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\
        );

    \I__4111\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22539\
        );

    \I__4110\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22534\
        );

    \I__4109\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22534\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__22539\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__22534\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__22529\,
            I => \N__22524\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \N__22521\
        );

    \I__4104\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22516\
        );

    \I__4103\ : InMux
    port map (
            O => \N__22524\,
            I => \N__22516\
        );

    \I__4102\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22513\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__22516\,
            I => \N__22510\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__22513\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__22510\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__22505\,
            I => \N__22501\
        );

    \I__4097\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22497\
        );

    \I__4096\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22494\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22491\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22488\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__22494\,
            I => \N__22485\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22478\
        );

    \I__4091\ : Sp12to4
    port map (
            O => \N__22488\,
            I => \N__22473\
        );

    \I__4090\ : Span12Mux_s4_h
    port map (
            O => \N__22485\,
            I => \N__22473\
        );

    \I__4089\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22468\
        );

    \I__4088\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22468\
        );

    \I__4087\ : InMux
    port map (
            O => \N__22482\,
            I => \N__22465\
        );

    \I__4086\ : InMux
    port map (
            O => \N__22481\,
            I => \N__22462\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__22478\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__4084\ : Odrv12
    port map (
            O => \N__22473\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22468\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__22465\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__22462\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__22451\,
            I => \N__22447\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22443\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22438\
        );

    \I__4077\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22438\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__22443\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22438\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\
        );

    \I__4074\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22429\
        );

    \I__4073\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22426\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__22429\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__22426\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22418\,
            I => \N__22414\
        );

    \I__4068\ : InMux
    port map (
            O => \N__22417\,
            I => \N__22411\
        );

    \I__4067\ : Span4Mux_h
    port map (
            O => \N__22414\,
            I => \N__22408\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22402\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__22408\,
            I => \N__22398\
        );

    \I__4064\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22395\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__22406\,
            I => \N__22392\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__22405\,
            I => \N__22389\
        );

    \I__4061\ : Span12Mux_s6_v
    port map (
            O => \N__22402\,
            I => \N__22386\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22383\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__22398\,
            I => \N__22378\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22378\
        );

    \I__4057\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22375\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22372\
        );

    \I__4055\ : Odrv12
    port map (
            O => \N__22386\,
            I => \ppm_encoder_1.N_227\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__22383\,
            I => \ppm_encoder_1.N_227\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__22378\,
            I => \ppm_encoder_1.N_227\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22375\,
            I => \ppm_encoder_1.N_227\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__22372\,
            I => \ppm_encoder_1.N_227\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__22361\,
            I => \N__22355\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__22360\,
            I => \N__22350\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__22359\,
            I => \N__22347\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \N__22344\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22338\
        );

    \I__4045\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22333\
        );

    \I__4044\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22333\
        );

    \I__4043\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22330\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22327\
        );

    \I__4041\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22324\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22321\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__22342\,
            I => \N__22318\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__22341\,
            I => \N__22315\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__22338\,
            I => \N__22311\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__22333\,
            I => \N__22308\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22305\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__22327\,
            I => \N__22302\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22299\
        );

    \I__4032\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22296\
        );

    \I__4031\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22291\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22315\,
            I => \N__22291\
        );

    \I__4029\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22288\
        );

    \I__4028\ : Span4Mux_s2_h
    port map (
            O => \N__22311\,
            I => \N__22283\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__22308\,
            I => \N__22283\
        );

    \I__4026\ : Span4Mux_s3_h
    port map (
            O => \N__22305\,
            I => \N__22280\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__22302\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__22299\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__22296\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__22291\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__22288\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__22283\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__22280\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__22265\,
            I => \N__22257\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__22264\,
            I => \N__22253\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22246\
        );

    \I__4015\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22243\
        );

    \I__4014\ : InMux
    port map (
            O => \N__22261\,
            I => \N__22240\
        );

    \I__4013\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22237\
        );

    \I__4012\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22228\
        );

    \I__4011\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22228\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22228\
        );

    \I__4009\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22228\
        );

    \I__4008\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22225\
        );

    \I__4007\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22219\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22216\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__22246\,
            I => \N__22209\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__22243\,
            I => \N__22209\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22209\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22206\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22203\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__22225\,
            I => \N__22199\
        );

    \I__3999\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22194\
        );

    \I__3998\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22194\
        );

    \I__3997\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22191\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__22219\,
            I => \N__22188\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22179\
        );

    \I__3994\ : Span4Mux_v
    port map (
            O => \N__22209\,
            I => \N__22179\
        );

    \I__3993\ : Span4Mux_v
    port map (
            O => \N__22206\,
            I => \N__22179\
        );

    \I__3992\ : Span4Mux_s2_h
    port map (
            O => \N__22203\,
            I => \N__22179\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22176\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__22199\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__22194\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__22191\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3987\ : Odrv4
    port map (
            O => \N__22188\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__22179\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__22176\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0\
        );

    \I__3984\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22156\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22159\,
            I => \N__22153\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__22156\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__22153\,
            I => \ppm_encoder_1.un1_init_pulses_0_8\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__22148\,
            I => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__3977\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__22133\,
            I => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__22130\,
            I => \N__22126\
        );

    \I__3972\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22120\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22117\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__22125\,
            I => \N__22114\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__22124\,
            I => \N__22111\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__22123\,
            I => \N__22107\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__22120\,
            I => \N__22102\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__22117\,
            I => \N__22099\
        );

    \I__3965\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22096\
        );

    \I__3964\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22092\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22089\
        );

    \I__3962\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22086\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__22106\,
            I => \N__22083\
        );

    \I__3960\ : CascadeMux
    port map (
            O => \N__22105\,
            I => \N__22079\
        );

    \I__3959\ : Span4Mux_s3_h
    port map (
            O => \N__22102\,
            I => \N__22075\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__22099\,
            I => \N__22070\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22070\
        );

    \I__3956\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22067\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22064\
        );

    \I__3954\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22061\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__22086\,
            I => \N__22058\
        );

    \I__3952\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22055\
        );

    \I__3951\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22048\
        );

    \I__3950\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22048\
        );

    \I__3949\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22048\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__22075\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__22070\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__22067\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__22064\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__22061\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__22058\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__22055\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__22048\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__22031\,
            I => \N__22027\
        );

    \I__3939\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22023\
        );

    \I__3938\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22020\
        );

    \I__3937\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22017\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22013\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__22020\,
            I => \N__22010\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__22017\,
            I => \N__22007\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__22016\,
            I => \N__22003\
        );

    \I__3932\ : Span4Mux_s3_h
    port map (
            O => \N__22013\,
            I => \N__21993\
        );

    \I__3931\ : Span4Mux_s3_h
    port map (
            O => \N__22010\,
            I => \N__21990\
        );

    \I__3930\ : Span4Mux_s3_h
    port map (
            O => \N__22007\,
            I => \N__21987\
        );

    \I__3929\ : InMux
    port map (
            O => \N__22006\,
            I => \N__21984\
        );

    \I__3928\ : InMux
    port map (
            O => \N__22003\,
            I => \N__21979\
        );

    \I__3927\ : InMux
    port map (
            O => \N__22002\,
            I => \N__21979\
        );

    \I__3926\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21976\
        );

    \I__3925\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21973\
        );

    \I__3924\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21970\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21963\
        );

    \I__3922\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21963\
        );

    \I__3921\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21963\
        );

    \I__3920\ : Odrv4
    port map (
            O => \N__21993\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__21990\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__21987\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__21984\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__21979\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__21976\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__21973\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__21970\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__21963\,
            I => \ppm_encoder_1.init_pulses_2_sqmuxa_0\
        );

    \I__3911\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__21941\,
            I => \ppm_encoder_1.un2_throttle_iv_1_8\
        );

    \I__3909\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21929\
        );

    \I__3908\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21929\
        );

    \I__3907\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21929\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__21929\,
            I => \ppm_encoder_1.elevatorZ0Z_8\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__3904\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21919\
        );

    \I__3903\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__21916\,
            I => \N__21910\
        );

    \I__3900\ : Span4Mux_h
    port map (
            O => \N__21913\,
            I => \N__21904\
        );

    \I__3899\ : Span4Mux_s3_h
    port map (
            O => \N__21910\,
            I => \N__21904\
        );

    \I__3898\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21901\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__21904\,
            I => \N__21898\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__21901\,
            I => throttle_command_8
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__21898\,
            I => throttle_command_8
        );

    \I__3894\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__21887\,
            I => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\
        );

    \I__3891\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21875\
        );

    \I__3890\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21875\
        );

    \I__3889\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21875\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__21875\,
            I => \ppm_encoder_1.throttleZ0Z_8\
        );

    \I__3887\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21868\
        );

    \I__3886\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21865\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21860\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21860\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__21857\,
            I => scaler_2_data_8
        );

    \I__3881\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__21848\,
            I => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\
        );

    \I__3878\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21840\
        );

    \I__3877\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21837\
        );

    \I__3876\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21834\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21829\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__21837\,
            I => \N__21829\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__21834\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__21829\,
            I => \ppm_encoder_1.throttleZ0Z_4\
        );

    \I__3871\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__21818\,
            I => \ppm_encoder_1.N_296\
        );

    \I__3868\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21808\
        );

    \I__3866\ : InMux
    port map (
            O => \N__21811\,
            I => \N__21805\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__21808\,
            I => throttle_command_4
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__21805\,
            I => throttle_command_4
        );

    \I__3863\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__21791\,
            I => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__21782\,
            I => \N__21778\
        );

    \I__3856\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21775\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__21778\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__21775\,
            I => \ppm_encoder_1.un1_init_pulses_0_12\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__21770\,
            I => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__3851\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__3849\ : Span4Mux_v
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__21755\,
            I => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\
        );

    \I__3847\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__21749\,
            I => \ppm_encoder_1.un2_throttle_iv_1_12\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \ppm_encoder_1.N_304_cascade_\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__21743\,
            I => \N__21739\
        );

    \I__3843\ : InMux
    port map (
            O => \N__21742\,
            I => \N__21736\
        );

    \I__3842\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21733\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21730\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__21733\,
            I => \N__21727\
        );

    \I__3839\ : Span4Mux_v
    port map (
            O => \N__21730\,
            I => \N__21724\
        );

    \I__3838\ : Odrv12
    port map (
            O => \N__21727\,
            I => scaler_2_data_12
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__21724\,
            I => scaler_2_data_12
        );

    \I__3836\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21713\
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__21713\,
            I => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\
        );

    \I__3833\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21701\
        );

    \I__3832\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21701\
        );

    \I__3831\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21701\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__21701\,
            I => \ppm_encoder_1.aileronZ0Z_12\
        );

    \I__3829\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21689\
        );

    \I__3828\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21689\
        );

    \I__3827\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21689\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__21689\,
            I => \ppm_encoder_1.elevatorZ0Z_12\
        );

    \I__3825\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21682\
        );

    \I__3824\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21679\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21676\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21673\
        );

    \I__3821\ : Span4Mux_h
    port map (
            O => \N__21676\,
            I => \N__21670\
        );

    \I__3820\ : Span4Mux_s2_h
    port map (
            O => \N__21673\,
            I => \N__21667\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__21670\,
            I => throttle_command_12
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__21667\,
            I => throttle_command_12
        );

    \I__3817\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__21653\,
            I => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\
        );

    \I__3813\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21641\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21641\
        );

    \I__3811\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21641\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__21641\,
            I => \ppm_encoder_1.throttleZ0Z_12\
        );

    \I__3809\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21614\
        );

    \I__3808\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21614\
        );

    \I__3807\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21614\
        );

    \I__3806\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21614\
        );

    \I__3805\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21611\
        );

    \I__3804\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21608\
        );

    \I__3803\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21605\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21592\
        );

    \I__3801\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21592\
        );

    \I__3800\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21592\
        );

    \I__3799\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21592\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21592\
        );

    \I__3797\ : InMux
    port map (
            O => \N__21626\,
            I => \N__21592\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21589\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21586\
        );

    \I__3794\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21583\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21566\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__21611\,
            I => \N__21563\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21560\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__21605\,
            I => \N__21557\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21554\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21551\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__21586\,
            I => \N__21548\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21545\
        );

    \I__3785\ : SRMux
    port map (
            O => \N__21582\,
            I => \N__21500\
        );

    \I__3784\ : SRMux
    port map (
            O => \N__21581\,
            I => \N__21500\
        );

    \I__3783\ : SRMux
    port map (
            O => \N__21580\,
            I => \N__21500\
        );

    \I__3782\ : SRMux
    port map (
            O => \N__21579\,
            I => \N__21500\
        );

    \I__3781\ : SRMux
    port map (
            O => \N__21578\,
            I => \N__21500\
        );

    \I__3780\ : SRMux
    port map (
            O => \N__21577\,
            I => \N__21500\
        );

    \I__3779\ : SRMux
    port map (
            O => \N__21576\,
            I => \N__21500\
        );

    \I__3778\ : SRMux
    port map (
            O => \N__21575\,
            I => \N__21500\
        );

    \I__3777\ : SRMux
    port map (
            O => \N__21574\,
            I => \N__21500\
        );

    \I__3776\ : SRMux
    port map (
            O => \N__21573\,
            I => \N__21500\
        );

    \I__3775\ : SRMux
    port map (
            O => \N__21572\,
            I => \N__21500\
        );

    \I__3774\ : SRMux
    port map (
            O => \N__21571\,
            I => \N__21500\
        );

    \I__3773\ : SRMux
    port map (
            O => \N__21570\,
            I => \N__21500\
        );

    \I__3772\ : SRMux
    port map (
            O => \N__21569\,
            I => \N__21500\
        );

    \I__3771\ : Glb2LocalMux
    port map (
            O => \N__21566\,
            I => \N__21500\
        );

    \I__3770\ : Glb2LocalMux
    port map (
            O => \N__21563\,
            I => \N__21500\
        );

    \I__3769\ : Glb2LocalMux
    port map (
            O => \N__21560\,
            I => \N__21500\
        );

    \I__3768\ : Glb2LocalMux
    port map (
            O => \N__21557\,
            I => \N__21500\
        );

    \I__3767\ : Glb2LocalMux
    port map (
            O => \N__21554\,
            I => \N__21500\
        );

    \I__3766\ : Glb2LocalMux
    port map (
            O => \N__21551\,
            I => \N__21500\
        );

    \I__3765\ : Glb2LocalMux
    port map (
            O => \N__21548\,
            I => \N__21500\
        );

    \I__3764\ : Glb2LocalMux
    port map (
            O => \N__21545\,
            I => \N__21500\
        );

    \I__3763\ : GlobalMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__3762\ : gio2CtrlBuf
    port map (
            O => \N__21497\,
            I => \N_423_g\
        );

    \I__3761\ : IoInMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__3759\ : Span12Mux_s11_v
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__3758\ : Odrv12
    port map (
            O => \N__21485\,
            I => \pid_alt.N_422_0\
        );

    \I__3757\ : CEMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__21479\,
            I => \pid_alt.state_1_0_0\
        );

    \I__3755\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21472\
        );

    \I__3754\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21465\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__21469\,
            I => \N__21462\
        );

    \I__3751\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21459\
        );

    \I__3750\ : Span12Mux_s4_h
    port map (
            O => \N__21465\,
            I => \N__21456\
        );

    \I__3749\ : Span4Mux_h
    port map (
            O => \N__21462\,
            I => \N__21453\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__21459\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3747\ : Odrv12
    port map (
            O => \N__21456\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__21453\,
            I => \ppm_encoder_1.rudderZ0Z_11\
        );

    \I__3745\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21442\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__21445\,
            I => \N__21439\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__21442\,
            I => \N__21436\
        );

    \I__3742\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21433\
        );

    \I__3741\ : Span4Mux_v
    port map (
            O => \N__21436\,
            I => \N__21427\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21427\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21424\
        );

    \I__3738\ : Span4Mux_v
    port map (
            O => \N__21427\,
            I => \N__21421\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__21424\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__21421\,
            I => \ppm_encoder_1.rudderZ0Z_7\
        );

    \I__3735\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21412\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__21415\,
            I => \N__21408\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21405\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21402\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21399\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__21405\,
            I => \N__21396\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21393\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__21399\,
            I => throttle_command_10
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__21396\,
            I => throttle_command_10
        );

    \I__3726\ : Odrv12
    port map (
            O => \N__21393\,
            I => throttle_command_10
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__21386\,
            I => \N__21383\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21380\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21377\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__21377\,
            I => \N__21374\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__21374\,
            I => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\
        );

    \I__3720\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21367\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21364\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21361\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21358\
        );

    \I__3716\ : Span4Mux_v
    port map (
            O => \N__21361\,
            I => \N__21353\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__21358\,
            I => \N__21353\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__21353\,
            I => throttle_command_13
        );

    \I__3713\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21347\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21347\,
            I => \N__21344\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__21344\,
            I => \N__21341\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__21341\,
            I => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__3707\ : Span4Mux_h
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__21329\,
            I => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21326\,
            I => \N__21323\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21319\
        );

    \I__3703\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21316\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21313\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21310\
        );

    \I__3700\ : Span4Mux_v
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__3699\ : Span4Mux_s3_h
    port map (
            O => \N__21310\,
            I => \N__21304\
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__21307\,
            I => throttle_command_2
        );

    \I__3697\ : Odrv4
    port map (
            O => \N__21304\,
            I => throttle_command_2
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__21299\,
            I => \N__21296\
        );

    \I__3695\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21290\
        );

    \I__3694\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21290\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21287\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__21287\,
            I => \N__21284\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__21284\,
            I => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21281\,
            I => \scaler_2.un2_source_data_0_cry_5\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21269\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21269\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__21263\,
            I => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__3682\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21253\
        );

    \I__3681\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21250\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21247\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21244\
        );

    \I__3678\ : Span12Mux_s4_h
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__3677\ : Span4Mux_v
    port map (
            O => \N__21244\,
            I => \N__21238\
        );

    \I__3676\ : Odrv12
    port map (
            O => \N__21241\,
            I => scaler_2_data_11
        );

    \I__3675\ : Odrv4
    port map (
            O => \N__21238\,
            I => scaler_2_data_11
        );

    \I__3674\ : InMux
    port map (
            O => \N__21233\,
            I => \scaler_2.un2_source_data_0_cry_6\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__3672\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21221\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21221\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__21215\,
            I => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21212\,
            I => \scaler_2.un2_source_data_0_cry_7\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21205\
        );

    \I__3665\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21202\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21205\,
            I => \N__21199\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21196\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__21199\,
            I => \N__21193\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__21196\,
            I => \N__21190\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__21193\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__3659\ : Odrv4
    port map (
            O => \N__21190\,
            I => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\
        );

    \I__3658\ : CascadeMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__3657\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21176\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__21173\,
            I => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21170\,
            I => \bfn_4_17_0_\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21167\,
            I => \scaler_2.un2_source_data_0_cry_9\
        );

    \I__3651\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__3649\ : Span4Mux_h
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__3648\ : Span4Mux_v
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__21152\,
            I => scaler_2_data_14
        );

    \I__3646\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__3644\ : Span12Mux_v
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__3643\ : Odrv12
    port map (
            O => \N__21140\,
            I => alt_ki_7
        );

    \I__3642\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__21131\,
            I => \N__21127\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21124\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__21127\,
            I => \pid_alt.un1_pid_prereg_0_axb_1\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__21124\,
            I => \pid_alt.un1_pid_prereg_0_axb_1\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__3635\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__21107\,
            I => \pid_alt.un1_pid_prereg_0_cry_0_THRU_CO\
        );

    \I__3631\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__3629\ : Span4Mux_h
    port map (
            O => \N__21098\,
            I => \N__21093\
        );

    \I__3628\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21090\
        );

    \I__3627\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21087\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__21093\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__21090\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__21087\,
            I => \pid_alt.pid_preregZ0Z_1\
        );

    \I__3623\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__21074\,
            I => \scaler_2.N_881_i_l_ofxZ0\
        );

    \I__3620\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21065\
        );

    \I__3619\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21065\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__21065\,
            I => \frame_decoder_CH2data_7\
        );

    \I__3617\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21059\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__21056\,
            I => \N__21053\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__21053\,
            I => \scaler_2.un3_source_data_0_axb_7\
        );

    \I__3613\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__21047\,
            I => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__21044\,
            I => \N__21038\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__21043\,
            I => \N__21035\
        );

    \I__3609\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21032\
        );

    \I__3608\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21029\
        );

    \I__3607\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21026\
        );

    \I__3606\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21023\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__21020\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21017\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21012\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__21023\,
            I => \N__21012\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__21020\,
            I => \N__21009\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__21017\,
            I => \N__21004\
        );

    \I__3599\ : Span4Mux_h
    port map (
            O => \N__21012\,
            I => \N__21004\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__21009\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__21004\,
            I => \scaler_2.un2_source_data_0\
        );

    \I__3596\ : InMux
    port map (
            O => \N__20999\,
            I => \scaler_2.un2_source_data_0_cry_1\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__3594\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20987\
        );

    \I__3593\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20987\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__20981\,
            I => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\
        );

    \I__3589\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20971\
        );

    \I__3587\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20968\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__20971\,
            I => \N__20963\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__20968\,
            I => \N__20963\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__20960\,
            I => scaler_2_data_7
        );

    \I__3582\ : InMux
    port map (
            O => \N__20957\,
            I => \scaler_2.un2_source_data_0_cry_2\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__3580\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20945\
        );

    \I__3579\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20945\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__20939\,
            I => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\
        );

    \I__3575\ : InMux
    port map (
            O => \N__20936\,
            I => \scaler_2.un2_source_data_0_cry_3\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__3573\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20924\
        );

    \I__3572\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20924\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__20918\,
            I => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\
        );

    \I__3568\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20912\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__20909\,
            I => \N__20905\
        );

    \I__3565\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20902\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__20905\,
            I => \N__20899\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__20902\,
            I => \N__20896\
        );

    \I__3562\ : Span4Mux_v
    port map (
            O => \N__20899\,
            I => \N__20893\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__20893\,
            I => scaler_2_data_9
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__20890\,
            I => scaler_2_data_9
        );

    \I__3558\ : InMux
    port map (
            O => \N__20885\,
            I => \scaler_2.un2_source_data_0_cry_4\
        );

    \I__3557\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20878\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__20881\,
            I => \N__20875\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__20878\,
            I => \N__20870\
        );

    \I__3554\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20867\
        );

    \I__3553\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20862\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20862\
        );

    \I__3551\ : Span4Mux_v
    port map (
            O => \N__20870\,
            I => \N__20856\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20856\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20853\
        );

    \I__3548\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20850\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__20856\,
            I => \N__20847\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__20853\,
            I => \N__20841\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20838\
        );

    \I__3544\ : Sp12to4
    port map (
            O => \N__20847\,
            I => \N__20835\
        );

    \I__3543\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20828\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20828\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20844\,
            I => \N__20828\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__20841\,
            I => \N__20825\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__20838\,
            I => \N__20822\
        );

    \I__3538\ : Span12Mux_s1_h
    port map (
            O => \N__20835\,
            I => \N__20817\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__20828\,
            I => \N__20817\
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__20825\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__20822\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__20817\,
            I => \pid_alt.error_i_regZ0Z_20\
        );

    \I__3533\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__3530\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20796\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__20800\,
            I => \N__20793\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__20799\,
            I => \N__20790\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20785\
        );

    \I__3526\ : Sp12to4
    port map (
            O => \N__20793\,
            I => \N__20782\
        );

    \I__3525\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20775\
        );

    \I__3524\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20775\
        );

    \I__3523\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20775\
        );

    \I__3522\ : Span4Mux_v
    port map (
            O => \N__20785\,
            I => \N__20772\
        );

    \I__3521\ : Span12Mux_h
    port map (
            O => \N__20782\,
            I => \N__20767\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__20775\,
            I => \N__20767\
        );

    \I__3519\ : Span4Mux_h
    port map (
            O => \N__20772\,
            I => \N__20764\
        );

    \I__3518\ : Span12Mux_v
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__20764\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3516\ : Odrv12
    port map (
            O => \N__20761\,
            I => \pid_alt.error_p_regZ0Z_20\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__20756\,
            I => \N__20753\
        );

    \I__3514\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__20750\,
            I => \N__20747\
        );

    \I__3512\ : Span4Mux_h
    port map (
            O => \N__20747\,
            I => \N__20744\
        );

    \I__3511\ : Sp12to4
    port map (
            O => \N__20744\,
            I => \N__20741\
        );

    \I__3510\ : Odrv12
    port map (
            O => \N__20741\,
            I => \pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20\
        );

    \I__3509\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__20732\,
            I => \frame_decoder_CH2data_1\
        );

    \I__3506\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__20723\,
            I => \frame_decoder_CH2data_2\
        );

    \I__3503\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__20714\,
            I => \frame_decoder_CH2data_3\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__20711\,
            I => \N__20708\
        );

    \I__3499\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__20702\,
            I => \frame_decoder_CH2data_4\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__3495\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__3493\ : Odrv4
    port map (
            O => \N__20690\,
            I => \frame_decoder_CH2data_5\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__3491\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__20678\,
            I => \frame_decoder_CH2data_6\
        );

    \I__3488\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__20672\,
            I => \dron_frame_decoder_1.drone_altitude_11\
        );

    \I__3486\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__20666\,
            I => \dron_frame_decoder_1.drone_altitude_9\
        );

    \I__3484\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__20660\,
            I => \dron_frame_decoder_1.drone_altitude_10\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__20654\,
            I => \dron_frame_decoder_1.drone_altitude_8\
        );

    \I__3480\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__20648\,
            I => drone_altitude_14
        );

    \I__3478\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__20642\,
            I => drone_altitude_2
        );

    \I__3476\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__20636\,
            I => drone_altitude_3
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__3473\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20626\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20623\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20626\,
            I => \N__20615\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__20623\,
            I => \N__20615\
        );

    \I__3469\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20612\
        );

    \I__3468\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20607\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20607\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__20615\,
            I => \N__20604\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20601\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20598\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__20604\,
            I => \N__20595\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20590\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__20598\,
            I => \N__20590\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__20595\,
            I => \pid_alt.error_i_regZ0Z_18\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__20590\,
            I => \pid_alt.error_i_regZ0Z_18\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__3457\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20576\
        );

    \I__3456\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20576\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20573\
        );

    \I__3454\ : Span4Mux_h
    port map (
            O => \N__20573\,
            I => \N__20569\
        );

    \I__3453\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20566\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__20569\,
            I => \N__20561\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20561\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__20561\,
            I => \N__20558\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__20558\,
            I => \N__20555\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__20555\,
            I => \pid_alt.error_p_regZ0Z_18\
        );

    \I__3447\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20546\
        );

    \I__3445\ : Span4Mux_h
    port map (
            O => \N__20546\,
            I => \N__20543\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__20543\,
            I => \N__20540\
        );

    \I__3443\ : Odrv4
    port map (
            O => \N__20540\,
            I => \pid_alt.error_p_reg_esr_RNIF43KZ0Z_18\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20530\
        );

    \I__3440\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20525\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__20530\,
            I => \N__20522\
        );

    \I__3438\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20519\
        );

    \I__3437\ : InMux
    port map (
            O => \N__20528\,
            I => \N__20516\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__20525\,
            I => \N__20513\
        );

    \I__3435\ : Span4Mux_s1_v
    port map (
            O => \N__20522\,
            I => \N__20508\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20508\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__20516\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__20513\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__20508\,
            I => \ppm_encoder_1.init_pulsesZ0Z_2\
        );

    \I__3430\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20498\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__3428\ : Span4Mux_h
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__20492\,
            I => alt_kp_7
        );

    \I__3426\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20486\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20482\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__3423\ : Span4Mux_h
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__20479\,
            I => alt_kp_4
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__20476\,
            I => alt_kp_4
        );

    \I__3420\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__3418\ : Span4Mux_h
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__20462\,
            I => \pid_alt.O_10\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20455\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20446\
        );

    \I__3412\ : Span4Mux_v
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__3411\ : Span12Mux_v
    port map (
            O => \N__20446\,
            I => \N__20440\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__20443\,
            I => \pid_alt.error_p_regZ0Z_6\
        );

    \I__3409\ : Odrv12
    port map (
            O => \N__20440\,
            I => \pid_alt.error_p_regZ0Z_6\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__20435\,
            I => \N__20431\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20428\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20425\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20422\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20425\,
            I => \N__20418\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__20422\,
            I => \N__20415\
        );

    \I__3402\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20412\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__20418\,
            I => \N__20409\
        );

    \I__3400\ : Span4Mux_v
    port map (
            O => \N__20415\,
            I => \N__20406\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__20412\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__20409\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__20406\,
            I => \pid_alt.error_i_regZ0Z_6\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20399\,
            I => \N__20394\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20391\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20387\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20394\,
            I => \N__20384\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20381\
        );

    \I__3391\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20378\
        );

    \I__3390\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20375\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__20384\,
            I => \N__20372\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__20381\,
            I => \N__20367\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20367\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20375\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__20372\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__20367\,
            I => \pid_alt.error_i_acummZ0Z_6\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__3379\ : Sp12to4
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__3378\ : Odrv12
    port map (
            O => \N__20345\,
            I => \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6\
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_\
        );

    \I__3376\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20333\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__20327\,
            I => \pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7\
        );

    \I__3371\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20321\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__20321\,
            I => \N__20318\
        );

    \I__3369\ : Span4Mux_h
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__20315\,
            I => \pid_alt.O_11\
        );

    \I__3367\ : CEMux
    port map (
            O => \N__20312\,
            I => \N__20270\
        );

    \I__3366\ : CEMux
    port map (
            O => \N__20311\,
            I => \N__20270\
        );

    \I__3365\ : CEMux
    port map (
            O => \N__20310\,
            I => \N__20270\
        );

    \I__3364\ : CEMux
    port map (
            O => \N__20309\,
            I => \N__20270\
        );

    \I__3363\ : CEMux
    port map (
            O => \N__20308\,
            I => \N__20270\
        );

    \I__3362\ : CEMux
    port map (
            O => \N__20307\,
            I => \N__20270\
        );

    \I__3361\ : CEMux
    port map (
            O => \N__20306\,
            I => \N__20270\
        );

    \I__3360\ : CEMux
    port map (
            O => \N__20305\,
            I => \N__20270\
        );

    \I__3359\ : CEMux
    port map (
            O => \N__20304\,
            I => \N__20270\
        );

    \I__3358\ : CEMux
    port map (
            O => \N__20303\,
            I => \N__20270\
        );

    \I__3357\ : CEMux
    port map (
            O => \N__20302\,
            I => \N__20270\
        );

    \I__3356\ : CEMux
    port map (
            O => \N__20301\,
            I => \N__20270\
        );

    \I__3355\ : CEMux
    port map (
            O => \N__20300\,
            I => \N__20270\
        );

    \I__3354\ : CEMux
    port map (
            O => \N__20299\,
            I => \N__20270\
        );

    \I__3353\ : GlobalMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__3352\ : gio2CtrlBuf
    port map (
            O => \N__20267\,
            I => \pid_alt.N_422_0_g\
        );

    \I__3351\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20258\
        );

    \I__3350\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20258\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__3348\ : Span4Mux_v
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__20252\,
            I => \pid_alt.error_p_regZ0Z_7\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__3345\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__3343\ : Span4Mux_h
    port map (
            O => \N__20240\,
            I => \N__20235\
        );

    \I__3342\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20230\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20230\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__20235\,
            I => \pid_alt.error_i_regZ0Z_7\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__20230\,
            I => \pid_alt.error_i_regZ0Z_7\
        );

    \I__3338\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20217\
        );

    \I__3337\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20217\
        );

    \I__3336\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20214\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__20222\,
            I => \N__20211\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__20217\,
            I => \N__20208\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20205\
        );

    \I__3332\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20202\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__20208\,
            I => \N__20197\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__20205\,
            I => \N__20197\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__20202\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__20197\,
            I => \pid_alt.error_i_acummZ0Z_7\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__20192\,
            I => \N__20188\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \N__20185\
        );

    \I__3325\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20182\
        );

    \I__3324\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20179\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20176\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__20179\,
            I => \N__20171\
        );

    \I__3321\ : Span12Mux_v
    port map (
            O => \N__20176\,
            I => \N__20171\
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__20171\,
            I => \pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20161\
        );

    \I__3317\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20158\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20155\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__20158\,
            I => \N__20152\
        );

    \I__3314\ : Span4Mux_s3_h
    port map (
            O => \N__20155\,
            I => \N__20149\
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__20152\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__20149\,
            I => \ppm_encoder_1.un1_init_pulses_0_4\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__20141\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_4\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20129\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20129\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20129\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__20129\,
            I => \ppm_encoder_1.init_pulsesZ0Z_4\
        );

    \I__3305\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20114\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20114\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20114\
        );

    \I__3302\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20109\
        );

    \I__3301\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20109\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20102\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__20114\,
            I => \N__20095\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__20109\,
            I => \N__20095\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20092\
        );

    \I__3296\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20085\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20085\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20085\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20079\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20074\
        );

    \I__3291\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20074\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__20095\,
            I => \N__20068\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__20092\,
            I => \N__20065\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__20085\,
            I => \N__20062\
        );

    \I__3287\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20059\
        );

    \I__3286\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20054\
        );

    \I__3285\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20054\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__20079\,
            I => \N__20049\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__20074\,
            I => \N__20049\
        );

    \I__3282\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20042\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20042\
        );

    \I__3280\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20042\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__20068\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__20065\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3277\ : Odrv12
    port map (
            O => \N__20062\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__20059\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__20054\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__20049\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__20042\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1\
        );

    \I__3272\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__20024\,
            I => \ppm_encoder_1.un1_init_pulses_11_5\
        );

    \I__3270\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__3268\ : Span4Mux_s2_v
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__20012\,
            I => \ppm_encoder_1.un1_init_pulses_10_5\
        );

    \I__3266\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20000\
        );

    \I__3265\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20000\
        );

    \I__3264\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20000\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__19994\,
            I => \ppm_encoder_1.init_pulsesZ0Z_5\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__3259\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__19985\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_14\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__19982\,
            I => \ppm_encoder_1.N_319_cascade_\
        );

    \I__3256\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__19976\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_12\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__3253\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__19967\,
            I => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__3250\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__19955\,
            I => \ppm_encoder_1.un1_init_pulses_10_2\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__19949\,
            I => \ppm_encoder_1.un1_init_pulses_11_2\
        );

    \I__3245\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19942\
        );

    \I__3244\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19939\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19930\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19930\
        );

    \I__3241\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19923\
        );

    \I__3240\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19923\
        );

    \I__3239\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19923\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__19935\,
            I => \N__19918\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__19930\,
            I => \N__19914\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19911\
        );

    \I__3235\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19906\
        );

    \I__3234\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19906\
        );

    \I__3233\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19901\
        );

    \I__3232\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19901\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__19914\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__19911\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__19906\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19901\,
            I => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__3226\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__19886\,
            I => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__19883\,
            I => \N__19880\
        );

    \I__3223\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__19871\,
            I => \ppm_encoder_1.un1_init_pulses_10_6\
        );

    \I__3219\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__19865\,
            I => \ppm_encoder_1.un1_init_pulses_11_6\
        );

    \I__3217\ : InMux
    port map (
            O => \N__19862\,
            I => \N__19858\
        );

    \I__3216\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19855\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19852\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__19855\,
            I => \N__19849\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__19849\,
            I => \N__19843\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__19846\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__19843\,
            I => \ppm_encoder_1.un1_init_pulses_0_6\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__19838\,
            I => \N__19834\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \N__19830\
        );

    \I__3207\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19825\
        );

    \I__3206\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19825\
        );

    \I__3205\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19822\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19817\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__19822\,
            I => \N__19817\
        );

    \I__3202\ : Span4Mux_s3_h
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__19814\,
            I => \ppm_encoder_1.un1_init_pulses_0\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__3199\ : InMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__19802\,
            I => \ppm_encoder_1.un1_init_pulses_10_16\
        );

    \I__3196\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__19796\,
            I => \ppm_encoder_1.un1_init_pulses_11_16\
        );

    \I__3194\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__19790\,
            I => \ppm_encoder_1.un1_init_pulses_11_4\
        );

    \I__3192\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__3190\ : Span4Mux_s2_v
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__19778\,
            I => \ppm_encoder_1.un1_init_pulses_10_4\
        );

    \I__3188\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19771\
        );

    \I__3187\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19768\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19765\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__19768\,
            I => \N__19762\
        );

    \I__3184\ : Odrv12
    port map (
            O => \N__19765\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__19762\,
            I => \ppm_encoder_1.aileronZ0Z_4\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__19754\,
            I => \ppm_encoder_1.un1_init_pulses_11_3\
        );

    \I__3180\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__19745\,
            I => \ppm_encoder_1.un1_init_pulses_10_3\
        );

    \I__3177\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__19739\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_3\
        );

    \I__3175\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19733\,
            I => \ppm_encoder_1.un1_init_pulses_11_7\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__19721\,
            I => \ppm_encoder_1.un1_init_pulses_10_7\
        );

    \I__3169\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__19715\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_7\
        );

    \I__3167\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__19709\,
            I => \N__19705\
        );

    \I__3165\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19702\
        );

    \I__3164\ : Span4Mux_s3_h
    port map (
            O => \N__19705\,
            I => \N__19697\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19697\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__19697\,
            I => \ppm_encoder_1.un1_init_pulses_0_7\
        );

    \I__3161\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19685\
        );

    \I__3160\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19685\
        );

    \I__3159\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19685\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__19685\,
            I => \ppm_encoder_1.init_pulsesZ0Z_7\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19676\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__19676\,
            I => \ppm_encoder_1.un1_init_pulses_11_8\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__3153\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__19667\,
            I => \ppm_encoder_1.un1_init_pulses_10_8\
        );

    \I__3151\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__3149\ : Span4Mux_s3_h
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__19655\,
            I => \ppm_encoder_1.un1_init_pulses_11_0\
        );

    \I__3147\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19648\
        );

    \I__3146\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19645\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__19648\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__19645\,
            I => \ppm_encoder_1.un1_init_pulses_0_3\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__3142\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__19634\,
            I => \ppm_encoder_1.throttle_RNI82223Z0Z_3\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__3138\ : Span4Mux_h
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__19622\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__19619\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__3133\ : Span4Mux_v
    port map (
            O => \N__19610\,
            I => \N__19606\
        );

    \I__3132\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19603\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__19606\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__19603\,
            I => \ppm_encoder_1.un1_init_pulses_0_10\
        );

    \I__3129\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19593\
        );

    \I__3128\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19588\
        );

    \I__3127\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19588\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__19593\,
            I => \N__19585\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19588\,
            I => \N__19580\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__19585\,
            I => \N__19580\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__19580\,
            I => \ppm_encoder_1.init_pulsesZ0Z_9\
        );

    \I__3122\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19573\
        );

    \I__3121\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19570\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__19573\,
            I => \N__19565\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__19570\,
            I => \N__19565\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__19565\,
            I => \ppm_encoder_1.un1_init_pulses_0_9\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__3114\ : Span4Mux_s3_h
    port map (
            O => \N__19553\,
            I => \N__19549\
        );

    \I__3113\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19546\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__19549\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__19546\,
            I => \ppm_encoder_1.un1_init_pulses_0_2\
        );

    \I__3110\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19538\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__3108\ : Span4Mux_h
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__19532\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_10\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__19529\,
            I => \ppm_encoder_1.un2_throttle_iv_1_4_cascade_\
        );

    \I__3105\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__19523\,
            I => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__19517\,
            I => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__19511\,
            I => \ppm_encoder_1.un2_throttle_iv_0_4\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__19508\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__19505\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__3096\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__19496\,
            I => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__19493\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\
        );

    \I__3093\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19485\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19482\
        );

    \I__3091\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19477\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__19485\,
            I => \N__19472\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__19482\,
            I => \N__19472\
        );

    \I__3088\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19469\
        );

    \I__3087\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19466\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19463\
        );

    \I__3085\ : Span4Mux_v
    port map (
            O => \N__19472\,
            I => \N__19456\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19456\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19456\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__19463\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__19456\,
            I => \pid_alt.pid_preregZ0Z_4\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__19451\,
            I => \pid_alt.N_88_cascade_\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19442\
        );

    \I__3078\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19442\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19438\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__19438\,
            I => \pid_alt.N_90\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__19435\,
            I => \pid_alt.N_90\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__19430\,
            I => \N__19427\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19420\
        );

    \I__3071\ : InMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__19425\,
            I => \N__19416\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__19420\,
            I => \N__19410\
        );

    \I__3068\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19403\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19403\
        );

    \I__3066\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19403\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__19414\,
            I => \N__19399\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__19413\,
            I => \N__19395\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__19410\,
            I => \N__19391\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19388\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19381\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19381\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19381\
        );

    \I__3058\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19378\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19375\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__19391\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__19388\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__19381\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__19378\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__19375\,
            I => \pid_alt.pid_preregZ0Z_22\
        );

    \I__3051\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__19357\,
            I => \N__19349\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19354\,
            I => \N__19349\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__19349\,
            I => \pid_alt.pid_preregZ0Z_2\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__19346\,
            I => \pid_alt.N_90_cascade_\
        );

    \I__3044\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19337\
        );

    \I__3043\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19337\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19327\
        );

    \I__3041\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19324\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19319\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19310\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19310\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19310\
        );

    \I__3036\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19310\
        );

    \I__3035\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19307\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__19327\,
            I => \N__19302\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19324\,
            I => \N__19302\
        );

    \I__3032\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19297\
        );

    \I__3031\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19297\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__19319\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19310\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__19307\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__19302\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__19297\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\
        );

    \I__3025\ : CEMux
    port map (
            O => \N__19286\,
            I => \N__19281\
        );

    \I__3024\ : CEMux
    port map (
            O => \N__19285\,
            I => \N__19278\
        );

    \I__3023\ : CEMux
    port map (
            O => \N__19284\,
            I => \N__19275\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19281\,
            I => \N__19270\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19270\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19265\
        );

    \I__3019\ : Span4Mux_v
    port map (
            O => \N__19270\,
            I => \N__19265\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__19265\,
            I => \pid_alt.N_60_i_1\
        );

    \I__3017\ : SRMux
    port map (
            O => \N__19262\,
            I => \N__19257\
        );

    \I__3016\ : SRMux
    port map (
            O => \N__19261\,
            I => \N__19253\
        );

    \I__3015\ : SRMux
    port map (
            O => \N__19260\,
            I => \N__19250\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19246\
        );

    \I__3013\ : SRMux
    port map (
            O => \N__19256\,
            I => \N__19243\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19240\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19237\
        );

    \I__3010\ : SRMux
    port map (
            O => \N__19249\,
            I => \N__19234\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__19246\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__19243\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__3007\ : Odrv12
    port map (
            O => \N__19240\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__3006\ : Odrv12
    port map (
            O => \N__19237\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__19234\,
            I => \pid_alt.un1_reset_0_i\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19219\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19216\
        );

    \I__3002\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19213\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__19216\,
            I => \N__19210\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__19213\,
            I => \N__19207\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__19210\,
            I => \N__19204\
        );

    \I__2998\ : Odrv12
    port map (
            O => \N__19207\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__19204\,
            I => \pid_alt.pid_preregZ0Z_5\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19192\
        );

    \I__2995\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19192\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19189\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19185\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19182\
        );

    \I__2991\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19179\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__19185\,
            I => \N__19176\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__19182\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__19179\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__19176\,
            I => \pid_alt.pid_preregZ0Z_12\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__2985\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19161\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19158\
        );

    \I__2983\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19155\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__19161\,
            I => \N__19151\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__19158\,
            I => \N__19146\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19146\
        );

    \I__2979\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19143\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__19151\,
            I => \N__19138\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__19146\,
            I => \N__19138\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__19143\,
            I => \pid_alt.N_130\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__19138\,
            I => \pid_alt.N_130\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19123\
        );

    \I__2971\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19120\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__19123\,
            I => \N__19117\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19114\
        );

    \I__2968\ : Span4Mux_v
    port map (
            O => \N__19117\,
            I => \N__19111\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__19114\,
            I => \N__19108\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__19111\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__19108\,
            I => \ppm_encoder_1.un1_init_pulses_0_1\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__19103\,
            I => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__2962\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__19094\,
            I => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\
        );

    \I__2960\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__2958\ : Span4Mux_s3_h
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__2957\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__19079\,
            I => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19076\,
            I => \ppm_encoder_1.un1_aileron_cry_8\
        );

    \I__2954\ : InMux
    port map (
            O => \N__19073\,
            I => \ppm_encoder_1.un1_aileron_cry_9\
        );

    \I__2953\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__19067\,
            I => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\
        );

    \I__2951\ : InMux
    port map (
            O => \N__19064\,
            I => \ppm_encoder_1.un1_aileron_cry_10\
        );

    \I__2950\ : InMux
    port map (
            O => \N__19061\,
            I => \ppm_encoder_1.un1_aileron_cry_11\
        );

    \I__2949\ : InMux
    port map (
            O => \N__19058\,
            I => \ppm_encoder_1.un1_aileron_cry_12\
        );

    \I__2948\ : InMux
    port map (
            O => \N__19055\,
            I => \bfn_3_22_0_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19048\
        );

    \I__2946\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19045\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19042\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__2942\ : Odrv12
    port map (
            O => \N__19039\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__19036\,
            I => \ppm_encoder_1.aileronZ0Z_14\
        );

    \I__2940\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19027\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__19021\
        );

    \I__2937\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19018\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__19021\,
            I => \N__19013\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__19018\,
            I => \N__19013\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__19013\,
            I => \pid_alt.pid_preregZ0Z_3\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__19010\,
            I => \N__19006\
        );

    \I__2932\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19002\
        );

    \I__2931\ : InMux
    port map (
            O => \N__19006\,
            I => \N__18995\
        );

    \I__2930\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18995\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__19002\,
            I => \N__18991\
        );

    \I__2928\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18986\
        );

    \I__2927\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18986\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__18995\,
            I => \N__18983\
        );

    \I__2925\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18980\
        );

    \I__2924\ : Span4Mux_v
    port map (
            O => \N__18991\,
            I => \N__18975\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__18986\,
            I => \N__18975\
        );

    \I__2922\ : Odrv12
    port map (
            O => \N__18983\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18980\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__18975\,
            I => \pid_alt.pid_preregZ0Z_13\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__18965\,
            I => \N__18961\
        );

    \I__2917\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__2916\ : Odrv12
    port map (
            O => \N__18961\,
            I => \pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__18958\,
            I => \pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6\
        );

    \I__2914\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18947\
        );

    \I__2913\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18947\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__18944\,
            I => \pid_alt.N_88\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\
        );

    \I__2909\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18934\
        );

    \I__2908\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18931\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__18934\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__18931\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__18926\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__18923\,
            I => \pid_alt.N_92_cascade_\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \pid_alt.un1_reset_1_cascade_\
        );

    \I__2902\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__18914\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__18911\,
            I => \pid_alt.un1_reset_0_i_cascade_\
        );

    \I__2899\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__2897\ : Sp12to4
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__2896\ : Odrv12
    port map (
            O => \N__18899\,
            I => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\
        );

    \I__2895\ : InMux
    port map (
            O => \N__18896\,
            I => \ppm_encoder_1.un1_aileron_cry_6\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18893\,
            I => \ppm_encoder_1.un1_aileron_cry_7\
        );

    \I__2893\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__18884\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__2889\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18874\
        );

    \I__2888\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18871\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18865\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18865\
        );

    \I__2885\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18862\
        );

    \I__2884\ : Span4Mux_v
    port map (
            O => \N__18865\,
            I => \N__18857\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__18862\,
            I => \N__18854\
        );

    \I__2882\ : InMux
    port map (
            O => \N__18861\,
            I => \N__18849\
        );

    \I__2881\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18849\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__18857\,
            I => \N__18846\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__18854\,
            I => \N__18841\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__18849\,
            I => \N__18841\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__18846\,
            I => \pid_alt.error_i_regZ0Z_17\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__18841\,
            I => \pid_alt.error_i_regZ0Z_17\
        );

    \I__2875\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18830\
        );

    \I__2874\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18830\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__18830\,
            I => \pid_alt.error_i_acumm_preregZ0Z_17\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__2870\ : Odrv12
    port map (
            O => \N__18821\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO\
        );

    \I__2869\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18812\
        );

    \I__2868\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18812\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__18812\,
            I => \pid_alt.error_i_acumm_preregZ0Z_18\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2865\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18791\
        );

    \I__2864\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18791\
        );

    \I__2863\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18791\
        );

    \I__2862\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18791\
        );

    \I__2861\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18791\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__18785\,
            I => \pid_alt.source_pid_9_0_tz_6\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \pid_alt.source_pid_9_0_tz_6_cascade_\
        );

    \I__2856\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__18776\,
            I => \N__18771\
        );

    \I__2854\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18766\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18766\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__18771\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__18766\,
            I => \pid_alt.pid_preregZ0Z_8\
        );

    \I__2850\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__2848\ : Span4Mux_s2_h
    port map (
            O => \N__18755\,
            I => \N__18750\
        );

    \I__2847\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18747\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18744\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__18750\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__18747\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__18744\,
            I => \pid_alt.pid_preregZ0Z_11\
        );

    \I__2842\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18733\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__18736\,
            I => \N__18730\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18726\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18723\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18720\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__18726\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__18723\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__18720\,
            I => \pid_alt.pid_preregZ0Z_9\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__18713\,
            I => \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18702\
        );

    \I__2831\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18699\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__18705\,
            I => \N__18696\
        );

    \I__2829\ : Span4Mux_v
    port map (
            O => \N__18702\,
            I => \N__18693\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__18699\,
            I => \N__18690\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18696\,
            I => \N__18687\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__18693\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__18690\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__18687\,
            I => \pid_alt.pid_preregZ0Z_6\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18673\
        );

    \I__2821\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18670\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__2818\ : Odrv12
    port map (
            O => \N__18667\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__18664\,
            I => \pid_alt.pid_preregZ0Z_0\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__18656\,
            I => \N__18651\
        );

    \I__2814\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18646\
        );

    \I__2813\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18646\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__18651\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__18646\,
            I => \pid_alt.pid_preregZ0Z_10\
        );

    \I__2810\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18633\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18628\
        );

    \I__2807\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18628\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__18633\,
            I => \pid_alt.pid_preregZ0Z_7\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__18628\,
            I => \pid_alt.pid_preregZ0Z_7\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__18614\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18608\,
            I => \N__18605\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__18605\,
            I => \N__18601\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18598\
        );

    \I__2796\ : Span4Mux_v
    port map (
            O => \N__18601\,
            I => \N__18591\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__18598\,
            I => \N__18591\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18597\,
            I => \N__18586\
        );

    \I__2793\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18586\
        );

    \I__2792\ : Span4Mux_v
    port map (
            O => \N__18591\,
            I => \N__18582\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__18586\,
            I => \N__18579\
        );

    \I__2790\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18576\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__18582\,
            I => \N__18573\
        );

    \I__2788\ : Odrv12
    port map (
            O => \N__18579\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__18576\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__18573\,
            I => \pid_alt.error_i_regZ0Z_19\
        );

    \I__2785\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__18563\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__18560\,
            I => \N__18556\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__18559\,
            I => \N__18553\
        );

    \I__2781\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18549\
        );

    \I__2780\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18544\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18544\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__18549\,
            I => \pid_alt.error_i_acumm_preregZ0Z_19\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__18544\,
            I => \pid_alt.error_i_acumm_preregZ0Z_19\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18535\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18538\,
            I => \N__18532\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__18535\,
            I => \N__18529\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__18532\,
            I => \N__18526\
        );

    \I__2772\ : Span4Mux_v
    port map (
            O => \N__18529\,
            I => \N__18522\
        );

    \I__2771\ : Span12Mux_v
    port map (
            O => \N__18526\,
            I => \N__18519\
        );

    \I__2770\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18516\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__18522\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__2768\ : Odrv12
    port map (
            O => \N__18519\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__18516\,
            I => \pid_alt.error_p_regZ0Z_16\
        );

    \I__2766\ : InMux
    port map (
            O => \N__18509\,
            I => \N__18504\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18499\
        );

    \I__2764\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18499\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__18504\,
            I => \N__18493\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__18499\,
            I => \N__18493\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__18498\,
            I => \N__18490\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__18493\,
            I => \N__18486\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18490\,
            I => \N__18483\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18489\,
            I => \N__18480\
        );

    \I__2757\ : Span4Mux_h
    port map (
            O => \N__18486\,
            I => \N__18477\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__18483\,
            I => \N__18474\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__18480\,
            I => \N__18471\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__18477\,
            I => \N__18468\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__18474\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__18471\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__18468\,
            I => \pid_alt.error_i_regZ0Z_16\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__2747\ : Span4Mux_h
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__18449\,
            I => \pid_alt.error_p_reg_esr_RNIB03KZ0Z_16\
        );

    \I__2745\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__2743\ : Span4Mux_v
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__18434\,
            I => \ppm_encoder_1.N_306\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__18431\,
            I => \dron_frame_decoder_1.N_194_4_cascade_\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \N__18424\
        );

    \I__2738\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__2737\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__18421\,
            I => \pid_alt.error_i_acumm_preregZ0Z_20\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__18418\,
            I => \pid_alt.error_i_acumm_preregZ0Z_20\
        );

    \I__2734\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18407\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18407\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__18407\,
            I => \pid_alt.m7_e_4\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__18398\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__2727\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18389\,
            I => \N__18385\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__18388\,
            I => \N__18382\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__18385\,
            I => \N__18378\
        );

    \I__2723\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18375\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18372\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__18378\,
            I => \N__18367\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__18375\,
            I => \N__18364\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18357\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18357\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18357\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__18367\,
            I => \N__18352\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__18364\,
            I => \N__18352\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__18357\,
            I => \N__18349\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__18352\,
            I => \pid_alt.error_i_regZ0Z_15\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__18349\,
            I => \pid_alt.error_i_regZ0Z_15\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18338\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18343\,
            I => \N__18338\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__18338\,
            I => \pid_alt.error_i_acumm_preregZ0Z_15\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18335\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_16\
        );

    \I__2707\ : InMux
    port map (
            O => \N__18332\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_17\
        );

    \I__2706\ : InMux
    port map (
            O => \N__18329\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_18\
        );

    \I__2705\ : InMux
    port map (
            O => \N__18326\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18323\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_20\
        );

    \I__2703\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18312\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18312\
        );

    \I__2701\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18307\
        );

    \I__2700\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18307\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__18312\,
            I => \N__18304\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18307\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__18304\,
            I => \pid_alt.error_i_acumm_preregZ0Z_21\
        );

    \I__2696\ : CEMux
    port map (
            O => \N__18299\,
            I => \N__18281\
        );

    \I__2695\ : CEMux
    port map (
            O => \N__18298\,
            I => \N__18281\
        );

    \I__2694\ : CEMux
    port map (
            O => \N__18297\,
            I => \N__18281\
        );

    \I__2693\ : CEMux
    port map (
            O => \N__18296\,
            I => \N__18281\
        );

    \I__2692\ : CEMux
    port map (
            O => \N__18295\,
            I => \N__18281\
        );

    \I__2691\ : CEMux
    port map (
            O => \N__18294\,
            I => \N__18281\
        );

    \I__2690\ : GlobalMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__2689\ : gio2CtrlBuf
    port map (
            O => \N__18278\,
            I => \pid_alt.state_0_g_0\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__18272\,
            I => \N__18268\
        );

    \I__2686\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18265\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__18268\,
            I => \N__18259\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__18265\,
            I => \N__18259\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18264\,
            I => \N__18256\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__18259\,
            I => \N__18253\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__18256\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__18253\,
            I => \pid_alt.error_i_acummZ0Z_0\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__18248\,
            I => \N__18244\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18237\
        );

    \I__2676\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18234\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__18240\,
            I => \N__18231\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18228\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18225\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18222\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__18228\,
            I => \N__18219\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__18225\,
            I => \N__18214\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__18222\,
            I => \N__18214\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__18219\,
            I => \N__18211\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__18214\,
            I => \N__18208\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__18211\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__18208\,
            I => \pid_alt.error_i_regZ0Z_0\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18199\
        );

    \I__2663\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18196\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__18199\,
            I => \N__18192\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__18196\,
            I => \N__18189\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18186\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__18192\,
            I => \N__18183\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__18189\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18186\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__18183\,
            I => \pid_alt.error_i_acumm_preregZ0Z_0\
        );

    \I__2655\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__18170\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__18164\,
            I => \N__18161\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__18161\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__18158\,
            I => \N__18154\
        );

    \I__2648\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18151\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18148\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__18151\,
            I => \N__18145\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__18148\,
            I => \N__18140\
        );

    \I__2644\ : Span4Mux_h
    port map (
            O => \N__18145\,
            I => \N__18137\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__18144\,
            I => \N__18134\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18130\
        );

    \I__2641\ : Span12Mux_v
    port map (
            O => \N__18140\,
            I => \N__18127\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__18137\,
            I => \N__18124\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18119\
        );

    \I__2638\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18119\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__18130\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2636\ : Odrv12
    port map (
            O => \N__18127\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__18124\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18119\,
            I => \pid_alt.error_i_regZ0Z_14\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18105\
        );

    \I__2632\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18100\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18100\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__18105\,
            I => \pid_alt.error_i_acumm_preregZ0Z_14\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__18100\,
            I => \pid_alt.error_i_acumm_preregZ0Z_14\
        );

    \I__2628\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__18092\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18081\
        );

    \I__2624\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18076\
        );

    \I__2623\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18076\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__18081\,
            I => \pid_alt.error_i_acumm_preregZ0Z_16\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__18076\,
            I => \pid_alt.error_i_acumm_preregZ0Z_16\
        );

    \I__2620\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__18065\,
            I => \N__18060\
        );

    \I__2617\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18055\
        );

    \I__2616\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18055\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__18060\,
            I => \pid_alt.error_i_regZ0Z_9\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__18055\,
            I => \pid_alt.error_i_regZ0Z_9\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \N__18044\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__18049\,
            I => \N__18041\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18036\
        );

    \I__2610\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18036\
        );

    \I__2609\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18033\
        );

    \I__2608\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18030\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__18036\,
            I => \N__18027\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__18033\,
            I => \N__18022\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__18030\,
            I => \N__18022\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__18027\,
            I => \N__18019\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__18022\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__18019\,
            I => \pid_alt.error_i_acummZ0Z_9\
        );

    \I__2601\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18011\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__18011\,
            I => \N__18006\
        );

    \I__2599\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18001\
        );

    \I__2598\ : InMux
    port map (
            O => \N__18009\,
            I => \N__18001\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__18006\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__18001\,
            I => \pid_alt.error_i_acumm_preregZ0Z_9\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17996\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_8\
        );

    \I__2594\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__17987\,
            I => \N__17982\
        );

    \I__2591\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17977\
        );

    \I__2590\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17977\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__17982\,
            I => \pid_alt.error_i_regZ0Z_10\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__17977\,
            I => \pid_alt.error_i_regZ0Z_10\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__17972\,
            I => \N__17968\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17963\
        );

    \I__2585\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17960\
        );

    \I__2584\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17955\
        );

    \I__2583\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17955\
        );

    \I__2582\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17952\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__17960\,
            I => \N__17949\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__17955\,
            I => \N__17946\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__17952\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__17949\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__17946\,
            I => \pid_alt.error_i_acummZ0Z_10\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17935\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__17938\,
            I => \N__17932\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__17935\,
            I => \N__17928\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17923\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17923\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__17928\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__17923\,
            I => \pid_alt.error_i_acumm_preregZ0Z_10\
        );

    \I__2569\ : InMux
    port map (
            O => \N__17918\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_9\
        );

    \I__2568\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__17909\,
            I => \N__17904\
        );

    \I__2565\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17899\
        );

    \I__2564\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17899\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__17904\,
            I => \pid_alt.error_i_regZ0Z_11\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__17899\,
            I => \pid_alt.error_i_regZ0Z_11\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17889\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__17893\,
            I => \N__17885\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__17892\,
            I => \N__17882\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17889\,
            I => \N__17879\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17874\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17874\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17871\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__17879\,
            I => \N__17868\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17874\,
            I => \N__17865\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__17871\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__17868\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__17865\,
            I => \pid_alt.error_i_acummZ0Z_11\
        );

    \I__2549\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17854\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__17857\,
            I => \N__17850\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__17854\,
            I => \N__17847\
        );

    \I__2546\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17842\
        );

    \I__2545\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17842\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__17847\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__17842\,
            I => \pid_alt.error_i_acumm_preregZ0Z_11\
        );

    \I__2542\ : InMux
    port map (
            O => \N__17837\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_10\
        );

    \I__2541\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17831\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__17828\,
            I => \N__17823\
        );

    \I__2538\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17818\
        );

    \I__2537\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17818\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__17823\,
            I => \pid_alt.error_i_regZ0Z_12\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__17818\,
            I => \pid_alt.error_i_regZ0Z_12\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__17813\,
            I => \N__17809\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \N__17804\
        );

    \I__2532\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17801\
        );

    \I__2531\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17796\
        );

    \I__2530\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17796\
        );

    \I__2529\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17793\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__17801\,
            I => \N__17790\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__17796\,
            I => \N__17787\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__17793\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__17790\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__17787\,
            I => \pid_alt.error_i_acummZ0Z_12\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__2522\ : InMux
    port map (
            O => \N__17777\,
            I => \N__17773\
        );

    \I__2521\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17770\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__17773\,
            I => \N__17767\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17763\
        );

    \I__2518\ : Span4Mux_h
    port map (
            O => \N__17767\,
            I => \N__17760\
        );

    \I__2517\ : InMux
    port map (
            O => \N__17766\,
            I => \N__17757\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__17763\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__17760\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__17757\,
            I => \pid_alt.error_i_acumm7lto12\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17750\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_11\
        );

    \I__2512\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__2511\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17741\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17737\
        );

    \I__2509\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__17737\,
            I => \N__17731\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__17731\,
            I => \N__17725\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__17728\,
            I => \pid_alt.error_i_acummZ0Z_13\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__17725\,
            I => \pid_alt.error_i_acummZ0Z_13\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__2502\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__17711\,
            I => \N__17706\
        );

    \I__2499\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17703\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17700\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__17706\,
            I => \N__17697\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__17703\,
            I => \N__17692\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__17700\,
            I => \N__17692\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__17697\,
            I => \pid_alt.error_i_regZ0Z_13\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__17692\,
            I => \pid_alt.error_i_regZ0Z_13\
        );

    \I__2492\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17678\
        );

    \I__2491\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17678\
        );

    \I__2490\ : InMux
    port map (
            O => \N__17685\,
            I => \N__17678\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__17675\,
            I => \pid_alt.error_i_acumm7lto13\
        );

    \I__2487\ : InMux
    port map (
            O => \N__17672\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_12\
        );

    \I__2486\ : InMux
    port map (
            O => \N__17669\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_13\
        );

    \I__2485\ : InMux
    port map (
            O => \N__17666\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_14\
        );

    \I__2484\ : InMux
    port map (
            O => \N__17663\,
            I => \bfn_3_15_0_\
        );

    \I__2483\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17652\
        );

    \I__2481\ : InMux
    port map (
            O => \N__17656\,
            I => \N__17647\
        );

    \I__2480\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17647\
        );

    \I__2479\ : Span4Mux_h
    port map (
            O => \N__17652\,
            I => \N__17644\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__17644\,
            I => \pid_alt.error_i_regZ0Z_2\
        );

    \I__2476\ : Odrv12
    port map (
            O => \N__17641\,
            I => \pid_alt.error_i_regZ0Z_2\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__2474\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__17630\,
            I => \N__17626\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__17629\,
            I => \N__17623\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__17626\,
            I => \N__17619\
        );

    \I__2470\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17614\
        );

    \I__2469\ : InMux
    port map (
            O => \N__17622\,
            I => \N__17614\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__17619\,
            I => \pid_alt.error_i_acummZ0Z_2\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__17614\,
            I => \pid_alt.error_i_acummZ0Z_2\
        );

    \I__2466\ : InMux
    port map (
            O => \N__17609\,
            I => \N__17606\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__2464\ : Span4Mux_s3_h
    port map (
            O => \N__17603\,
            I => \N__17599\
        );

    \I__2463\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17596\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__17599\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__17596\,
            I => \pid_alt.error_i_acumm_preregZ0Z_2\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17591\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_1\
        );

    \I__2459\ : InMux
    port map (
            O => \N__17588\,
            I => \N__17583\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17578\
        );

    \I__2457\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17578\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__17583\,
            I => \N__17575\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17572\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__17575\,
            I => \pid_alt.error_i_regZ0Z_3\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__17572\,
            I => \pid_alt.error_i_regZ0Z_3\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__2451\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__17561\,
            I => \N__17557\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__17560\,
            I => \N__17554\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__17557\,
            I => \N__17550\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17545\
        );

    \I__2446\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17545\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__17550\,
            I => \pid_alt.error_i_acummZ0Z_3\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__17545\,
            I => \pid_alt.error_i_acummZ0Z_3\
        );

    \I__2443\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__17534\,
            I => \N__17530\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17527\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__17530\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__17527\,
            I => \pid_alt.error_i_acumm_preregZ0Z_3\
        );

    \I__2437\ : InMux
    port map (
            O => \N__17522\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_2\
        );

    \I__2436\ : InMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__17513\,
            I => \N__17508\
        );

    \I__2433\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17503\
        );

    \I__2432\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17503\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__17508\,
            I => \pid_alt.error_i_acummZ0Z_4\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__17503\,
            I => \pid_alt.error_i_acummZ0Z_4\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__17498\,
            I => \N__17494\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \N__17491\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17487\
        );

    \I__2426\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17482\
        );

    \I__2425\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17482\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__17487\,
            I => \N__17479\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__17482\,
            I => \N__17476\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__17479\,
            I => \pid_alt.error_i_regZ0Z_4\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__17476\,
            I => \pid_alt.error_i_regZ0Z_4\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__17471\,
            I => \N__17467\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__17470\,
            I => \N__17461\
        );

    \I__2418\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17456\
        );

    \I__2417\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17456\
        );

    \I__2416\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17453\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17464\,
            I => \N__17450\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17447\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__17456\,
            I => \N__17442\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__17453\,
            I => \N__17442\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17437\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17437\
        );

    \I__2409\ : Span4Mux_s3_h
    port map (
            O => \N__17442\,
            I => \N__17433\
        );

    \I__2408\ : Span4Mux_s3_h
    port map (
            O => \N__17437\,
            I => \N__17430\
        );

    \I__2407\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17427\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__17433\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__17430\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__17427\,
            I => \pid_alt.error_i_acumm7lto4\
        );

    \I__2403\ : InMux
    port map (
            O => \N__17420\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_3\
        );

    \I__2402\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17412\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17408\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__17415\,
            I => \N__17405\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17412\,
            I => \N__17402\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17399\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__17408\,
            I => \N__17396\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17393\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__17402\,
            I => \N__17390\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__17399\,
            I => \N__17385\
        );

    \I__2393\ : Span12Mux_s8_v
    port map (
            O => \N__17396\,
            I => \N__17385\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__17393\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__17390\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__17385\,
            I => \pid_alt.error_i_acummZ0Z_5\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__17378\,
            I => \N__17374\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17370\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17367\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17364\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__17370\,
            I => \N__17361\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17358\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__17364\,
            I => \N__17355\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__17361\,
            I => \N__17352\
        );

    \I__2381\ : Odrv12
    port map (
            O => \N__17358\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__2380\ : Odrv12
    port map (
            O => \N__17355\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__17352\,
            I => \pid_alt.error_i_regZ0Z_5\
        );

    \I__2378\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17340\
        );

    \I__2377\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17337\
        );

    \I__2376\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17334\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__17340\,
            I => \N__17329\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__17337\,
            I => \N__17329\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17334\,
            I => \N__17326\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__17329\,
            I => \N__17321\
        );

    \I__2371\ : Span4Mux_s3_h
    port map (
            O => \N__17326\,
            I => \N__17318\
        );

    \I__2370\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17313\
        );

    \I__2369\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17313\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__17321\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__17318\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__17313\,
            I => \pid_alt.error_i_acumm7lto5\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17306\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_4\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17300\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__17300\,
            I => \N__17297\
        );

    \I__2362\ : Span4Mux_s3_h
    port map (
            O => \N__17297\,
            I => \N__17292\
        );

    \I__2361\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17287\
        );

    \I__2360\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17287\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__17292\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__17287\,
            I => \pid_alt.error_i_acumm_preregZ0Z_6\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17282\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_5\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17272\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__17272\,
            I => \N__17265\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17260\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17260\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__17265\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__17260\,
            I => \pid_alt.error_i_acumm_preregZ0Z_7\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17255\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_6\
        );

    \I__2347\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17249\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__17246\,
            I => \N__17241\
        );

    \I__2344\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17236\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17236\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__17241\,
            I => \pid_alt.error_i_regZ0Z_8\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__17236\,
            I => \pid_alt.error_i_regZ0Z_8\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \N__17227\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__17230\,
            I => \N__17222\
        );

    \I__2338\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17217\
        );

    \I__2337\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17217\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__17225\,
            I => \N__17214\
        );

    \I__2335\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17211\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__17217\,
            I => \N__17208\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17205\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17211\,
            I => \N__17202\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__17208\,
            I => \N__17199\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__17205\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__2329\ : Odrv12
    port map (
            O => \N__17202\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__17199\,
            I => \pid_alt.error_i_acummZ0Z_8\
        );

    \I__2327\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17184\
        );

    \I__2325\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17179\
        );

    \I__2324\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17179\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__17184\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__17179\,
            I => \pid_alt.error_i_acumm_preregZ0Z_8\
        );

    \I__2321\ : InMux
    port map (
            O => \N__17174\,
            I => \bfn_3_14_0_\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17168\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__17168\,
            I => \pid_alt.error_axbZ0Z_12\
        );

    \I__2318\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__17162\,
            I => drone_altitude_12
        );

    \I__2316\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17156\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__17156\,
            I => \pid_alt.error_axbZ0Z_13\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__17150\,
            I => drone_altitude_13
        );

    \I__2312\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__17144\,
            I => \pid_alt.error_axbZ0Z_14\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__17141\,
            I => \N__17138\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17135\,
            I => \pid_alt.error_axbZ0Z_2\
        );

    \I__2307\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17129\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__17129\,
            I => \pid_alt.error_axbZ0Z_3\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17120\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__17120\,
            I => \N__17115\
        );

    \I__2302\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17110\
        );

    \I__2301\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17110\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__17115\,
            I => \pid_alt.error_i_acummZ0Z_1\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17110\,
            I => \pid_alt.error_i_acummZ0Z_1\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17097\
        );

    \I__2296\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17092\
        );

    \I__2295\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17092\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__17097\,
            I => \N__17089\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__17089\,
            I => \pid_alt.error_i_regZ0Z_1\
        );

    \I__2291\ : Odrv12
    port map (
            O => \N__17086\,
            I => \pid_alt.error_i_regZ0Z_1\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__17081\,
            I => \N__17078\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__2286\ : Span4Mux_s1_h
    port map (
            O => \N__17069\,
            I => \N__17065\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__17065\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__17062\,
            I => \pid_alt.error_i_acumm_preregZ0Z_1\
        );

    \I__2282\ : InMux
    port map (
            O => \N__17057\,
            I => \pid_alt.un1_error_i_acumm_prereg_cry_0\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__17054\,
            I => \Commands_frame_decoder.source_CH1data8_cascade_\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__17051\,
            I => \N__17047\
        );

    \I__2279\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__2278\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17041\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__17044\,
            I => alt_command_0
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__17041\,
            I => alt_command_0
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__2274\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__17030\,
            I => drone_altitude_i_7
        );

    \I__2272\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__17024\,
            I => \dron_frame_decoder_1.drone_altitude_7\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__17018\,
            I => drone_altitude_i_8
        );

    \I__2268\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__17012\,
            I => drone_altitude_i_9
        );

    \I__2266\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__17006\,
            I => drone_altitude_i_10
        );

    \I__2264\ : InMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__17000\,
            I => drone_altitude_i_11
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__2261\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__16991\,
            I => \pid_alt.error_axbZ0Z_1\
        );

    \I__2259\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__16985\,
            I => drone_altitude_1
        );

    \I__2257\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__16979\,
            I => \N__16976\
        );

    \I__2255\ : Span4Mux_s3_h
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__16973\,
            I => alt_kp_6
        );

    \I__2253\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__16967\,
            I => \N__16964\
        );

    \I__2251\ : Span4Mux_s3_h
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__16961\,
            I => alt_kp_5
        );

    \I__2249\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__2247\ : Span4Mux_s3_h
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__16949\,
            I => alt_kp_1
        );

    \I__2245\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16940\
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__16940\,
            I => alt_kp_0
        );

    \I__2242\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2240\ : Span4Mux_s3_h
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__16928\,
            I => drone_altitude_15
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__16925\,
            I => \N__16921\
        );

    \I__2237\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__2236\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16915\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__16918\,
            I => alt_command_2
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__16915\,
            I => alt_command_2
        );

    \I__2233\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16903\
        );

    \I__2231\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16900\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__16903\,
            I => \N__16897\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__16900\,
            I => alt_command_3
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__16897\,
            I => alt_command_3
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__16892\,
            I => \N__16888\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__2225\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__16885\,
            I => alt_command_1
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__16882\,
            I => alt_command_1
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__16874\,
            I => \N__16870\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \N__16867\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16859\
        );

    \I__2218\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16859\
        );

    \I__2217\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16859\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__16859\,
            I => \Commands_frame_decoder.source_CH1data8\
        );

    \I__2215\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__16853\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__16850\,
            I => \N__16847\
        );

    \I__2212\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__16844\,
            I => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__16838\,
            I => \ppm_encoder_1.un1_init_pulses_11_13\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16835\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_12\
        );

    \I__2207\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__16829\,
            I => \ppm_encoder_1.un1_init_pulses_11_14\
        );

    \I__2205\ : InMux
    port map (
            O => \N__16826\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_13\
        );

    \I__2204\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__16817\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_15\
        );

    \I__2201\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__16811\,
            I => \ppm_encoder_1.un1_init_pulses_11_15\
        );

    \I__2199\ : InMux
    port map (
            O => \N__16808\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_14\
        );

    \I__2198\ : InMux
    port map (
            O => \N__16805\,
            I => \bfn_2_30_0_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__16796\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_17\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__16787\,
            I => \ppm_encoder_1.un1_init_pulses_11_17\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16784\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_16\
        );

    \I__2190\ : InMux
    port map (
            O => \N__16781\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_17\
        );

    \I__2189\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__16775\,
            I => \ppm_encoder_1.un1_init_pulses_11_18\
        );

    \I__2187\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16769\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__2185\ : Span4Mux_s3_h
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__16763\,
            I => alt_kp_3
        );

    \I__2183\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__2181\ : Span4Mux_s3_v
    port map (
            O => \N__16754\,
            I => \N__16751\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__16751\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_5\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16748\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_4\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__16742\,
            I => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16739\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_5\
        );

    \I__2175\ : InMux
    port map (
            O => \N__16736\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_6\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__16727\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_8\
        );

    \I__2171\ : InMux
    port map (
            O => \N__16724\,
            I => \bfn_2_29_0_\
        );

    \I__2170\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__2168\ : Span4Mux_s2_v
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__16712\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_9\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__16703\,
            I => \ppm_encoder_1.un1_init_pulses_11_9\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16700\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_8\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16694\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__16694\,
            I => \ppm_encoder_1.un1_init_pulses_11_10\
        );

    \I__2160\ : InMux
    port map (
            O => \N__16691\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_9\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__16685\,
            I => \ppm_encoder_1.un1_init_pulses_11_11\
        );

    \I__2157\ : InMux
    port map (
            O => \N__16682\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_10\
        );

    \I__2156\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__16676\,
            I => \ppm_encoder_1.un1_init_pulses_11_12\
        );

    \I__2154\ : InMux
    port map (
            O => \N__16673\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_11\
        );

    \I__2153\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__16667\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_18\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__16661\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_16\
        );

    \I__2149\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__16655\,
            I => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__16646\,
            I => \ppm_encoder_1.un1_init_pulses_3_axb_1\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__16640\,
            I => \ppm_encoder_1.un1_init_pulses_11_1\
        );

    \I__2142\ : InMux
    port map (
            O => \N__16637\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_0\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16634\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_1\
        );

    \I__2140\ : InMux
    port map (
            O => \N__16631\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_2\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16628\,
            I => \ppm_encoder_1.un1_init_pulses_3_cry_3\
        );

    \I__2138\ : InMux
    port map (
            O => \N__16625\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_10\
        );

    \I__2137\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__2135\ : Span4Mux_s2_v
    port map (
            O => \N__16616\,
            I => \N__16613\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__16613\,
            I => \ppm_encoder_1.un1_init_pulses_10_12\
        );

    \I__2133\ : InMux
    port map (
            O => \N__16610\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_11\
        );

    \I__2132\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__16604\,
            I => \N__16600\
        );

    \I__2130\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16597\
        );

    \I__2129\ : Span4Mux_v
    port map (
            O => \N__16600\,
            I => \N__16592\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__16597\,
            I => \N__16592\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__16589\,
            I => \ppm_encoder_1.un1_init_pulses_0_13\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__16586\,
            I => \N__16583\
        );

    \I__2124\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__16577\,
            I => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\
        );

    \I__2121\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16568\
        );

    \I__2119\ : Span4Mux_s1_v
    port map (
            O => \N__16568\,
            I => \N__16565\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__16565\,
            I => \ppm_encoder_1.un1_init_pulses_10_13\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16562\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_12\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16556\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__16556\,
            I => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__16553\,
            I => \N__16549\
        );

    \I__2113\ : InMux
    port map (
            O => \N__16552\,
            I => \N__16546\
        );

    \I__2112\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16543\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16546\,
            I => \N__16538\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__16543\,
            I => \N__16538\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__16535\,
            I => \ppm_encoder_1.un1_init_pulses_0_14\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__2106\ : InMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__16523\,
            I => \ppm_encoder_1.un1_init_pulses_10_14\
        );

    \I__2103\ : InMux
    port map (
            O => \N__16520\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_13\
        );

    \I__2102\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__16511\,
            I => \N__16508\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__16508\,
            I => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__2097\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__2095\ : Span4Mux_h
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__16493\,
            I => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__2091\ : Span4Mux_s1_v
    port map (
            O => \N__16484\,
            I => \N__16481\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__16481\,
            I => \ppm_encoder_1.un1_init_pulses_10_15\
        );

    \I__2089\ : InMux
    port map (
            O => \N__16478\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_14\
        );

    \I__2088\ : InMux
    port map (
            O => \N__16475\,
            I => \bfn_2_27_0_\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__16466\,
            I => \ppm_encoder_1.un1_init_pulses_10_17\
        );

    \I__2084\ : InMux
    port map (
            O => \N__16463\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_16\
        );

    \I__2083\ : InMux
    port map (
            O => \N__16460\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_17\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \N__16454\
        );

    \I__2081\ : InMux
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__16448\,
            I => \ppm_encoder_1.un1_init_pulses_10_18\
        );

    \I__2078\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16442\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__16442\,
            I => \ppm_encoder_1.un1_init_pulses_0_axb_17\
        );

    \I__2076\ : InMux
    port map (
            O => \N__16439\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_2\
        );

    \I__2075\ : InMux
    port map (
            O => \N__16436\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_3\
        );

    \I__2074\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16429\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16426\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__16429\,
            I => \N__16423\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16420\
        );

    \I__2070\ : Span4Mux_h
    port map (
            O => \N__16423\,
            I => \N__16417\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__16420\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__16417\,
            I => \ppm_encoder_1.un1_init_pulses_0_5\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__16412\,
            I => \N__16409\
        );

    \I__2066\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__16406\,
            I => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\
        );

    \I__2064\ : InMux
    port map (
            O => \N__16403\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_4\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2062\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16394\,
            I => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16391\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_5\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__2058\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__16382\,
            I => \N__16379\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__16379\,
            I => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\
        );

    \I__2055\ : InMux
    port map (
            O => \N__16376\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_6\
        );

    \I__2054\ : InMux
    port map (
            O => \N__16373\,
            I => \bfn_2_26_0_\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__16364\,
            I => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__2049\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16355\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__16355\,
            I => \ppm_encoder_1.un1_init_pulses_10_9\
        );

    \I__2047\ : InMux
    port map (
            O => \N__16352\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_8\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__2045\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16343\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__16343\,
            I => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\
        );

    \I__2043\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__16334\,
            I => \ppm_encoder_1.un1_init_pulses_10_10\
        );

    \I__2040\ : InMux
    port map (
            O => \N__16331\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_9\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__16328\,
            I => \N__16325\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16325\,
            I => \N__16322\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__2036\ : Odrv12
    port map (
            O => \N__16319\,
            I => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__16316\,
            I => \N__16313\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16310\,
            I => \N__16307\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__16307\,
            I => \ppm_encoder_1.un1_init_pulses_10_11\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__16304\,
            I => \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__16301\,
            I => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\
        );

    \I__2029\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16295\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__16295\,
            I => \ppm_encoder_1.un2_throttle_iv_1_6\
        );

    \I__2027\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16289\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__16289\,
            I => \ppm_encoder_1.un2_throttle_iv_0_13\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16282\
        );

    \I__2024\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16279\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__16282\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__16279\,
            I => \ppm_encoder_1.aileronZ0Z_5\
        );

    \I__2021\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16270\
        );

    \I__2020\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16267\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__16270\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__16267\,
            I => \ppm_encoder_1.elevatorZ0Z_5\
        );

    \I__2017\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16259\,
            I => \ppm_encoder_1.un2_throttle_iv_1_5\
        );

    \I__2015\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__16253\,
            I => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\
        );

    \I__2013\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16247\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__2011\ : Span4Mux_s3_v
    port map (
            O => \N__16244\,
            I => \N__16241\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__16241\,
            I => \ppm_encoder_1.un1_init_pulses_10_1\
        );

    \I__2009\ : InMux
    port map (
            O => \N__16238\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_0\
        );

    \I__2008\ : InMux
    port map (
            O => \N__16235\,
            I => \ppm_encoder_1.un1_init_pulses_0_cry_1\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__16232\,
            I => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16226\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__16226\,
            I => \ppm_encoder_1.un2_throttle_iv_1_7\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__16223\,
            I => \ppm_encoder_1.N_299_cascade_\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16211\
        );

    \I__2002\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16211\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16218\,
            I => \N__16211\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16211\,
            I => \ppm_encoder_1.aileronZ0Z_7\
        );

    \I__1999\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16199\
        );

    \I__1998\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16199\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16199\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__16199\,
            I => \ppm_encoder_1.elevatorZ0Z_7\
        );

    \I__1995\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__16190\,
            I => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16179\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16176\
        );

    \I__1989\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16173\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16179\,
            I => \N__16168\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16168\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__16173\,
            I => \N__16165\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__16168\,
            I => throttle_command_7
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__16165\,
            I => throttle_command_7
        );

    \I__1983\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16151\
        );

    \I__1982\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16151\
        );

    \I__1981\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16151\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__16151\,
            I => \ppm_encoder_1.throttleZ0Z_7\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\
        );

    \I__1978\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__16142\,
            I => \ppm_encoder_1.un2_throttle_iv_1_11\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__16139\,
            I => \ppm_encoder_1.N_303_cascade_\
        );

    \I__1975\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16127\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16127\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16127\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16127\,
            I => \ppm_encoder_1.aileronZ0Z_11\
        );

    \I__1971\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16115\
        );

    \I__1970\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16115\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16115\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16115\,
            I => \ppm_encoder_1.elevatorZ0Z_11\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__16109\,
            I => \N__16104\
        );

    \I__1965\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16101\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16098\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__16104\,
            I => \N__16095\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__16101\,
            I => \N__16092\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__16098\,
            I => throttle_command_11
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__16095\,
            I => throttle_command_11
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__16092\,
            I => throttle_command_11
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__16085\,
            I => \N__16082\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16079\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__16079\,
            I => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\
        );

    \I__1955\ : InMux
    port map (
            O => \N__16076\,
            I => \N__16067\
        );

    \I__1954\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16067\
        );

    \I__1953\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16067\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__16067\,
            I => \ppm_encoder_1.throttleZ0Z_11\
        );

    \I__1951\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16061\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__16058\,
            I => \pid_alt.pid_preregZ0Z_14\
        );

    \I__1948\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16052\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__16052\,
            I => \pid_alt.pid_preregZ0Z_19\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__16049\,
            I => \N__16046\
        );

    \I__1945\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__16043\,
            I => \pid_alt.pid_preregZ0Z_20\
        );

    \I__1943\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__16037\,
            I => \pid_alt.pid_preregZ0Z_21\
        );

    \I__1941\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__16031\,
            I => \pid_alt.pid_preregZ0Z_16\
        );

    \I__1939\ : InMux
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__16025\,
            I => \pid_alt.pid_preregZ0Z_15\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__16022\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__16019\,
            I => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_\
        );

    \I__1935\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__16013\,
            I => \pid_alt.pid_preregZ0Z_17\
        );

    \I__1933\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__16007\,
            I => \pid_alt.pid_preregZ0Z_18\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16004\,
            I => \N__16001\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__16001\,
            I => \pid_alt.source_pid_1_sqmuxa_0_a2_2_3\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__1928\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15992\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__15992\,
            I => \pid_alt.source_pid_9_0_0_4\
        );

    \I__1926\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15986\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__15986\,
            I => \N__15982\
        );

    \I__1924\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15979\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__15982\,
            I => throttle_command_5
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__15979\,
            I => throttle_command_5
        );

    \I__1921\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__1919\ : Span12Mux_v
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__15965\,
            I => \pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__1916\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15956\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__1914\ : Span12Mux_h
    port map (
            O => \N__15953\,
            I => \N__15950\
        );

    \I__1913\ : Span12Mux_v
    port map (
            O => \N__15950\,
            I => \N__15947\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__15947\,
            I => \pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14\
        );

    \I__1911\ : InMux
    port map (
            O => \N__15944\,
            I => \bfn_2_19_0_\
        );

    \I__1910\ : InMux
    port map (
            O => \N__15941\,
            I => \N__15938\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__15938\,
            I => \N__15935\
        );

    \I__1908\ : Span12Mux_s3_h
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__1907\ : Span12Mux_v
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__1906\ : Odrv12
    port map (
            O => \N__15929\,
            I => \pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__1904\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__1902\ : Span12Mux_v
    port map (
            O => \N__15917\,
            I => \N__15914\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__15914\,
            I => \pid_alt.error_p_reg_esr_RNIKU581Z0Z_15\
        );

    \I__1900\ : InMux
    port map (
            O => \N__15911\,
            I => \pid_alt.un1_pid_prereg_0_cry_15\
        );

    \I__1899\ : InMux
    port map (
            O => \N__15908\,
            I => \N__15905\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__15905\,
            I => \N__15902\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__15899\,
            I => \pid_alt.error_p_reg_esr_RNIO2681Z0Z_16\
        );

    \I__1895\ : InMux
    port map (
            O => \N__15896\,
            I => \pid_alt.un1_pid_prereg_0_cry_16\
        );

    \I__1894\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__15887\,
            I => \N__15884\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__15881\,
            I => \pid_alt.error_p_reg_esr_RNID23KZ0Z_17\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__1888\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15872\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__15872\,
            I => \N__15869\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__15869\,
            I => \pid_alt.error_p_reg_esr_RNIS6681Z0Z_17\
        );

    \I__1885\ : InMux
    port map (
            O => \N__15866\,
            I => \pid_alt.un1_pid_prereg_0_cry_17\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \N__15860\
        );

    \I__1883\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15857\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__15857\,
            I => \N__15854\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__15854\,
            I => \pid_alt.error_p_reg_esr_RNI0B681Z0Z_18\
        );

    \I__1880\ : InMux
    port map (
            O => \N__15851\,
            I => \pid_alt.un1_pid_prereg_0_cry_18\
        );

    \I__1879\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15845\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__15845\,
            I => \N__15842\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__15842\,
            I => \N__15839\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__15839\,
            I => \pid_alt.error_p_reg_esr_RNIIU781Z0Z_19\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__15836\,
            I => \N__15833\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15833\,
            I => \N__15830\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15830\,
            I => \N__15827\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__15827\,
            I => \N__15824\
        );

    \I__1871\ : Span4Mux_v
    port map (
            O => \N__15824\,
            I => \N__15821\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__15821\,
            I => \pid_alt.error_p_reg_esr_RNIH63KZ0Z_19\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15818\,
            I => \pid_alt.un1_pid_prereg_0_cry_19\
        );

    \I__1868\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__15809\,
            I => \pid_alt.error_p_reg_esr_RNI2G981Z0Z_20\
        );

    \I__1865\ : InMux
    port map (
            O => \N__15806\,
            I => \pid_alt.un1_pid_prereg_0_cry_20\
        );

    \I__1864\ : InMux
    port map (
            O => \N__15803\,
            I => \pid_alt.un1_pid_prereg_0_cry_21\
        );

    \I__1863\ : InMux
    port map (
            O => \N__15800\,
            I => \bfn_2_18_0_\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__15794\,
            I => \N__15791\
        );

    \I__1860\ : Odrv12
    port map (
            O => \N__15791\,
            I => \pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15788\,
            I => \pid_alt.un1_pid_prereg_0_cry_7\
        );

    \I__1858\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15782\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__15779\,
            I => \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__1854\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__15770\,
            I => \N__15767\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__15764\,
            I => \N__15761\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__15761\,
            I => \pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9\
        );

    \I__1849\ : InMux
    port map (
            O => \N__15758\,
            I => \pid_alt.un1_pid_prereg_0_cry_8\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__15755\,
            I => \N__15751\
        );

    \I__1847\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15748\
        );

    \I__1846\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15745\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15742\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15739\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__15742\,
            I => \N__15736\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__15739\,
            I => \N__15733\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__15736\,
            I => \N__15730\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__15733\,
            I => \pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__15730\,
            I => \pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__15725\,
            I => \N__15722\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15719\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15716\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__15713\,
            I => \pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15710\,
            I => \pid_alt.un1_pid_prereg_0_cry_9\
        );

    \I__1832\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15704\,
            I => \N__15701\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__15701\,
            I => \N__15697\
        );

    \I__1829\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15694\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__15694\,
            I => \pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__15691\,
            I => \pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__1824\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__15680\,
            I => \N__15677\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__15671\,
            I => \pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11\
        );

    \I__1819\ : InMux
    port map (
            O => \N__15668\,
            I => \pid_alt.un1_pid_prereg_0_cry_10\
        );

    \I__1818\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__15653\,
            I => \pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \N__15647\
        );

    \I__1812\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15644\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15644\,
            I => \N__15641\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__15638\,
            I => \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11\
        );

    \I__1808\ : InMux
    port map (
            O => \N__15635\,
            I => \pid_alt.un1_pid_prereg_0_cry_11\
        );

    \I__1807\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__15620\,
            I => \N__15617\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__15617\,
            I => \pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__15614\,
            I => \N__15610\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__15613\,
            I => \N__15607\
        );

    \I__1799\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15604\
        );

    \I__1798\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15601\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__15604\,
            I => \N__15598\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__15601\,
            I => \N__15595\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__15598\,
            I => \N__15592\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__15595\,
            I => \N__15587\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__15592\,
            I => \N__15587\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__15587\,
            I => \pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12\
        );

    \I__1791\ : InMux
    port map (
            O => \N__15584\,
            I => \pid_alt.un1_pid_prereg_0_cry_12\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15578\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__15578\,
            I => \N__15575\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__15572\,
            I => \N__15569\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__15569\,
            I => \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__1784\ : InMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__15560\,
            I => \N__15557\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__15554\,
            I => \N__15551\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__15548\,
            I => \pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13\
        );

    \I__1778\ : InMux
    port map (
            O => \N__15545\,
            I => \pid_alt.un1_pid_prereg_0_cry_13\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \N__15539\
        );

    \I__1776\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15536\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__15536\,
            I => \N__15532\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15535\,
            I => \N__15529\
        );

    \I__1773\ : Span4Mux_h
    port map (
            O => \N__15532\,
            I => \N__15524\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15529\,
            I => \N__15524\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__15515\,
            I => \pid_alt.error_p_regZ0Z_0\
        );

    \I__1767\ : InMux
    port map (
            O => \N__15512\,
            I => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\
        );

    \I__1766\ : InMux
    port map (
            O => \N__15509\,
            I => \pid_alt.un1_pid_prereg_0_cry_0\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15503\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__15503\,
            I => \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15494\,
            I => \pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2\
        );

    \I__1760\ : InMux
    port map (
            O => \N__15491\,
            I => \pid_alt.un1_pid_prereg_0_cry_1\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__1758\ : InMux
    port map (
            O => \N__15485\,
            I => \N__15481\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__15481\,
            I => \pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__15478\,
            I => \pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \N__15470\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15464\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__15464\,
            I => \pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3\
        );

    \I__1750\ : InMux
    port map (
            O => \N__15461\,
            I => \pid_alt.un1_pid_prereg_0_cry_2\
        );

    \I__1749\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__15452\,
            I => \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__1745\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__15437\,
            I => \pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4\
        );

    \I__1741\ : InMux
    port map (
            O => \N__15434\,
            I => \pid_alt.un1_pid_prereg_0_cry_3\
        );

    \I__1740\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__15422\,
            I => \N__15419\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__15419\,
            I => \pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15410\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__15410\,
            I => \N__15406\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15397\
        );

    \I__1729\ : Span4Mux_v
    port map (
            O => \N__15400\,
            I => \N__15394\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15397\,
            I => \N__15391\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__15394\,
            I => \pid_alt.error_p_reg_esr_RNI91H61Z0Z_4\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__15391\,
            I => \pid_alt.error_p_reg_esr_RNI91H61Z0Z_4\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15386\,
            I => \pid_alt.un1_pid_prereg_0_cry_4\
        );

    \I__1724\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15380\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__15377\,
            I => \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__15368\,
            I => \pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6\
        );

    \I__1718\ : InMux
    port map (
            O => \N__15365\,
            I => \pid_alt.un1_pid_prereg_0_cry_5\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15359\,
            I => \N__15355\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15352\
        );

    \I__1714\ : Span4Mux_s2_h
    port map (
            O => \N__15355\,
            I => \N__15349\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__15349\,
            I => \N__15342\
        );

    \I__1711\ : Span4Mux_s2_h
    port map (
            O => \N__15346\,
            I => \N__15339\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15336\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__15342\,
            I => drone_altitude_0
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__15339\,
            I => drone_altitude_0
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15336\,
            I => drone_altitude_0
        );

    \I__1706\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15314\
        );

    \I__1705\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15314\
        );

    \I__1704\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15314\
        );

    \I__1703\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15314\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15314\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__15314\,
            I => \N__15310\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__1699\ : Span4Mux_s3_h
    port map (
            O => \N__15310\,
            I => \N__15301\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__15307\,
            I => \N__15298\
        );

    \I__1697\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15293\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15293\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15290\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__15301\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\
        );

    \I__1693\ : Odrv12
    port map (
            O => \N__15298\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__15293\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__15290\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15278\,
            I => \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__15275\,
            I => \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15265\
        );

    \I__1685\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15262\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__15265\,
            I => \N__15255\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__15262\,
            I => \N__15255\
        );

    \I__1682\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15250\
        );

    \I__1681\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15250\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__15255\,
            I => \pid_alt.N_9_0\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__15250\,
            I => \pid_alt.N_9_0\
        );

    \I__1678\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__15239\,
            I => \pid_alt.m21_e_9\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__15236\,
            I => \pid_alt.N_9_0_cascade_\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__15227\,
            I => \pid_alt.m21_e_10\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_\
        );

    \I__1670\ : SRMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__15218\,
            I => \N__15213\
        );

    \I__1668\ : SRMux
    port map (
            O => \N__15217\,
            I => \N__15209\
        );

    \I__1667\ : SRMux
    port map (
            O => \N__15216\,
            I => \N__15205\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__15213\,
            I => \N__15202\
        );

    \I__1665\ : SRMux
    port map (
            O => \N__15212\,
            I => \N__15199\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__15209\,
            I => \N__15196\
        );

    \I__1663\ : SRMux
    port map (
            O => \N__15208\,
            I => \N__15193\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15205\,
            I => \N__15190\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__15202\,
            I => \N__15185\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15185\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__15196\,
            I => \N__15180\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15180\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__15190\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__15185\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__15180\,
            I => \pid_alt.un1_reset_1_0_i\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \pid_alt.un1_reset_1_0_i_cascade_\
        );

    \I__1653\ : CEMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15163\
        );

    \I__1651\ : CEMux
    port map (
            O => \N__15166\,
            I => \N__15160\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__15163\,
            I => \N__15154\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15160\,
            I => \N__15154\
        );

    \I__1648\ : CEMux
    port map (
            O => \N__15159\,
            I => \N__15151\
        );

    \I__1647\ : Span4Mux_h
    port map (
            O => \N__15154\,
            I => \N__15148\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__15151\,
            I => \N__15143\
        );

    \I__1645\ : Span4Mux_s1_h
    port map (
            O => \N__15148\,
            I => \N__15143\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__15143\,
            I => \pid_alt.N_60_i_0\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15140\,
            I => \scaler_2.un3_source_data_0_cry_1\
        );

    \I__1642\ : InMux
    port map (
            O => \N__15137\,
            I => \scaler_2.un3_source_data_0_cry_2\
        );

    \I__1641\ : InMux
    port map (
            O => \N__15134\,
            I => \scaler_2.un3_source_data_0_cry_3\
        );

    \I__1640\ : InMux
    port map (
            O => \N__15131\,
            I => \scaler_2.un3_source_data_0_cry_4\
        );

    \I__1639\ : InMux
    port map (
            O => \N__15128\,
            I => \scaler_2.un3_source_data_0_cry_5\
        );

    \I__1638\ : InMux
    port map (
            O => \N__15125\,
            I => \scaler_2.un3_source_data_0_cry_6\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15122\,
            I => \bfn_2_15_0_\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15119\,
            I => \scaler_2.un3_source_data_0_cry_8\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15106\
        );

    \I__1632\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15103\
        );

    \I__1631\ : Span4Mux_s3_h
    port map (
            O => \N__15106\,
            I => \N__15100\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__15103\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__15100\,
            I => \pid_alt.drone_altitude_i_0\
        );

    \I__1628\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15089\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15089\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__15089\,
            I => \N__15086\
        );

    \I__1625\ : Span4Mux_s2_h
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__15083\,
            I => \pid_alt.m35_e_2\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__15080\,
            I => \pid_alt.m35_e_2_cascade_\
        );

    \I__1622\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15074\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__15068\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__15065\,
            I => \N__15061\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__15064\,
            I => \N__15058\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15053\
        );

    \I__1615\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15053\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__15050\,
            I => \N__15046\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15043\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__15046\,
            I => \pid_alt.m35_e_3\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__15043\,
            I => \pid_alt.m35_e_3\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__15038\,
            I => \pid_alt.m21_e_2_cascade_\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \pid_alt.m21_e_0_cascade_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__15029\,
            I => \pid_alt.m21_e_8\
        );

    \I__1605\ : InMux
    port map (
            O => \N__15026\,
            I => \scaler_2.un3_source_data_0_cry_0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__15020\,
            I => \N__15016\
        );

    \I__1602\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15013\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__15010\,
            I => \N__15002\
        );

    \I__1598\ : Span4Mux_s1_h
    port map (
            O => \N__15007\,
            I => \N__15002\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__15002\,
            I => \pid_alt.error_8\
        );

    \I__1596\ : InMux
    port map (
            O => \N__14999\,
            I => \bfn_2_12_0_\
        );

    \I__1595\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14989\
        );

    \I__1593\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14986\
        );

    \I__1592\ : Span4Mux_v
    port map (
            O => \N__14989\,
            I => \N__14983\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__14986\,
            I => \N__14980\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__14983\,
            I => \N__14975\
        );

    \I__1589\ : Span4Mux_s1_h
    port map (
            O => \N__14980\,
            I => \N__14975\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__14975\,
            I => \pid_alt.error_9\
        );

    \I__1587\ : InMux
    port map (
            O => \N__14972\,
            I => \pid_alt.error_cry_8\
        );

    \I__1586\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14962\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__14962\,
            I => \N__14956\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__14956\,
            I => \N__14948\
        );

    \I__1580\ : Span4Mux_s1_h
    port map (
            O => \N__14953\,
            I => \N__14948\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__14948\,
            I => \pid_alt.error_10\
        );

    \I__1578\ : InMux
    port map (
            O => \N__14945\,
            I => \pid_alt.error_cry_9\
        );

    \I__1577\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14939\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14939\,
            I => \N__14936\
        );

    \I__1575\ : Span4Mux_v
    port map (
            O => \N__14936\,
            I => \N__14932\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__14932\,
            I => \N__14924\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__14929\,
            I => \N__14924\
        );

    \I__1571\ : Span4Mux_s1_h
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__14921\,
            I => \pid_alt.error_11\
        );

    \I__1569\ : InMux
    port map (
            O => \N__14918\,
            I => \pid_alt.error_cry_10\
        );

    \I__1568\ : InMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__14909\,
            I => \N__14905\
        );

    \I__1565\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14902\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__14905\,
            I => \N__14897\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__14902\,
            I => \N__14897\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__14897\,
            I => \pid_alt.error_12\
        );

    \I__1561\ : InMux
    port map (
            O => \N__14894\,
            I => \pid_alt.error_cry_11\
        );

    \I__1560\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__14885\,
            I => \N__14881\
        );

    \I__1557\ : InMux
    port map (
            O => \N__14884\,
            I => \N__14878\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__14881\,
            I => \N__14873\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14873\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__14873\,
            I => \pid_alt.error_13\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14870\,
            I => \pid_alt.error_cry_12\
        );

    \I__1552\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__14861\,
            I => \N__14857\
        );

    \I__1549\ : InMux
    port map (
            O => \N__14860\,
            I => \N__14854\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__14857\,
            I => \N__14849\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__14854\,
            I => \N__14849\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__14849\,
            I => \pid_alt.error_14\
        );

    \I__1545\ : InMux
    port map (
            O => \N__14846\,
            I => \pid_alt.error_cry_13\
        );

    \I__1544\ : InMux
    port map (
            O => \N__14843\,
            I => \pid_alt.error_cry_14\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__14834\,
            I => \N__14830\
        );

    \I__1540\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14827\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__14830\,
            I => \N__14822\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__14827\,
            I => \N__14822\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__14822\,
            I => \pid_alt.error_15\
        );

    \I__1536\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14813\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14818\,
            I => \N__14813\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14810\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__14807\,
            I => \pid_alt.error_p_regZ0Z_9\
        );

    \I__1531\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14800\
        );

    \I__1530\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14797\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__14800\,
            I => \N__14794\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__1527\ : Span4Mux_s2_h
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__1526\ : Span4Mux_s3_h
    port map (
            O => \N__14791\,
            I => \N__14785\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__14788\,
            I => \pid_alt.error_1\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__14785\,
            I => \pid_alt.error_1\
        );

    \I__1523\ : InMux
    port map (
            O => \N__14780\,
            I => \pid_alt.error_cry_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14773\
        );

    \I__1521\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14770\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__14773\,
            I => \N__14767\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__14770\,
            I => \N__14764\
        );

    \I__1518\ : Span4Mux_s3_h
    port map (
            O => \N__14767\,
            I => \N__14761\
        );

    \I__1517\ : Span4Mux_s2_h
    port map (
            O => \N__14764\,
            I => \N__14758\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__14761\,
            I => \pid_alt.error_2\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__14758\,
            I => \pid_alt.error_2\
        );

    \I__1514\ : InMux
    port map (
            O => \N__14753\,
            I => \pid_alt.error_cry_1\
        );

    \I__1513\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14746\
        );

    \I__1512\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14743\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14740\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__14743\,
            I => \N__14737\
        );

    \I__1509\ : Span4Mux_s2_h
    port map (
            O => \N__14740\,
            I => \N__14734\
        );

    \I__1508\ : Span4Mux_s2_h
    port map (
            O => \N__14737\,
            I => \N__14731\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__14734\,
            I => \pid_alt.error_3\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__14731\,
            I => \pid_alt.error_3\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14726\,
            I => \pid_alt.error_cry_2\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14719\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14716\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__14719\,
            I => \N__14713\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__14716\,
            I => \N__14710\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__14713\,
            I => \N__14707\
        );

    \I__1499\ : Span4Mux_s3_h
    port map (
            O => \N__14710\,
            I => \N__14704\
        );

    \I__1498\ : Span4Mux_s0_h
    port map (
            O => \N__14707\,
            I => \N__14701\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__14704\,
            I => \pid_alt.error_4\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__14701\,
            I => \pid_alt.error_4\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14696\,
            I => \pid_alt.error_cry_3\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14689\
        );

    \I__1493\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14686\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14689\,
            I => \N__14683\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__14686\,
            I => \N__14680\
        );

    \I__1490\ : Span4Mux_s2_h
    port map (
            O => \N__14683\,
            I => \N__14677\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__14680\,
            I => \N__14674\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__14677\,
            I => \pid_alt.error_5\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__14674\,
            I => \pid_alt.error_5\
        );

    \I__1486\ : InMux
    port map (
            O => \N__14669\,
            I => \pid_alt.error_cry_4\
        );

    \I__1485\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14663\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14659\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14656\
        );

    \I__1482\ : Span4Mux_s1_h
    port map (
            O => \N__14659\,
            I => \N__14653\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14656\,
            I => \N__14650\
        );

    \I__1480\ : Span4Mux_v
    port map (
            O => \N__14653\,
            I => \N__14647\
        );

    \I__1479\ : Span4Mux_s2_h
    port map (
            O => \N__14650\,
            I => \N__14644\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__14647\,
            I => \pid_alt.error_6\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__14644\,
            I => \pid_alt.error_6\
        );

    \I__1476\ : InMux
    port map (
            O => \N__14639\,
            I => \pid_alt.error_cry_5\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__14633\,
            I => \N__14629\
        );

    \I__1473\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14626\
        );

    \I__1472\ : Span4Mux_s1_h
    port map (
            O => \N__14629\,
            I => \N__14623\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__14626\,
            I => \N__14620\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__14623\,
            I => \N__14617\
        );

    \I__1469\ : Span4Mux_s2_h
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__14617\,
            I => \pid_alt.error_7\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__14614\,
            I => \pid_alt.error_7\
        );

    \I__1466\ : InMux
    port map (
            O => \N__14609\,
            I => \pid_alt.error_cry_6\
        );

    \I__1465\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__1462\ : Span4Mux_s1_h
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__14594\,
            I => alt_ki_2
        );

    \I__1460\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14588\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__1458\ : Span4Mux_s3_h
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__14582\,
            I => alt_ki_3
        );

    \I__1456\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14576\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__1454\ : Span4Mux_s3_h
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__14570\,
            I => alt_ki_5
        );

    \I__1452\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14564\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__14564\,
            I => \N__14561\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__14561\,
            I => \N__14558\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__14558\,
            I => alt_ki_6
        );

    \I__1448\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14552\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__14552\,
            I => \N__14549\
        );

    \I__1446\ : Span4Mux_h
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__14546\,
            I => \pid_alt.O_12\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14537\
        );

    \I__1443\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14537\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__14537\,
            I => \N__14534\
        );

    \I__1441\ : Span4Mux_v
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__14531\,
            I => \pid_alt.error_p_regZ0Z_8\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__14528\,
            I => \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__14516\,
            I => \pid_alt.O_13\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__14510\,
            I => \N__14507\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__14507\,
            I => \N__14504\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__14504\,
            I => \pid_alt.O_0_8\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14495\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14495\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__14495\,
            I => \N__14492\
        );

    \I__1427\ : Sp12to4
    port map (
            O => \N__14492\,
            I => \N__14489\
        );

    \I__1426\ : Span12Mux_v
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__1425\ : Odrv12
    port map (
            O => \N__14486\,
            I => \pid_alt.error_p_regZ0Z_4\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14480\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__14480\,
            I => \N__14477\
        );

    \I__1422\ : Span4Mux_s3_h
    port map (
            O => \N__14477\,
            I => \N__14474\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__14474\,
            I => alt_kp_2
        );

    \I__1420\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__14468\,
            I => \N__14465\
        );

    \I__1418\ : Span4Mux_s2_h
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__14462\,
            I => alt_ki_4
        );

    \I__1416\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__1414\ : Span12Mux_s2_h
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__1413\ : Odrv12
    port map (
            O => \N__14450\,
            I => alt_ki_1
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__14447\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__14444\,
            I => \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\
        );

    \I__1410\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__14438\,
            I => \ppm_encoder_1.un2_throttle_iv_0_9\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14430\
        );

    \I__1407\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14425\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14425\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__14430\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__14425\,
            I => \ppm_encoder_1.elevatorZ0Z_9\
        );

    \I__1403\ : InMux
    port map (
            O => \N__14420\,
            I => \N__14417\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__1401\ : Odrv12
    port map (
            O => \N__14414\,
            I => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14403\
        );

    \I__1398\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14400\
        );

    \I__1397\ : InMux
    port map (
            O => \N__14406\,
            I => \N__14397\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__14403\,
            I => \N__14392\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__14400\,
            I => \N__14392\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__14397\,
            I => throttle_command_9
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__14392\,
            I => throttle_command_9
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14379\
        );

    \I__1390\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14374\
        );

    \I__1389\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14374\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__14379\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__14374\,
            I => \ppm_encoder_1.throttleZ0Z_9\
        );

    \I__1386\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14364\
        );

    \I__1385\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14359\
        );

    \I__1384\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14359\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__14364\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14359\,
            I => \ppm_encoder_1.rudderZ0Z_9\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__14354\,
            I => \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\
        );

    \I__1380\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14348\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__14348\,
            I => \ppm_encoder_1.un2_throttle_iv_0_10\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14341\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14338\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14341\,
            I => \N__14335\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__14338\,
            I => \N__14332\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__14335\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__14332\,
            I => \ppm_encoder_1.throttleZ0Z_14\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__14327\,
            I => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\
        );

    \I__1371\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14321\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__14321\,
            I => \ppm_encoder_1.un2_throttle_iv_1_14\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__14318\,
            I => \ppm_encoder_1.un1_init_pulses_10_0_cascade_\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__14315\,
            I => \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14312\,
            I => \ppm_encoder_1.un1_throttle_cry_13\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__14309\,
            I => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \N__14301\
        );

    \I__1364\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14298\
        );

    \I__1363\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14295\
        );

    \I__1362\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14292\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14287\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__14295\,
            I => \N__14287\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14292\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__14287\,
            I => \ppm_encoder_1.throttleZ0Z_5\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__14282\,
            I => \ppm_encoder_1.N_297_cascade_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14276\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__1354\ : Span4Mux_v
    port map (
            O => \N__14273\,
            I => \N__14270\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__14270\,
            I => scaler_2_data_5
        );

    \I__1352\ : InMux
    port map (
            O => \N__14267\,
            I => \ppm_encoder_1.un1_throttle_cry_4\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14259\
        );

    \I__1350\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14256\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14253\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14250\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__14256\,
            I => throttle_command_6
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__14253\,
            I => throttle_command_6
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__14250\,
            I => throttle_command_6
        );

    \I__1344\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__14240\,
            I => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14237\,
            I => \ppm_encoder_1.un1_throttle_cry_5\
        );

    \I__1341\ : InMux
    port map (
            O => \N__14234\,
            I => \ppm_encoder_1.un1_throttle_cry_6\
        );

    \I__1340\ : InMux
    port map (
            O => \N__14231\,
            I => \bfn_1_23_0_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14228\,
            I => \ppm_encoder_1.un1_throttle_cry_8\
        );

    \I__1338\ : InMux
    port map (
            O => \N__14225\,
            I => \ppm_encoder_1.un1_throttle_cry_9\
        );

    \I__1337\ : InMux
    port map (
            O => \N__14222\,
            I => \ppm_encoder_1.un1_throttle_cry_10\
        );

    \I__1336\ : InMux
    port map (
            O => \N__14219\,
            I => \ppm_encoder_1.un1_throttle_cry_11\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14216\,
            I => \ppm_encoder_1.un1_throttle_cry_12\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14213\,
            I => \ppm_encoder_1.un1_throttle_cry_0\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14210\,
            I => \ppm_encoder_1.un1_throttle_cry_1\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14207\,
            I => \ppm_encoder_1.un1_throttle_cry_2\
        );

    \I__1331\ : InMux
    port map (
            O => \N__14204\,
            I => \ppm_encoder_1.un1_throttle_cry_3\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14201\,
            I => \N__14198\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__14198\,
            I => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14188\
        );

    \I__1326\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14185\
        );

    \I__1325\ : Odrv12
    port map (
            O => \N__14188\,
            I => \pid_alt.error_p_regZ0Z_5\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__14185\,
            I => \pid_alt.error_p_regZ0Z_5\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__14180\,
            I => \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__14177\,
            I => \N__14174\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14169\
        );

    \I__1320\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14166\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14163\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__14169\,
            I => \N__14158\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__14166\,
            I => \N__14158\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__14163\,
            I => \N__14155\
        );

    \I__1315\ : Span12Mux_v
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__1314\ : Span4Mux_v
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__14152\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__1312\ : Odrv4
    port map (
            O => \N__14149\,
            I => \pid_alt.error_p_regZ0Z_19\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14141\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__1309\ : Span12Mux_v
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__14135\,
            I => alt_ki_0
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \pid_alt.N_37_cascade_\
        );

    \I__1306\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14122\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14117\
        );

    \I__1304\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14117\
        );

    \I__1303\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14114\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14111\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__14122\,
            I => \pid_alt.N_62_mux\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__14117\,
            I => \pid_alt.N_62_mux\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14114\,
            I => \pid_alt.N_62_mux\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__14111\,
            I => \pid_alt.N_62_mux\
        );

    \I__1297\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14097\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14092\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14092\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__14097\,
            I => \pid_alt.N_37\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__14092\,
            I => \pid_alt.N_37\
        );

    \I__1292\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14081\
        );

    \I__1291\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14081\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__1289\ : Odrv12
    port map (
            O => \N__14078\,
            I => \pid_alt.error_p_regZ0Z_1\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__14075\,
            I => \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_\
        );

    \I__1287\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14066\
        );

    \I__1286\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14066\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__14066\,
            I => \N__14063\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__1283\ : Sp12to4
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__14057\,
            I => \pid_alt.error_p_regZ0Z_2\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__14054\,
            I => \N__14051\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14048\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__1278\ : Sp12to4
    port map (
            O => \N__14045\,
            I => \N__14040\
        );

    \I__1277\ : InMux
    port map (
            O => \N__14044\,
            I => \N__14035\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14043\,
            I => \N__14035\
        );

    \I__1275\ : Span12Mux_v
    port map (
            O => \N__14040\,
            I => \N__14030\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__14035\,
            I => \N__14030\
        );

    \I__1273\ : Odrv12
    port map (
            O => \N__14030\,
            I => \pid_alt.error_p_regZ0Z_17\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__14027\,
            I => \pid_alt.N_62_mux_cascade_\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__14024\,
            I => \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_\
        );

    \I__1270\ : InMux
    port map (
            O => \N__14021\,
            I => \N__14015\
        );

    \I__1269\ : InMux
    port map (
            O => \N__14020\,
            I => \N__14015\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__14006\,
            I => \pid_alt.error_p_regZ0Z_3\
        );

    \I__1264\ : InMux
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__14000\,
            I => \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5\
        );

    \I__1262\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__13991\,
            I => \pid_alt.O_9\
        );

    \I__1259\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__13982\,
            I => \pid_alt.O_8\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__13979\,
            I => \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13973\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__13973\,
            I => \pid_alt.O_16\
        );

    \I__1253\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13964\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13964\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__1250\ : Span4Mux_v
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__13958\,
            I => \pid_alt.error_p_regZ0Z_12\
        );

    \I__1248\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13952\,
            I => \pid_alt.O_14\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13943\
        );

    \I__1245\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13943\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__13940\,
            I => \pid_alt.error_p_regZ0Z_10\
        );

    \I__1242\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__13928\,
            I => \pid_alt.O_5\
        );

    \I__1238\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13919\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__13916\,
            I => \pid_alt.O_7\
        );

    \I__1234\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13910\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__13907\,
            I => \pid_alt.O_19\
        );

    \I__1231\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__13898\,
            I => \pid_alt.O_20\
        );

    \I__1228\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__13889\,
            I => \pid_alt.O_21\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__13880\,
            I => \pid_alt.O_22\
        );

    \I__1222\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__13874\,
            I => \pid_alt.O_6\
        );

    \I__1220\ : InMux
    port map (
            O => \N__13871\,
            I => \N__13868\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__13865\,
            I => \pid_alt.O_24\
        );

    \I__1217\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__13859\,
            I => \pid_alt.O_15\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__1214\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13847\
        );

    \I__1213\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13847\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__13844\,
            I => \N__13841\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__13841\,
            I => \pid_alt.error_p_regZ0Z_11\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__13838\,
            I => \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_\
        );

    \I__1208\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13829\
        );

    \I__1207\ : InMux
    port map (
            O => \N__13834\,
            I => \N__13829\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__13826\,
            I => \pid_alt.error_p_regZ0Z_13\
        );

    \I__1204\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13820\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__13820\,
            I => \N__13817\
        );

    \I__1202\ : Span4Mux_h
    port map (
            O => \N__13817\,
            I => \N__13814\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__13814\,
            I => \pid_alt.O_18\
        );

    \I__1200\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13804\
        );

    \I__1199\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__1198\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13801\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__13801\,
            I => \pid_alt.error_p_regZ0Z_14\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__13798\,
            I => \pid_alt.error_p_regZ0Z_14\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13790\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__13790\,
            I => \N__13787\
        );

    \I__1192\ : Span4Mux_h
    port map (
            O => \N__13787\,
            I => \N__13784\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__13784\,
            I => \pid_alt.O_23\
        );

    \I__1190\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13778\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__13778\,
            I => \pid_alt.O_4\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13772\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13769\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__13769\,
            I => \pid_alt.O_17\
        );

    \I__1185\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__13763\,
            I => \pid_alt.O_0_13\
        );

    \I__1183\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13757\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__13757\,
            I => \N__13754\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__13754\,
            I => \pid_alt.O_0_24\
        );

    \I__1180\ : InMux
    port map (
            O => \N__13751\,
            I => \N__13748\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__13748\,
            I => \pid_alt.O_0_19\
        );

    \I__1178\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13742\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__13742\,
            I => \pid_alt.O_0_20\
        );

    \I__1176\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__13736\,
            I => \pid_alt.O_0_18\
        );

    \I__1174\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__13730\,
            I => \pid_alt.O_0_9\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__13727\,
            I => \N__13722\
        );

    \I__1171\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13719\
        );

    \I__1170\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13714\
        );

    \I__1169\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13714\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__13719\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__13714\,
            I => \pid_alt.error_p_regZ0Z_15\
        );

    \I__1166\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__13703\,
            I => \pid_alt.O_0_17\
        );

    \I__1163\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13697\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__13697\,
            I => \pid_alt.O_0_15\
        );

    \I__1161\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__13688\,
            I => \pid_alt.O_0_16\
        );

    \I__1158\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13682\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__13682\,
            I => \pid_alt.O_0_5\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13676\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__13676\,
            I => \N__13673\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__13673\,
            I => \pid_alt.O_0_22\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__13667\,
            I => \pid_alt.O_0_4\
        );

    \I__1151\ : InMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__13661\,
            I => \pid_alt.O_0_10\
        );

    \I__1149\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__13655\,
            I => \pid_alt.O_0_23\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__13649\,
            I => \pid_alt.O_0_11\
        );

    \I__1145\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13643\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__13640\,
            I => \pid_alt.O_0_6\
        );

    \I__1142\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13634\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__13631\,
            I => \pid_alt.O_0_14\
        );

    \I__1139\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13625\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__13622\,
            I => \pid_alt.O_0_12\
        );

    \I__1136\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13616\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__13613\,
            I => \pid_alt.O_0_21\
        );

    \I__1133\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__13607\,
            I => \pid_alt.O_0_7\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_6\,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_pid_prereg_0_cry_14\,
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un3_source_data_0_cry_7\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_4.un2_source_data_0_cry_8\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un3_source_data_0_cry_7\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_3.un2_source_data_0_cry_8\,
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un3_source_data_0_cry_7\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \scaler_2.un2_source_data_0_cry_8\,
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_8\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \reset_module_System.count_1_cry_16\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_throttle_cry_7\,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_5_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_29_0_\
        );

    \IN_MUX_bfv_5_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_rudder_cry_13\,
            carryinitout => \bfn_5_30_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_elevator_cry_13\,
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_3_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_aileron_cry_13\,
            carryinitout => \bfn_3_22_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            carryinitout => \bfn_2_27_0_\
        );

    \IN_MUX_bfv_2_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_28_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_5_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.counter24_0_data_tmp_7\,
            carryinitout => \bfn_5_28_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pid_alt.error_cry_7\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_10_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_11_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_7\,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ppm_encoder_1.un1_counter_13_cry_15\,
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \dron_frame_decoder_1.un1_WDT_cry_7\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \Commands_frame_decoder.un1_WDT_cry_7\,
            carryinitout => \bfn_11_16_0_\
        );

    \reset_module_System.reset_RNITC69_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26141\,
            GLOBALBUFFEROUTPUT => \N_423_g\
        );

    \reset_module_System.reset_RNITC69\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__35079\,
            GLOBALBUFFEROUTPUT => reset_system_g
        );

    \pid_alt.state_RNICP2N1_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21494\,
            GLOBALBUFFEROUTPUT => \pid_alt.N_422_0_g\
        );

    \debug_CH3_20A_c_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__36377\,
            GLOBALBUFFEROUTPUT => \debug_CH3_20A_c_0_g\
        );

    \pid_alt.state_RNIH1EN_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34076\,
            GLOBALBUFFEROUTPUT => \pid_alt.state_0_g_0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25313\,
            GLOBALBUFFEROUTPUT => \ppm_encoder_1.N_320_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_2_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13646\,
            lcout => \pid_alt.error_p_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36167\,
            ce => \N__20312\,
            sr => \N__21582\
        );

    \pid_alt.error_p_reg_esr_10_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13637\,
            lcout => \pid_alt.error_p_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36166\,
            ce => \N__20311\,
            sr => \N__21581\
        );

    \pid_alt.error_p_reg_esr_8_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13628\,
            lcout => \pid_alt.error_p_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36166\,
            ce => \N__20311\,
            sr => \N__21581\
        );

    \pid_alt.error_p_reg_esr_17_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13619\,
            lcout => \pid_alt.error_p_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36166\,
            ce => \N__20311\,
            sr => \N__21581\
        );

    \pid_alt.error_p_reg_esr_3_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13610\,
            lcout => \pid_alt.error_p_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36166\,
            ce => \N__20311\,
            sr => \N__21581\
        );

    \pid_alt.error_p_reg_esr_13_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13709\,
            lcout => \pid_alt.error_p_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_11_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13700\,
            lcout => \pid_alt.error_p_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_12_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13694\,
            lcout => \pid_alt.error_p_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_1_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13685\,
            lcout => \pid_alt.error_p_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_18_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13679\,
            lcout => \pid_alt.error_p_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_0_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13670\,
            lcout => \pid_alt.error_p_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36165\,
            ce => \N__20310\,
            sr => \N__21580\
        );

    \pid_alt.error_p_reg_esr_6_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13664\,
            lcout => \pid_alt.error_p_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_19_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13658\,
            lcout => \pid_alt.error_p_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_7_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13652\,
            lcout => \pid_alt.error_p_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_9_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13766\,
            lcout => \pid_alt.error_p_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_20_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13760\,
            lcout => \pid_alt.error_p_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_15_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13751\,
            lcout => \pid_alt.error_p_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_16_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13745\,
            lcout => \pid_alt.error_p_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_14_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13739\,
            lcout => \pid_alt.error_p_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36163\,
            ce => \N__20308\,
            sr => \N__21578\
        );

    \pid_alt.error_p_reg_esr_RNIC74E2_5_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17377\,
            in1 => \N__17416\,
            in2 => \N__15416\,
            in3 => \N__14191\,
            lcout => \pid_alt.error_p_reg_esr_RNIC74E2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_5_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13733\,
            lcout => \pid_alt.error_p_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36161\,
            ce => \N__20307\,
            sr => \N__21577\
        );

    \pid_alt.error_p_reg_esr_RNIGQ581_14_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__13809\,
            in1 => \N__18370\,
            in2 => \N__13727\,
            in3 => \N__18143\,
            lcout => \pid_alt.error_p_reg_esr_RNIGQ581Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI9U2K_15_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18371\,
            lcout => \pid_alt.error_p_reg_esr_RNI9U2KZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIKU581_15_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__13726\,
            in1 => \N__18489\,
            in2 => \N__18381\,
            in3 => \N__18525\,
            lcout => \pid_alt.error_p_reg_esr_RNIKU581Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI6JDH1_13_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13834\,
            in1 => \N__17710\,
            in2 => \N__15613\,
            in3 => \N__17746\,
            lcout => \pid_alt.error_p_reg_esr_RNI6JDH1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI7S2K_0_14_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18133\,
            in2 => \_gnd_net_\,
            in3 => \N__13810\,
            lcout => \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14\,
            ltout => \pid_alt.error_p_reg_esr_RNI7S2K_0Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI0R7B1_13_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__17747\,
            in1 => \N__17709\,
            in2 => \N__13838\,
            in3 => \N__13835\,
            lcout => \pid_alt.error_p_reg_esr_RNI0R7B1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_14_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13823\,
            lcout => \pid_alt.error_i_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36157\,
            ce => \N__20306\,
            sr => \N__21576\
        );

    \pid_alt.error_p_reg_esr_RNI7S2K_14_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13811\,
            in1 => \_gnd_net_\,
            in2 => \N__18144\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.error_p_reg_esr_RNI7S2KZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIH63K_19_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18585\,
            in2 => \_gnd_net_\,
            in3 => \N__14172\,
            lcout => \pid_alt.error_p_reg_esr_RNIH63KZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_19_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13793\,
            lcout => \pid_alt.error_i_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36154\,
            ce => \N__20305\,
            sr => \N__21575\
        );

    \pid_alt.error_i_reg_esr_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13781\,
            lcout => \pid_alt.error_i_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_13_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13775\,
            lcout => \pid_alt.error_i_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_15_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13913\,
            lcout => \pid_alt.error_i_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_16_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13904\,
            lcout => \pid_alt.error_i_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_17_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13895\,
            lcout => \pid_alt.error_i_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_18_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13886\,
            lcout => \pid_alt.error_i_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_2_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13877\,
            lcout => \pid_alt.error_i_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_i_reg_esr_20_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13871\,
            lcout => \pid_alt.error_i_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36151\,
            ce => \N__20304\,
            sr => \N__21574\
        );

    \pid_alt.error_p_reg_esr_RNIHVGK1_11_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__15700\,
            in1 => \N__13852\,
            in2 => \N__17893\,
            in3 => \N__17907\,
            lcout => \pid_alt.error_p_reg_esr_RNIHVGK1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_11_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13862\,
            lcout => \pid_alt.error_i_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36147\,
            ce => \N__20302\,
            sr => \N__21572\
        );

    \pid_alt.error_p_reg_esr_RNIAH8Q_11_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17908\,
            in1 => \_gnd_net_\,
            in2 => \N__13856\,
            in3 => \N__17888\,
            lcout => \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11\,
            ltout => \pid_alt.error_p_reg_esr_RNIAH8QZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIN5HK1_12_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__13969\,
            in1 => \N__17807\,
            in2 => \N__13979\,
            in3 => \N__17826\,
            lcout => \pid_alt.error_p_reg_esr_RNIN5HK1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_12_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13976\,
            lcout => \pid_alt.error_i_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36147\,
            ce => \N__20302\,
            sr => \N__21572\
        );

    \pid_alt.error_p_reg_esr_RNIDK8Q_12_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__13970\,
            in1 => \N__17808\,
            in2 => \_gnd_net_\,
            in3 => \N__17827\,
            lcout => \pid_alt.error_p_reg_esr_RNIDK8QZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIM0S12_10_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17966\,
            in1 => \N__17985\,
            in2 => \N__15755\,
            in3 => \N__13948\,
            lcout => \pid_alt.error_p_reg_esr_RNIM0S12Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_10_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13955\,
            lcout => \pid_alt.error_i_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36144\,
            ce => \N__20301\,
            sr => \N__21571\
        );

    \pid_alt.error_p_reg_esr_RNI7E8Q_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__17967\,
            in1 => \N__13949\,
            in2 => \_gnd_net_\,
            in3 => \N__17986\,
            lcout => \pid_alt.error_p_reg_esr_RNI7E8QZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIO2681_16_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__18860\,
            in1 => \N__14044\,
            in2 => \N__18498\,
            in3 => \N__18539\,
            lcout => \pid_alt.error_p_reg_esr_RNIO2681Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNID23K_17_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14043\,
            lcout => \pid_alt.error_p_reg_esr_RNID23KZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_1_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13937\,
            lcout => \pid_alt.error_i_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36140\,
            ce => \N__20299\,
            sr => \N__21569\
        );

    \pid_alt.error_i_reg_esr_3_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13925\,
            lcout => \pid_alt.error_i_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36140\,
            ce => \N__20299\,
            sr => \N__21569\
        );

    \pid_alt.error_i_reg_esr_5_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13997\,
            lcout => \pid_alt.error_i_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36140\,
            ce => \N__20299\,
            sr => \N__21569\
        );

    \pid_alt.error_i_reg_esr_4_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13988\,
            lcout => \pid_alt.error_i_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36140\,
            ce => \N__20299\,
            sr => \N__21569\
        );

    \pid_alt.error_i_acumm_10_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__15325\,
            in1 => \N__23950\,
            in2 => \N__17971\,
            in3 => \N__17939\,
            lcout => \pid_alt.error_i_acummZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_11_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__23947\,
            in1 => \N__15328\,
            in2 => \N__17892\,
            in3 => \N__17858\,
            lcout => \pid_alt.error_i_acummZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_6_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__15326\,
            in1 => \N__23951\,
            in2 => \N__20397\,
            in3 => \N__17303\,
            lcout => \pid_alt.error_i_acummZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_9_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__23949\,
            in1 => \N__15329\,
            in2 => \N__18050\,
            in3 => \N__18014\,
            lcout => \pid_alt.error_i_acummZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_8_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__15327\,
            in1 => \N__23952\,
            in2 => \N__17225\,
            in3 => \N__17192\,
            lcout => \pid_alt.error_i_acummZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_12_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__17776\,
            in1 => \N__15269\,
            in2 => \N__17812\,
            in3 => \N__23953\,
            lcout => \pid_alt.error_i_acummZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_5_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__17344\,
            in2 => \N__17415\,
            in3 => \N__14125\,
            lcout => \pid_alt.error_i_acummZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36135\,
            ce => 'H',
            sr => \N__15216\
        );

    \pid_alt.error_i_acumm_esr_3_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__14126\,
            in1 => \N__14102\,
            in2 => \N__17470\,
            in3 => \N__17540\,
            lcout => \pid_alt.error_i_acummZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36131\,
            ce => \N__15170\,
            sr => \N__15217\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI6M6T3_10_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__15095\,
            in1 => \N__15261\,
            in2 => \N__15065\,
            in3 => \N__15305\,
            lcout => \pid_alt.N_62_mux\,
            ltout => \pid_alt.N_62_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_4_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100011101"
        )
    port map (
            in0 => \N__15306\,
            in1 => \N__17345\,
            in2 => \N__14027\,
            in3 => \N__17464\,
            lcout => \pid_alt.error_i_acummZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36131\,
            ce => \N__15170\,
            sr => \N__15217\
        );

    \pid_alt.error_p_reg_esr_RNI6UG61_3_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17587\,
            in1 => \_gnd_net_\,
            in2 => \N__17560\,
            in3 => \N__14021\,
            lcout => \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3\,
            ltout => \pid_alt.error_p_reg_esr_RNI6UG61Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIFV1D2_4_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14500\,
            in1 => \N__17490\,
            in2 => \N__14024\,
            in3 => \N__17511\,
            lcout => \pid_alt.error_p_reg_esr_RNIFV1D2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI91H61_4_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17512\,
            in1 => \_gnd_net_\,
            in2 => \N__17497\,
            in3 => \N__14501\,
            lcout => \pid_alt.error_p_reg_esr_RNI91H61Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI9P1D2_3_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14020\,
            in1 => \N__17553\,
            in2 => \N__15488\,
            in3 => \N__17586\,
            lcout => \pid_alt.error_p_reg_esr_RNI9P1D2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0_5_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15094\,
            in1 => \N__17343\,
            in2 => \N__15064\,
            in3 => \N__15260\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_1_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__17466\,
            in1 => \N__14128\,
            in2 => \N__17081\,
            in3 => \N__14100\,
            lcout => \pid_alt.error_i_acummZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36125\,
            ce => \N__15159\,
            sr => \N__15212\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNISKMM7_5_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15077\,
            in1 => \N__14003\,
            in2 => \_gnd_net_\,
            in3 => \N__15304\,
            lcout => \pid_alt.N_37\,
            ltout => \pid_alt.N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_0_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__18202\,
            in1 => \N__14127\,
            in2 => \N__14132\,
            in3 => \N__17465\,
            lcout => \pid_alt.error_i_acummZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36125\,
            ce => \N__15159\,
            sr => \N__15212\
        );

    \pid_alt.error_p_reg_esr_RNI0OG61_0_1_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17118\,
            in1 => \N__14086\,
            in2 => \_gnd_net_\,
            in3 => \N__17100\,
            lcout => \pid_alt.un1_pid_prereg_0_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_2_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__14129\,
            in1 => \N__14101\,
            in2 => \N__17471\,
            in3 => \N__17609\,
            lcout => \pid_alt.error_i_acummZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36125\,
            ce => \N__15159\,
            sr => \N__15212\
        );

    \pid_alt.error_p_reg_esr_RNI0OG61_1_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__17119\,
            in1 => \N__14087\,
            in2 => \_gnd_net_\,
            in3 => \N__17101\,
            lcout => \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1\,
            ltout => \pid_alt.error_p_reg_esr_RNI0OG61Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI3J1D2_2_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14071\,
            in1 => \N__17622\,
            in2 => \N__14075\,
            in3 => \N__17655\,
            lcout => \pid_alt.error_p_reg_esr_RNI3J1D2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI3RG61_2_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17656\,
            in1 => \_gnd_net_\,
            in2 => \N__17629\,
            in3 => \N__14072\,
            lcout => \pid_alt.error_p_reg_esr_RNI3RG61Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI2G981_20_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111000"
        )
    port map (
            in0 => \N__20789\,
            in1 => \N__20844\,
            in2 => \N__20799\,
            in3 => \N__20846\,
            lcout => \pid_alt.error_p_reg_esr_RNI2G981Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIS6681_17_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__18870\,
            in1 => \N__20581\,
            in2 => \N__14054\,
            in3 => \N__20620\,
            lcout => \pid_alt.error_p_reg_esr_RNIS6681Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIIU781_19_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20788\,
            in1 => \N__18597\,
            in2 => \N__14177\,
            in3 => \N__20845\,
            lcout => \pid_alt.error_p_reg_esr_RNIIU781Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI36J71_5_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__14195\,
            in1 => \N__17373\,
            in2 => \_gnd_net_\,
            in3 => \N__17411\,
            lcout => \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5\,
            ltout => \pid_alt.error_p_reg_esr_RNI36J71Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI9F6F2_6_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20434\,
            in1 => \N__20458\,
            in2 => \N__14180\,
            in3 => \N__20390\,
            lcout => \pid_alt.error_p_reg_esr_RNI9F6F2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI0B681_18_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__20621\,
            in1 => \N__14173\,
            in2 => \N__20585\,
            in3 => \N__18596\,
            lcout => \pid_alt.error_p_reg_esr_RNI0B681Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_0_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31493\,
            in2 => \_gnd_net_\,
            in3 => \N__21625\,
            lcout => alt_ki_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36115\,
            ce => \N__28049\,
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_5_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23780\,
            in1 => \N__23818\,
            in2 => \_gnd_net_\,
            in3 => \N__21041\,
            lcout => scaler_2_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36109\,
            ce => \N__29572\,
            sr => \N__36739\
        );

    \pid_alt.source_pid_1_10_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__18659\,
            in1 => \N__18802\,
            in2 => \N__21415\,
            in3 => \N__23939\,
            lcout => throttle_command_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => 'H',
            sr => \N__19260\
        );

    \pid_alt.source_pid_1_11_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111010000"
        )
    port map (
            in0 => \N__18803\,
            in1 => \N__18761\,
            in2 => \N__23954\,
            in3 => \N__16107\,
            lcout => throttle_command_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => 'H',
            sr => \N__19260\
        );

    \pid_alt.source_pid_1_7_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__18641\,
            in1 => \N__18805\,
            in2 => \N__16187\,
            in3 => \N__23940\,
            lcout => throttle_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => 'H',
            sr => \N__19260\
        );

    \pid_alt.source_pid_1_6_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111010000"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__18710\,
            in2 => \N__23955\,
            in3 => \N__14263\,
            lcout => throttle_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => 'H',
            sr => \N__19260\
        );

    \pid_alt.source_pid_1_9_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001001110"
        )
    port map (
            in0 => \N__23932\,
            in1 => \N__14406\,
            in2 => \N__18809\,
            in3 => \N__18737\,
            lcout => throttle_command_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36103\,
            ce => 'H',
            sr => \N__19260\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_14_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__24300\,
            in1 => \N__23089\,
            in2 => \_gnd_net_\,
            in3 => \N__30099\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_14_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29426\,
            in1 => \N__14345\,
            in2 => \_gnd_net_\,
            in3 => \N__24407\,
            lcout => \ppm_encoder_1.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_5_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__24972\,
            in1 => \N__15989\,
            in2 => \N__14306\,
            in3 => \N__14201\,
            lcout => \ppm_encoder_1.throttleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36096\,
            ce => 'H',
            sr => \N__36750\
        );

    \ppm_encoder_1.throttle_6_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__14243\,
            in1 => \N__14262\,
            in2 => \N__29329\,
            in3 => \N__24973\,
            lcout => \ppm_encoder_1.throttleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36096\,
            ce => 'H',
            sr => \N__36750\
        );

    \ppm_encoder_1.un1_throttle_cry_0_c_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_0_THRU_LUT4_0_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25069\,
            in2 => \N__28567\,
            in3 => \N__14213\,
            lcout => \ppm_encoder_1.un1_throttle_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_0\,
            carryout => \ppm_encoder_1.un1_throttle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_1_THRU_LUT4_0_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21322\,
            in2 => \_gnd_net_\,
            in3 => \N__14210\,
            lcout => \ppm_encoder_1.un1_throttle_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_1\,
            carryout => \ppm_encoder_1.un1_throttle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_2_THRU_LUT4_0_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25021\,
            in2 => \N__28568\,
            in3 => \N__14207\,
            lcout => \ppm_encoder_1.un1_throttle_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_2\,
            carryout => \ppm_encoder_1.un1_throttle_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_3_THRU_LUT4_0_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21811\,
            in2 => \_gnd_net_\,
            in3 => \N__14204\,
            lcout => \ppm_encoder_1.un1_throttle_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_3\,
            carryout => \ppm_encoder_1.un1_throttle_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_4_THRU_LUT4_0_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15985\,
            in2 => \_gnd_net_\,
            in3 => \N__14267\,
            lcout => \ppm_encoder_1.un1_throttle_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_4\,
            carryout => \ppm_encoder_1.un1_throttle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_5_THRU_LUT4_0_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14264\,
            in2 => \N__28569\,
            in3 => \N__14237\,
            lcout => \ppm_encoder_1.un1_throttle_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_5\,
            carryout => \ppm_encoder_1.un1_throttle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_6_THRU_LUT4_0_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16182\,
            in2 => \_gnd_net_\,
            in3 => \N__14234\,
            lcout => \ppm_encoder_1.un1_throttle_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_6\,
            carryout => \ppm_encoder_1.un1_throttle_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_7_THRU_LUT4_0_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21922\,
            in2 => \_gnd_net_\,
            in3 => \N__14231\,
            lcout => \ppm_encoder_1.un1_throttle_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => \ppm_encoder_1.un1_throttle_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_8_THRU_LUT4_0_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14407\,
            in2 => \_gnd_net_\,
            in3 => \N__14228\,
            lcout => \ppm_encoder_1.un1_throttle_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_8\,
            carryout => \ppm_encoder_1.un1_throttle_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_9_THRU_LUT4_0_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21411\,
            in2 => \_gnd_net_\,
            in3 => \N__14225\,
            lcout => \ppm_encoder_1.un1_throttle_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_9\,
            carryout => \ppm_encoder_1.un1_throttle_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_10_THRU_LUT4_0_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16108\,
            in2 => \_gnd_net_\,
            in3 => \N__14222\,
            lcout => \ppm_encoder_1.un1_throttle_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_10\,
            carryout => \ppm_encoder_1.un1_throttle_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_11_THRU_LUT4_0_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21685\,
            in2 => \_gnd_net_\,
            in3 => \N__14219\,
            lcout => \ppm_encoder_1.un1_throttle_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_11\,
            carryout => \ppm_encoder_1.un1_throttle_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_throttle_cry_12_THRU_LUT4_0_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21370\,
            in2 => \N__28535\,
            in3 => \N__14216\,
            lcout => \ppm_encoder_1.un1_throttle_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_throttle_cry_12\,
            carryout => \ppm_encoder_1.un1_throttle_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_14_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14312\,
            lcout => \ppm_encoder_1.throttleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36081\,
            ce => \N__27302\,
            sr => \N__36757\
        );

    \CONSTANT_ONE_LUT4_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNIV1OJ2_5_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__14304\,
            in1 => \N__27319\,
            in2 => \N__22361\,
            in3 => \N__22262\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNI4FIN5_5_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__16432\,
            in1 => \_gnd_net_\,
            in2 => \N__14309\,
            in3 => \N__16262\,
            lcout => \ppm_encoder_1.aileron_esr_RNI4FIN5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_5_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14305\,
            in1 => \N__16274\,
            in2 => \_gnd_net_\,
            in3 => \N__22500\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_5_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29237\,
            in2 => \N__14282\,
            in3 => \N__16286\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_5_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14279\,
            lcout => \ppm_encoder_1.aileronZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36072\,
            ce => \N__27294\,
            sr => \N__36759\
        );

    \ppm_encoder_1.elevator_esr_5_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29588\,
            lcout => \ppm_encoder_1.elevatorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36072\,
            ce => \N__27294\,
            sr => \N__36759\
        );

    \ppm_encoder_1.aileron_esr_RNIOVDS2_14_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__24403\,
            in1 => \N__19052\,
            in2 => \N__22125\,
            in3 => \N__22026\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIU0DH2_10_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__24160\,
            in1 => \N__24103\,
            in2 => \N__22130\,
            in3 => \N__22030\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI5GRT5_10_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19616\,
            in2 => \N__14354\,
            in3 => \N__14351\,
            lcout => \ppm_encoder_1.elevator_RNI5GRT5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIE2JI2_10_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__22606\,
            in1 => \N__25456\,
            in2 => \N__22264\,
            in3 => \N__22353\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_esr_RNI81QU2_14_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__22354\,
            in1 => \N__14344\,
            in2 => \N__25784\,
            in3 => \N__22256\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNITH3L6_14_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \N__16552\,
            in1 => \_gnd_net_\,
            in2 => \N__14327\,
            in3 => \N__14324\,
            lcout => \ppm_encoder_1.aileron_esr_RNITH3L6Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIN3352_0_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24514\,
            in2 => \N__19838\,
            in3 => \N__22252\,
            lcout => \ppm_encoder_1.throttle_RNIN3352Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_0_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101100011"
        )
    port map (
            in0 => \N__24515\,
            in1 => \N__19833\,
            in2 => \N__22265\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_0_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__23230\,
            in1 => \N__19664\,
            in2 => \N__14318\,
            in3 => \N__20121\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36062\,
            ce => 'H',
            sr => \N__36762\
        );

    \ppm_encoder_1.elevator_RNIEMVN2_9_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__14433\,
            in1 => \N__23421\,
            in2 => \N__22031\,
            in3 => \N__22129\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNITSI96_9_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__19577\,
            in1 => \_gnd_net_\,
            in2 => \N__14315\,
            in3 => \N__14441\,
            lcout => \ppm_encoder_1.throttle_RNITSI96Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIU7KK2_9_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__14382\,
            in1 => \N__14367\,
            in2 => \N__22360\,
            in3 => \N__22260\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_9_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29483\,
            in1 => \N__14383\,
            in2 => \_gnd_net_\,
            in3 => \N__14434\,
            lcout => \ppm_encoder_1.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_9_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011100100"
        )
    port map (
            in0 => \N__24991\,
            in1 => \N__14435\,
            in2 => \N__24467\,
            in3 => \N__28907\,
            lcout => \ppm_encoder_1.elevatorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36055\,
            ce => 'H',
            sr => \N__36766\
        );

    \ppm_encoder_1.throttle_9_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__24996\,
            in1 => \N__14420\,
            in2 => \N__14387\,
            in3 => \N__14411\,
            lcout => \ppm_encoder_1.throttleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36055\,
            ce => 'H',
            sr => \N__36766\
        );

    \ppm_encoder_1.aileron_9_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__19091\,
            in1 => \N__20915\,
            in2 => \N__25001\,
            in3 => \N__23422\,
            lcout => \ppm_encoder_1.aileronZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36055\,
            ce => 'H',
            sr => \N__36766\
        );

    \ppm_encoder_1.rudder_9_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__14368\,
            in1 => \N__24992\,
            in2 => \N__25559\,
            in3 => \N__26477\,
            lcout => \ppm_encoder_1.rudderZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36055\,
            ce => 'H',
            sr => \N__36766\
        );

    \ppm_encoder_1.init_pulses_9_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__20108\,
            in1 => \N__23237\,
            in2 => \N__16361\,
            in3 => \N__16709\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36048\,
            ce => 'H',
            sr => \N__36769\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_0_9_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19596\,
            in1 => \N__23059\,
            in2 => \_gnd_net_\,
            in3 => \N__30048\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_9_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19597\,
            in1 => \N__27957\,
            in2 => \N__30583\,
            in3 => \N__14369\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_0_5_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__30047\,
            in1 => \_gnd_net_\,
            in2 => \N__23085\,
            in3 => \N__20008\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIDQUS_5_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20007\,
            in1 => \N__23055\,
            in2 => \_gnd_net_\,
            in3 => \N__30046\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_5_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__27956\,
            in1 => \N__20009\,
            in2 => \N__27326\,
            in3 => \N__30575\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_0_8_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__24259\,
            in1 => \N__23060\,
            in2 => \_gnd_net_\,
            in3 => \N__30049\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUPKO2_13_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23288\,
            in1 => \N__24580\,
            in2 => \N__30089\,
            in3 => \N__19945\,
            lcout => \ppm_encoder_1.init_pulses_RNIUPKO2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_0_1_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23284\,
            in2 => \_gnd_net_\,
            in3 => \N__30051\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30052\,
            in1 => \_gnd_net_\,
            in2 => \N__23296\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_0_1_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30050\,
            lcout => \ppm_encoder_1.N_1014_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_17_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23236\,
            in1 => \N__20083\,
            in2 => \N__16472\,
            in3 => \N__16793\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36041\,
            ce => 'H',
            sr => \N__36771\
        );

    \ppm_encoder_1.init_pulses_14_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__20082\,
            in1 => \N__23235\,
            in2 => \N__16532\,
            in3 => \N__16832\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36041\,
            ce => 'H',
            sr => \N__36771\
        );

    \ppm_encoder_1.PPM_STATE_RNI78NT_0_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__25298\,
            in1 => \N__22417\,
            in2 => \N__22505\,
            in3 => \N__25362\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIRCE81_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__25397\,
            in1 => \_gnd_net_\,
            in2 => \N__14447\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_1\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_1_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__23212\,
            in1 => \N__16643\,
            in2 => \N__14444\,
            in3 => \N__16250\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36032\,
            ce => 'H',
            sr => \N__36772\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_1_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__23361\,
            in1 => \N__23051\,
            in2 => \_gnd_net_\,
            in3 => \N__30044\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI9MUS_0_1_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__30045\,
            in1 => \_gnd_net_\,
            in2 => \N__23084\,
            in3 => \N__23362\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_10_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20071\,
            in1 => \N__16697\,
            in2 => \N__23231\,
            in3 => \N__16340\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36032\,
            ce => 'H',
            sr => \N__36772\
        );

    \ppm_encoder_1.init_pulses_11_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23211\,
            in1 => \N__20072\,
            in2 => \N__16316\,
            in3 => \N__16688\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36032\,
            ce => 'H',
            sr => \N__36772\
        );

    \ppm_encoder_1.init_pulses_12_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20073\,
            in1 => \N__16679\,
            in2 => \N__23232\,
            in3 => \N__16622\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36032\,
            ce => 'H',
            sr => \N__36772\
        );

    \ppm_encoder_1.init_pulses_RNI5ATG1_15_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__23075\,
            in2 => \N__30101\,
            in3 => \N__30153\,
            lcout => \ppm_encoder_1.init_pulses_RNI5ATG1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIUHRP_15_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__30154\,
            in1 => \N__23063\,
            in2 => \_gnd_net_\,
            in3 => \N__30092\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_15_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20101\,
            in1 => \N__16814\,
            in2 => \N__23234\,
            in3 => \N__16490\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36022\,
            ce => 'H',
            sr => \N__36773\
        );

    \ppm_encoder_1.init_pulses_18_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__16778\,
            in1 => \N__20084\,
            in2 => \N__16457\,
            in3 => \N__23227\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36022\,
            ce => 'H',
            sr => \N__36773\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_2_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23062\,
            in2 => \_gnd_net_\,
            in3 => \N__30091\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1NZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_13_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20100\,
            in1 => \N__16841\,
            in2 => \N__23233\,
            in3 => \N__16574\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36022\,
            ce => 'H',
            sr => \N__36773\
        );

    \ppm_encoder_1.init_pulses_RNISFRP_13_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__24573\,
            in1 => \N__23061\,
            in2 => \_gnd_net_\,
            in3 => \N__30090\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_4_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14513\,
            lcout => \pid_alt.error_p_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36164\,
            ce => \N__20309\,
            sr => \N__21579\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_2_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30869\,
            in2 => \_gnd_net_\,
            in3 => \N__21633\,
            lcout => alt_kp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36158\,
            ce => \N__25756\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_7_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__17279\,
            in1 => \N__15313\,
            in2 => \N__20222\,
            in3 => \N__23957\,
            lcout => \pid_alt.error_i_acummZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36155\,
            ce => 'H',
            sr => \N__15221\
        );

    \Commands_frame_decoder.source_alt_ki_4_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21629\,
            lcout => alt_ki_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31829\,
            in2 => \_gnd_net_\,
            in3 => \N__21626\,
            lcout => alt_ki_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_2_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30868\,
            lcout => alt_ki_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_3_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31220\,
            in2 => \_gnd_net_\,
            in3 => \N__21628\,
            lcout => alt_ki_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_5_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30745\,
            lcout => alt_ki_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_ki_6_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31369\,
            in2 => \_gnd_net_\,
            in3 => \N__21631\,
            lcout => alt_ki_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36152\,
            ce => \N__28045\,
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNILR6F2_8_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14543\,
            in1 => \N__17226\,
            in2 => \N__20191\,
            in3 => \N__17244\,
            lcout => \pid_alt.error_p_reg_esr_RNILR6F2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_8_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14555\,
            lcout => \pid_alt.error_i_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36148\,
            ce => \N__20303\,
            sr => \N__21573\
        );

    \pid_alt.error_p_reg_esr_RNICFJ71_8_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__17245\,
            in1 => \_gnd_net_\,
            in2 => \N__17231\,
            in3 => \N__14542\,
            lcout => \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8\,
            ltout => \pid_alt.error_p_reg_esr_RNICFJ71Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIR17F2_9_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14818\,
            in1 => \N__18047\,
            in2 => \N__14528\,
            in3 => \N__18063\,
            lcout => \pid_alt.error_p_reg_esr_RNIR17F2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_9_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14525\,
            lcout => \pid_alt.error_i_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36148\,
            ce => \N__20303\,
            sr => \N__21573\
        );

    \pid_alt.error_p_reg_esr_RNIFIJ71_9_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__14819\,
            in1 => \N__18048\,
            in2 => \_gnd_net_\,
            in3 => \N__18064\,
            lcout => \pid_alt.error_p_reg_esr_RNIFIJ71Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15116\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pid_alt.error_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_RNI1N2F_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16997\,
            in3 => \N__14780\,
            lcout => \pid_alt.error_1\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_0\,
            carryout => \pid_alt.error_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_1_c_RNI3Q3F_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17141\,
            in3 => \N__14753\,
            lcout => \pid_alt.error_2\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_1\,
            carryout => \pid_alt.error_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_2_c_RNI5T4F_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__14726\,
            lcout => \pid_alt.error_3\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_2\,
            carryout => \pid_alt.error_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_3_c_RNIKE1T_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23495\,
            in2 => \N__17051\,
            in3 => \N__14696\,
            lcout => \pid_alt.error_4\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_3\,
            carryout => \pid_alt.error_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_4_c_RNINI2T_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23480\,
            in2 => \N__16892\,
            in3 => \N__14669\,
            lcout => \pid_alt.error_5\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_4\,
            carryout => \pid_alt.error_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_5_c_RNIQM3T_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23465\,
            in2 => \N__16925\,
            in3 => \N__14639\,
            lcout => \pid_alt.error_6\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_5\,
            carryout => \pid_alt.error_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_6_c_RNITQ4T_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16910\,
            in2 => \N__17036\,
            in3 => \N__14609\,
            lcout => \pid_alt.error_7\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_6\,
            carryout => \pid_alt.error_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_7_c_RNI9LEM_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17021\,
            in2 => \N__23456\,
            in3 => \N__14999\,
            lcout => \pid_alt.error_8\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pid_alt.error_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_8_c_RNICPFM_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17015\,
            in2 => \N__23591\,
            in3 => \N__14972\,
            lcout => \pid_alt.error_9\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_8\,
            carryout => \pid_alt.error_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_9_c_RNIMMUJ_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17009\,
            in2 => \N__23579\,
            in3 => \N__14945\,
            lcout => \pid_alt.error_10\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_9\,
            carryout => \pid_alt.error_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_10_c_RNI0SDO_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17003\,
            in2 => \N__23567\,
            in3 => \N__14918\,
            lcout => \pid_alt.error_11\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_10\,
            carryout => \pid_alt.error_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_11_c_RNI5JAH_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17171\,
            in2 => \_gnd_net_\,
            in3 => \N__14894\,
            lcout => \pid_alt.error_12\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_11\,
            carryout => \pid_alt.error_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_12_c_RNI7MBH_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17159\,
            in2 => \_gnd_net_\,
            in3 => \N__14870\,
            lcout => \pid_alt.error_13\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_12\,
            carryout => \pid_alt.error_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_13_c_RNI9PCH_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17147\,
            in2 => \_gnd_net_\,
            in3 => \N__14846\,
            lcout => \pid_alt.error_14\,
            ltout => OPEN,
            carryin => \pid_alt.error_cry_13\,
            carryout => \pid_alt.error_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_14_c_RNIBSDH_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16937\,
            in2 => \_gnd_net_\,
            in3 => \N__14843\,
            lcout => \pid_alt.error_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNILF5T_6_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__17296\,
            in1 => \_gnd_net_\,
            in2 => \N__17275\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.m35_e_2\,
            ltout => \pid_alt.m35_e_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNID8TA3_5_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__17325\,
            in1 => \N__15049\,
            in2 => \N__15080\,
            in3 => \N__15268\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNID8TA3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI4CCV_10_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17188\,
            in1 => \N__17853\,
            in2 => \N__17938\,
            in3 => \N__18010\,
            lcout => \pid_alt.m35_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNICP62_10_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17931\,
            in2 => \_gnd_net_\,
            in3 => \N__17766\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI56PT1_1_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17068\,
            in1 => \N__18203\,
            in2 => \N__15038\,
            in3 => \N__15032\,
            lcout => \pid_alt.m21_e_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNID75T_2_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__17602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17533\,
            lcout => OPEN,
            ltout => \pid_alt.m21_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI9BT82_7_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__17268\,
            in1 => \N__17324\,
            in2 => \N__15035\,
            in3 => \N__17436\,
            lcout => \pid_alt.m21_e_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIPNRC1_11_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18009\,
            in1 => \N__17187\,
            in2 => \N__17857\,
            in3 => \N__17295\,
            lcout => \pid_alt.m21_e_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23769\,
            in2 => \N__23817\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_0_c_RNIUVGK_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20738\,
            in2 => \N__23549\,
            in3 => \N__15026\,
            lcout => \scaler_2.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_0\,
            carryout => \scaler_2.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_1_c_RNI14IK_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20729\,
            in2 => \N__23537\,
            in3 => \N__15140\,
            lcout => \scaler_2.un3_source_data_0_cry_1_c_RNI14IK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_1\,
            carryout => \scaler_2.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_2_c_RNI48JK_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20720\,
            in2 => \N__23525\,
            in3 => \N__15137\,
            lcout => \scaler_2.un3_source_data_0_cry_2_c_RNI48JK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_2\,
            carryout => \scaler_2.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_3_c_RNI7CKK_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23513\,
            in2 => \N__20711\,
            in3 => \N__15134\,
            lcout => \scaler_2.un3_source_data_0_cry_3_c_RNI7CKK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_3\,
            carryout => \scaler_2.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_4_c_RNIAGLK_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23669\,
            in2 => \N__20699\,
            in3 => \N__15131\,
            lcout => \scaler_2.un3_source_data_0_cry_4_c_RNIAGLK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_4\,
            carryout => \scaler_2.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_5_c_RNIDKMK_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23660\,
            in2 => \N__20687\,
            in3 => \N__15128\,
            lcout => \scaler_2.un3_source_data_0_cry_5_c_RNIDKMK\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_5\,
            carryout => \scaler_2.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_6_c_RNIIUTM_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21062\,
            in2 => \_gnd_net_\,
            in3 => \N__15125\,
            lcout => \scaler_2.un3_source_data_0_cry_6_c_RNIIUTM\,
            ltout => OPEN,
            carryin => \scaler_2.un3_source_data_0_cry_6\,
            carryout => \scaler_2.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_7_c_RNIJ0VM_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21080\,
            in2 => \N__28690\,
            in3 => \N__15122\,
            lcout => \scaler_2.un3_source_data_0_cry_7_c_RNIJ0VM\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \scaler_2.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_cry_8_c_RNIQL42_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15119\,
            lcout => \scaler_2.un3_source_data_0_cry_8_c_RNIQL42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_cry_0_c_inv_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__15109\,
            in1 => \N__28659\,
            in2 => \_gnd_net_\,
            in3 => \N__15345\,
            lcout => \pid_alt.drone_altitude_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_0_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26125\,
            lcout => drone_altitude_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36126\,
            ce => \N__25703\,
            sr => \N__36717\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNI24S01_12_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011101110"
        )
    port map (
            in0 => \N__18320\,
            in1 => \N__15281\,
            in2 => \N__17780\,
            in3 => \N__17686\,
            lcout => \pid_alt.error_i_acumm_prereg_esr_RNI24S01Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_RNISOGT_14_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18413\,
            in1 => \N__18085\,
            in2 => \N__18559\,
            in3 => \N__18109\,
            lcout => \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14\,
            ltout => \pid_alt.error_i_acumm_prereg_RNISOGTZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_esr_13_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18318\,
            in2 => \N__15275\,
            in3 => \N__17687\,
            lcout => \pid_alt.error_i_acummZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36121\,
            ce => \N__15166\,
            sr => \N__15208\
        );

    \pid_alt.error_i_acumm_prereg_RNINGKC_14_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18552\,
            in1 => \N__18084\,
            in2 => \_gnd_net_\,
            in3 => \N__18108\,
            lcout => OPEN,
            ltout => \pid_alt.error_i_acumm_prereg_RNINGKCZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIBMOV_13_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__18319\,
            in1 => \N__17685\,
            in2 => \N__15272\,
            in3 => \N__18412\,
            lcout => \pid_alt.N_9_0\,
            ltout => \pid_alt.N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75_21_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__18317\,
            in1 => \N__15245\,
            in2 => \N__15236\,
            in3 => \N__15233\,
            lcout => OPEN,
            ltout => \pid_alt.error_i_acumm_prereg_esr_RNIGMJ75Z0Z_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNI2P1V5_1_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23912\,
            in2 => \N__15224\,
            in3 => \N__35080\,
            lcout => \pid_alt.un1_reset_1_0_i\,
            ltout => \pid_alt.un1_reset_1_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNINE9D6_1_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__23913\,
            in1 => \_gnd_net_\,
            in2 => \N__15173\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.N_60_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CRY_0_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15535\,
            in2 => \N__15542\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_0_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18264\,
            in2 => \N__18248\,
            in3 => \N__15512\,
            lcout => \pid_alt.pid_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_un1_pid_prereg_0_cry_0_c_THRU_CO\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_0\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.un1_pid_prereg_0_cry_0_THRU_LUT4_0_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21130\,
            in2 => \_gnd_net_\,
            in3 => \N__15509\,
            lcout => \pid_alt.un1_pid_prereg_0_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_0\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_2_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15506\,
            in2 => \N__15500\,
            in3 => \N__15491\,
            lcout => \pid_alt.pid_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_1\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_2\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.pid_prereg_esr_3_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15484\,
            in2 => \N__15473\,
            in3 => \N__15461\,
            lcout => \pid_alt.pid_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_2\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_3\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.pid_prereg_esr_4_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15458\,
            in2 => \N__15449\,
            in3 => \N__15434\,
            lcout => \pid_alt.pid_preregZ0Z_4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_3\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_4\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.pid_prereg_esr_5_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15431\,
            in2 => \N__15409\,
            in3 => \N__15386\,
            lcout => \pid_alt.pid_preregZ0Z_5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_4\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_5\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.pid_prereg_esr_6_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15383\,
            in2 => \N__15374\,
            in3 => \N__15365\,
            lcout => \pid_alt.pid_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_5\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_6\,
            clk => \N__36116\,
            ce => \N__18297\,
            sr => \N__36726\
        );

    \pid_alt.pid_prereg_esr_7_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20339\,
            in2 => \N__20360\,
            in3 => \N__15800\,
            lcout => \pid_alt.pid_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_7\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_8_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15797\,
            in2 => \N__20192\,
            in3 => \N__15788\,
            lcout => \pid_alt.pid_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_7\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_8\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_9_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15785\,
            in2 => \N__15776\,
            in3 => \N__15758\,
            lcout => \pid_alt.pid_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_8\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_9\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_10_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15754\,
            in2 => \N__15725\,
            in3 => \N__15710\,
            lcout => \pid_alt.pid_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_9\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_10\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_11_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15707\,
            in2 => \N__15686\,
            in3 => \N__15668\,
            lcout => \pid_alt.pid_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_10\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_11\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_12_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15665\,
            in2 => \N__15650\,
            in3 => \N__15635\,
            lcout => \pid_alt.pid_preregZ0Z_12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_11\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_12\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_13_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15632\,
            in2 => \N__15614\,
            in3 => \N__15584\,
            lcout => \pid_alt.pid_preregZ0Z_13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_12\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_13\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_14_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15581\,
            in2 => \N__15566\,
            in3 => \N__15545\,
            lcout => \pid_alt.pid_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_13\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_14\,
            clk => \N__36110\,
            ce => \N__18298\,
            sr => \N__36729\
        );

    \pid_alt.pid_prereg_esr_15_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15974\,
            in2 => \N__15962\,
            in3 => \N__15944\,
            lcout => \pid_alt.pid_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_15\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_16_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15941\,
            in2 => \N__15926\,
            in3 => \N__15911\,
            lcout => \pid_alt.pid_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_15\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_16\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_17_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15908\,
            in2 => \N__18461\,
            in3 => \N__15896\,
            lcout => \pid_alt.pid_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_16\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_17\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_18_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15893\,
            in2 => \N__15878\,
            in3 => \N__15866\,
            lcout => \pid_alt.pid_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_17\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_18\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_19_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20552\,
            in2 => \N__15863\,
            in3 => \N__15851\,
            lcout => \pid_alt.pid_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_18\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_19\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_20_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15848\,
            in2 => \N__15836\,
            in3 => \N__15818\,
            lcout => \pid_alt.pid_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_19\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_20\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_21_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15815\,
            in2 => \N__20756\,
            in3 => \N__15806\,
            lcout => \pid_alt.pid_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \pid_alt.un1_pid_prereg_0_cry_20\,
            carryout => \pid_alt.un1_pid_prereg_0_cry_21\,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_22_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__20882\,
            in1 => \N__20810\,
            in2 => \_gnd_net_\,
            in3 => \N__15803\,
            lcout => \pid_alt.pid_preregZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36104\,
            ce => \N__18299\,
            sr => \N__36735\
        );

    \pid_alt.pid_prereg_esr_RNI8OUM_14_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16064\,
            in1 => \N__16055\,
            in2 => \N__16049\,
            in3 => \N__16040\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIQORD1_15_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16034\,
            in1 => \N__16028\,
            in2 => \N__16022\,
            in3 => \N__16004\,
            lcout => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15\,
            ltout => \pid_alt.pid_prereg_esr_RNIQORD1Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_RNO_0_4_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__19398\,
            in1 => \N__19488\,
            in2 => \N__16019\,
            in3 => \N__19165\,
            lcout => \pid_alt.source_pid_9_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIBIEB_17_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16016\,
            in2 => \_gnd_net_\,
            in3 => \N__16010\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_13_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19330\,
            in2 => \N__19414\,
            in3 => \N__19005\,
            lcout => throttle_command_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36097\,
            ce => \N__19284\,
            sr => \N__19249\
        );

    \pid_alt.source_pid_1_esr_12_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__19197\,
            in1 => \N__19402\,
            in2 => \N__19010\,
            in3 => \N__19335\,
            lcout => throttle_command_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36097\,
            ce => \N__19284\,
            sr => \N__19249\
        );

    \pid_alt.source_pid_1_esr_1_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__19331\,
            in1 => \N__19448\,
            in2 => \N__19425\,
            in3 => \N__21104\,
            lcout => throttle_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36090\,
            ce => \N__19285\,
            sr => \N__19256\
        );

    \pid_alt.source_pid_1_esr_4_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__18952\,
            in2 => \N__15998\,
            in3 => \N__19490\,
            lcout => throttle_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36090\,
            ce => \N__19285\,
            sr => \N__19256\
        );

    \pid_alt.source_pid_1_esr_5_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__19419\,
            in2 => \N__19223\,
            in3 => \N__19334\,
            lcout => throttle_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36090\,
            ce => \N__19285\,
            sr => \N__19256\
        );

    \pid_alt.source_pid_1_esr_0_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__19447\,
            in1 => \N__19415\,
            in2 => \N__18680\,
            in3 => \N__19333\,
            lcout => throttle_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36090\,
            ce => \N__19285\,
            sr => \N__19256\
        );

    \ppm_encoder_1.throttle_RNIG4JI2_11_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16074\,
            in1 => \N__21475\,
            in2 => \N__22358\,
            in3 => \N__22263\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIALRT5_11_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22628\,
            in2 => \N__16148\,
            in3 => \N__16145\,
            lcout => \ppm_encoder_1.elevator_RNIALRT5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI03DH2_11_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16122\,
            in1 => \N__16134\,
            in2 => \N__22123\,
            in3 => \N__22001\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_11_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29490\,
            in1 => \N__16075\,
            in2 => \_gnd_net_\,
            in3 => \N__16123\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_11_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29268\,
            in2 => \N__16139\,
            in3 => \N__16135\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_11_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__16136\,
            in1 => \N__24970\,
            in2 => \N__21260\,
            in3 => \N__19070\,
            lcout => \ppm_encoder_1.aileronZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36082\,
            ce => 'H',
            sr => \N__36751\
        );

    \ppm_encoder_1.elevator_11_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__16124\,
            in1 => \N__29738\,
            in2 => \N__24997\,
            in3 => \N__24440\,
            lcout => \ppm_encoder_1.elevatorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36082\,
            ce => 'H',
            sr => \N__36751\
        );

    \ppm_encoder_1.throttle_11_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__16112\,
            in1 => \N__16076\,
            in2 => \N__16085\,
            in3 => \N__24971\,
            lcout => \ppm_encoder_1.throttleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36082\,
            ce => 'H',
            sr => \N__36751\
        );

    \ppm_encoder_1.throttle_RNIQ3KK2_7_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16158\,
            in1 => \N__22314\,
            in2 => \N__21445\,
            in3 => \N__22261\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIJII96_7_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19712\,
            in2 => \N__16232\,
            in3 => \N__16229\,
            lcout => \ppm_encoder_1.throttle_RNIJII96Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIAIVN2_7_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16206\,
            in1 => \N__16218\,
            in2 => \N__22106\,
            in3 => \N__21999\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_7_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29462\,
            in1 => \N__16159\,
            in2 => \_gnd_net_\,
            in3 => \N__16207\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_7_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29262\,
            in1 => \_gnd_net_\,
            in2 => \N__16223\,
            in3 => \N__16219\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_7_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__16220\,
            in1 => \N__18908\,
            in2 => \N__24998\,
            in3 => \N__20978\,
            lcout => \ppm_encoder_1.aileronZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36073\,
            ce => 'H',
            sr => \N__36754\
        );

    \ppm_encoder_1.elevator_7_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__16208\,
            in1 => \N__24080\,
            in2 => \N__28988\,
            in3 => \N__24980\,
            lcout => \ppm_encoder_1.elevatorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36073\,
            ce => 'H',
            sr => \N__36754\
        );

    \ppm_encoder_1.throttle_7_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__16196\,
            in1 => \N__16183\,
            in2 => \N__24999\,
            in3 => \N__16160\,
            lcout => \ppm_encoder_1.throttleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36073\,
            ce => 'H',
            sr => \N__36754\
        );

    \ppm_encoder_1.elevator_RNI47DH2_13_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__24335\,
            in2 => \N__29534\,
            in3 => \N__22082\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIKVRT5_13_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16607\,
            in2 => \N__16304\,
            in3 => \N__16292\,
            lcout => \ppm_encoder_1.elevator_RNIKVRT5Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI8GVN2_6_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__21996\,
            in1 => \N__29302\,
            in2 => \N__29123\,
            in3 => \N__22078\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIO1KK2_6_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__29325\,
            in1 => \N__24607\,
            in2 => \N__22342\,
            in3 => \N__22224\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIEDI96_6_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19862\,
            in2 => \N__16301\,
            in3 => \N__16298\,
            lcout => \ppm_encoder_1.throttle_RNIEDI96Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIK8JI2_13_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__23693\,
            in1 => \N__24560\,
            in2 => \N__22341\,
            in3 => \N__22223\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIOIR62_5_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__16285\,
            in1 => \N__16273\,
            in2 => \N__22105\,
            in3 => \N__21997\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIVO123_0_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16256\,
            in2 => \N__19837\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_1_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19126\,
            in2 => \N__19100\,
            in3 => \N__16238\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_2_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19562\,
            in2 => \N__19502\,
            in3 => \N__16235\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_3_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19652\,
            in2 => \N__19640\,
            in3 => \N__16439\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_4_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19526\,
            in2 => \N__20168\,
            in3 => \N__16436\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_5_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16433\,
            in2 => \N__16412\,
            in3 => \N__16403\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_6_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19861\,
            in2 => \N__16400\,
            in3 => \N__16391\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_7_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19708\,
            in2 => \N__16388\,
            in3 => \N__16376\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_8_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22159\,
            in2 => \N__22145\,
            in3 => \N__16373\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_8\,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_9_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19576\,
            in2 => \N__16370\,
            in3 => \N__16352\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_10_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19609\,
            in2 => \N__16349\,
            in3 => \N__16331\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_11_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22627\,
            in2 => \N__16328\,
            in3 => \N__16625\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_12_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21781\,
            in2 => \N__21767\,
            in3 => \N__16610\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_13_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16603\,
            in2 => \N__16586\,
            in3 => \N__16562\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_14_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16559\,
            in2 => \N__16553\,
            in3 => \N__16520\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_15_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16517\,
            in2 => \N__16505\,
            in3 => \N__16478\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_16_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16664\,
            in2 => \_gnd_net_\,
            in3 => \N__16475\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_16\,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_17_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16445\,
            in2 => \_gnd_net_\,
            in3 => \N__16463\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_0_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_0_18_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16670\,
            in2 => \_gnd_net_\,
            in3 => \N__16460\,
            lcout => \ppm_encoder_1.un1_init_pulses_10_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_0_17_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__30342\,
            in1 => \_gnd_net_\,
            in2 => \N__30097\,
            in3 => \N__22985\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_2_18_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__19922\,
            in1 => \N__30304\,
            in2 => \N__23045\,
            in3 => \N__30072\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_0_16_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__30394\,
            in1 => \_gnd_net_\,
            in2 => \N__30096\,
            in3 => \N__22983\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI0KRP_17_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__22984\,
            in1 => \N__30065\,
            in2 => \_gnd_net_\,
            in3 => \N__30343\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIAVNR2_0_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23292\,
            in1 => \N__24374\,
            in2 => \N__30098\,
            in3 => \N__19921\,
            lcout => \ppm_encoder_1.init_pulses_RNIAVNR2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC9HQ4_0_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16658\,
            in2 => \N__22655\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_28_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_1_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16652\,
            in3 => \N__16637\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_0\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_2_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19631\,
            in2 => \N__19973\,
            in3 => \N__16634\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_1\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_3_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19742\,
            in2 => \_gnd_net_\,
            in3 => \N__16631\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_2\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_4_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20144\,
            in2 => \_gnd_net_\,
            in3 => \N__16628\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_3\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_5_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16760\,
            in2 => \_gnd_net_\,
            in3 => \N__16748\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_4\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_6_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16745\,
            in2 => \N__19892\,
            in3 => \N__16739\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_5\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_7_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19718\,
            in2 => \_gnd_net_\,
            in3 => \N__16736\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_6\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_8_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16733\,
            in2 => \_gnd_net_\,
            in3 => \N__16724\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_8\,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_9_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16721\,
            in2 => \_gnd_net_\,
            in3 => \N__16700\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_8\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_10_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19541\,
            in2 => \_gnd_net_\,
            in3 => \N__16691\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_9\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_11_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23306\,
            in2 => \_gnd_net_\,
            in3 => \N__16682\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_10\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_12_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19979\,
            in2 => \_gnd_net_\,
            in3 => \N__16673\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_11\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_13_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16856\,
            in2 => \N__16850\,
            in3 => \N__16835\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_12\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_14_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19991\,
            in3 => \N__16826\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_13\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_15_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16823\,
            in2 => \_gnd_net_\,
            in3 => \N__16808\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_14\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_16_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22871\,
            in2 => \_gnd_net_\,
            in3 => \N__16805\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_16\,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_17_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16802\,
            in2 => \_gnd_net_\,
            in3 => \N__16784\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_init_pulses_3_cry_16\,
            carryout => \ppm_encoder_1.un1_init_pulses_3_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNO_1_18_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__30294\,
            in1 => \N__23088\,
            in2 => \N__30100\,
            in3 => \N__16781\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__30076\,
            in1 => \N__29388\,
            in2 => \N__29279\,
            in3 => \N__36912\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_3_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31222\,
            in2 => \_gnd_net_\,
            in3 => \N__21637\,
            lcout => alt_kp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36162\,
            ce => \N__25757\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_5_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31373\,
            lcout => alt_kp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36162\,
            ce => \N__25757\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_0_e_0_4_LC_3_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30749\,
            in2 => \_gnd_net_\,
            in3 => \N__21635\,
            lcout => alt_kp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36162\,
            ce => \N__25757\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_1_LC_3_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31841\,
            lcout => alt_kp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36162\,
            ce => \N__25757\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_0_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31499\,
            in2 => \_gnd_net_\,
            in3 => \N__21632\,
            lcout => alt_kp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36159\,
            ce => \N__25754\,
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_15_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26183\,
            lcout => drone_altitude_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36149\,
            ce => \N__25652\,
            sr => \N__36693\
        );

    \Commands_frame_decoder.source_CH1data_2_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__30846\,
            in1 => \N__25843\,
            in2 => \N__16874\,
            in3 => \N__16924\,
            lcout => alt_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36145\,
            ce => 'H',
            sr => \N__36695\
        );

    \Commands_frame_decoder.source_CH1data_3_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__25844\,
            in1 => \N__16866\,
            in2 => \N__31221\,
            in3 => \N__16906\,
            lcout => alt_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36145\,
            ce => 'H',
            sr => \N__36695\
        );

    \Commands_frame_decoder.source_CH1data_1_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__31840\,
            in1 => \N__25842\,
            in2 => \N__16873\,
            in3 => \N__16891\,
            lcout => alt_command_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36145\,
            ce => 'H',
            sr => \N__36695\
        );

    \Commands_frame_decoder.source_CH1data8lto3_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__31210\,
            in1 => \N__30845\,
            in2 => \_gnd_net_\,
            in3 => \N__31839\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.source_CH1data8lt7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data8lto7_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__31360\,
            in1 => \N__31654\,
            in2 => \N__16877\,
            in3 => \N__28070\,
            lcout => \Commands_frame_decoder.source_CH1data8\,
            ltout => \Commands_frame_decoder.source_CH1data8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__25841\,
            in1 => \N__31498\,
            in2 => \N__17054\,
            in3 => \N__17050\,
            lcout => alt_command_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36145\,
            ce => 'H',
            sr => \N__36695\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIKLDC_7_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17027\,
            lcout => drone_altitude_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_7_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26179\,
            lcout => \dron_frame_decoder_1.drone_altitude_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36141\,
            ce => \N__25709\,
            sr => \N__36701\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNILMDC_8_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20657\,
            lcout => drone_altitude_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIMNDC_9_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20669\,
            lcout => drone_altitude_i_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIUHR9_10_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20663\,
            lcout => drone_altitude_i_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIVIR9_11_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20675\,
            lcout => drone_altitude_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_1_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16988\,
            lcout => \pid_alt.error_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_1_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26090\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => drone_altitude_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36141\,
            ce => \N__25709\,
            sr => \N__36701\
        );

    \pid_alt.error_axb_12_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17165\,
            lcout => \pid_alt.error_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_12_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25963\,
            lcout => drone_altitude_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36136\,
            ce => \N__25648\,
            sr => \N__36705\
        );

    \pid_alt.error_axb_13_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17153\,
            lcout => \pid_alt.error_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_13_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26261\,
            lcout => drone_altitude_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36136\,
            ce => \N__25648\,
            sr => \N__36705\
        );

    \pid_alt.error_axb_14_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20651\,
            lcout => \pid_alt.error_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_2_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20645\,
            lcout => \pid_alt.error_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_axb_3_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20639\,
            lcout => \pid_alt.error_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_un1_error_i_acumm_prereg_cry_0_c_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18271\,
            in2 => \N__18240\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_1_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17126\,
            in2 => \N__17105\,
            in3 => \N__17057\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_0\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17660\,
            in2 => \N__17636\,
            in3 => \N__17591\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_2\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_1\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_3_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17588\,
            in2 => \N__17567\,
            in3 => \N__17522\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_3\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_2\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_4_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17519\,
            in2 => \N__17498\,
            in3 => \N__17420\,
            lcout => \pid_alt.error_i_acumm7lto4\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_3\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_5_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17417\,
            in2 => \N__17378\,
            in3 => \N__17306\,
            lcout => \pid_alt.error_i_acumm7lto5\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_4\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_6_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20398\,
            in2 => \N__20435\,
            in3 => \N__17282\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_6\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_5\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_7_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20223\,
            in2 => \N__20249\,
            in3 => \N__17255\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_7\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_6\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_7\,
            clk => \N__36132\,
            ce => \N__18294\,
            sr => \N__36707\
        );

    \pid_alt.error_i_acumm_prereg_esr_8_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17252\,
            in2 => \N__17230\,
            in3 => \N__17174\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.error_i_acumm_prereg_esr_9_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18071\,
            in2 => \N__18049\,
            in3 => \N__17996\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_9\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_8\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.error_i_acumm_prereg_esr_10_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17993\,
            in2 => \N__17972\,
            in3 => \N__17918\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_10\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_9\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.error_i_acumm_prereg_esr_11_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17915\,
            in2 => \N__17894\,
            in3 => \N__17837\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_11\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_10\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.error_i_acumm_prereg_esr_12_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17834\,
            in2 => \N__17813\,
            in3 => \N__17750\,
            lcout => \pid_alt.error_i_acumm7lto12\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_11\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.error_i_acumm_prereg_esr_13_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17740\,
            in2 => \N__17720\,
            in3 => \N__17672\,
            lcout => \pid_alt.error_i_acumm7lto13\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_12\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            clk => \N__36127\,
            ce => \N__18295\,
            sr => \N__36711\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_LUT4_0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18157\,
            in2 => \_gnd_net_\,
            in3 => \N__17669\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_13\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_LUT4_0_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18388\,
            in3 => \N__17666\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_14\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_LUT4_0_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18509\,
            in2 => \_gnd_net_\,
            in3 => \N__17663\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_LUT4_0_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18877\,
            in2 => \_gnd_net_\,
            in3 => \N__18335\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_16\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_LUT4_0_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20629\,
            in2 => \_gnd_net_\,
            in3 => \N__18332\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_17\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_LUT4_0_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18604\,
            in2 => \_gnd_net_\,
            in3 => \N__18329\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_18\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_LUT4_0_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20873\,
            in2 => \_gnd_net_\,
            in3 => \N__18326\,
            lcout => \pid_alt.un1_error_i_acumm_prereg_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \pid_alt.un1_error_i_acumm_prereg_cry_19\,
            carryout => \pid_alt.un1_error_i_acumm_prereg_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_esr_21_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18323\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36122\,
            ce => \N__18296\,
            sr => \N__36713\
        );

    \pid_alt.error_i_acumm_prereg_0_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__18275\,
            in1 => \N__34163\,
            in2 => \N__18247\,
            in3 => \N__18195\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36117\,
            ce => 'H',
            sr => \N__36718\
        );

    \pid_alt.error_i_acumm_prereg_20_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__34162\,
            in1 => \N__18176\,
            in2 => \N__20881\,
            in3 => \N__18427\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36117\,
            ce => 'H',
            sr => \N__36718\
        );

    \pid_alt.error_i_acumm_prereg_14_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__18167\,
            in1 => \N__34164\,
            in2 => \N__18158\,
            in3 => \N__18110\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36117\,
            ce => 'H',
            sr => \N__36718\
        );

    \pid_alt.error_i_acumm_prereg_16_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__34161\,
            in1 => \N__18095\,
            in2 => \N__18089\,
            in3 => \N__18508\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36117\,
            ce => 'H',
            sr => \N__36718\
        );

    \pid_alt.error_i_acumm_prereg_19_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010010111000"
        )
    port map (
            in0 => \N__18611\,
            in1 => \N__34165\,
            in2 => \N__18560\,
            in3 => \N__18566\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36117\,
            ce => 'H',
            sr => \N__36718\
        );

    \pid_alt.error_p_reg_esr_RNIB03K_16_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18507\,
            lcout => \pid_alt.error_p_reg_esr_RNIB03KZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIC2521_1_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__29494\,
            in1 => \N__29275\,
            in2 => \_gnd_net_\,
            in3 => \N__22421\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_14_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29274\,
            in1 => \N__18446\,
            in2 => \_gnd_net_\,
            in3 => \N__19051\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_4_3_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26003\,
            in1 => \N__25962\,
            in2 => \N__26230\,
            in3 => \N__26082\,
            lcout => \dron_frame_decoder_1.N_194_4\,
            ltout => \dron_frame_decoder_1.N_194_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_0_3_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__24028\,
            in1 => \_gnd_net_\,
            in2 => \N__18431\,
            in3 => \_gnd_net_\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_RNI58SG_15_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18817\,
            in1 => \N__18835\,
            in2 => \N__18428\,
            in3 => \N__18343\,
            lcout => \pid_alt.m7_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_acumm_prereg_15_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010101010"
        )
    port map (
            in0 => \N__18344\,
            in1 => \N__18404\,
            in2 => \N__18395\,
            in3 => \N__34160\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36111\,
            ce => 'H',
            sr => \N__36723\
        );

    \pid_alt.error_i_acumm_prereg_17_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__34158\,
            in1 => \N__18890\,
            in2 => \N__18881\,
            in3 => \N__18836\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36111\,
            ce => 'H',
            sr => \N__36723\
        );

    \pid_alt.error_i_acumm_prereg_18_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__18827\,
            in1 => \N__34159\,
            in2 => \N__20633\,
            in3 => \N__18818\,
            lcout => \pid_alt.error_i_acumm_preregZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36111\,
            ce => 'H',
            sr => \N__36723\
        );

    \pid_alt.pid_prereg_esr_RNIC62V1_12_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__18994\,
            in1 => \N__19188\,
            in2 => \N__19413\,
            in3 => \N__19336\,
            lcout => \pid_alt.source_pid_9_0_tz_6\,
            ltout => \pid_alt.source_pid_9_0_tz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_8_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__21909\,
            in1 => \N__18775\,
            in2 => \N__18782\,
            in3 => \N__23886\,
            lcout => throttle_command_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36105\,
            ce => 'H',
            sr => \N__19261\
        );

    \pid_alt.pid_prereg_esr_RNIT3KA1_11_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18753\,
            in1 => \N__18774\,
            in2 => \N__18705\,
            in3 => \N__18729\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI8H141_10_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__18779\,
            in1 => \N__18754\,
            in2 => \N__18736\,
            in3 => \N__18654\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIFQKS1_6_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18636\,
            in2 => \N__18713\,
            in3 => \N__18706\,
            lcout => \pid_alt.pid_prereg_esr_RNIFQKS1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIHBUI1_0_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__19360\,
            in2 => \N__19030\,
            in3 => \N__18676\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI4GSA2_10_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18655\,
            in1 => \N__18637\,
            in2 => \N__18623\,
            in3 => \N__23868\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI845S4_4_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19481\,
            in1 => \N__18938\,
            in2 => \N__18941\,
            in3 => \N__19164\,
            lcout => \pid_alt.source_pid_1_sqmuxa_0_a2_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIP29I1_4_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19000\,
            in1 => \N__23869\,
            in2 => \N__19169\,
            in3 => \N__19480\,
            lcout => OPEN,
            ltout => \pid_alt.source_pid_1_sqmuxa_0_a2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIJ1OF6_4_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19322\,
            in1 => \N__18937\,
            in2 => \N__18926\,
            in3 => \N__18964\,
            lcout => OPEN,
            ltout => \pid_alt.N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNIM9UC7_22_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__19394\,
            in1 => \N__23870\,
            in2 => \N__18923\,
            in3 => \N__35081\,
            lcout => OPEN,
            ltout => \pid_alt.un1_reset_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI9BMSD_13_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__19323\,
            in1 => \N__19001\,
            in2 => \N__18920\,
            in3 => \N__18917\,
            lcout => \pid_alt.un1_reset_0_i\,
            ltout => \pid_alt.un1_reset_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIU0UAE_1_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18911\,
            in3 => \N__23871\,
            lcout => \pid_alt.N_60_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_c_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \ppm_encoder_1.un1_aileron_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_6_THRU_LUT4_0_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20974\,
            in2 => \_gnd_net_\,
            in3 => \N__18896\,
            lcout => \ppm_encoder_1.un1_aileron_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_6\,
            carryout => \ppm_encoder_1.un1_aileron_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_7_THRU_LUT4_0_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21871\,
            in2 => \_gnd_net_\,
            in3 => \N__18893\,
            lcout => \ppm_encoder_1.un1_aileron_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_7\,
            carryout => \ppm_encoder_1.un1_aileron_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_8_THRU_LUT4_0_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20908\,
            in2 => \_gnd_net_\,
            in3 => \N__19076\,
            lcout => \ppm_encoder_1.un1_aileron_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_8\,
            carryout => \ppm_encoder_1.un1_aileron_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_9_THRU_LUT4_0_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24199\,
            in2 => \_gnd_net_\,
            in3 => \N__19073\,
            lcout => \ppm_encoder_1.un1_aileron_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_9\,
            carryout => \ppm_encoder_1.un1_aileron_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_10_THRU_LUT4_0_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21256\,
            in2 => \_gnd_net_\,
            in3 => \N__19064\,
            lcout => \ppm_encoder_1.un1_aileron_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_10\,
            carryout => \ppm_encoder_1.un1_aileron_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_11_THRU_LUT4_0_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21742\,
            in2 => \_gnd_net_\,
            in3 => \N__19061\,
            lcout => \ppm_encoder_1.un1_aileron_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_11\,
            carryout => \ppm_encoder_1.un1_aileron_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_aileron_cry_12_THRU_LUT4_0_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24133\,
            in2 => \N__28602\,
            in3 => \N__19058\,
            lcout => \ppm_encoder_1.un1_aileron_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_aileron_cry_12\,
            carryout => \ppm_encoder_1.un1_aileron_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_14_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21164\,
            in2 => \_gnd_net_\,
            in3 => \N__19055\,
            lcout => \ppm_encoder_1.aileronZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36074\,
            ce => \N__27301\,
            sr => \N__36744\
        );

    \ppm_encoder_1.aileron_esr_4_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23741\,
            lcout => \ppm_encoder_1.aileronZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36074\,
            ce => \N__27301\,
            sr => \N__36744\
        );

    \pid_alt.source_pid_1_esr_3_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__19441\,
            in1 => \N__19031\,
            in2 => \N__19430\,
            in3 => \N__19343\,
            lcout => throttle_command_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36063\,
            ce => \N__19286\,
            sr => \N__19262\
        );

    \pid_alt.pid_prereg_esr_RNIG2382_12_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__19199\,
            in1 => \N__19009\,
            in2 => \_gnd_net_\,
            in3 => \N__18968\,
            lcout => \pid_alt.N_88\,
            ltout => \pid_alt.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_esr_RNI3BD63_4_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110010"
        )
    port map (
            in0 => \N__19154\,
            in1 => \N__19489\,
            in2 => \N__19451\,
            in3 => \_gnd_net_\,
            lcout => \pid_alt.N_90\,
            ltout => \pid_alt.N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_pid_1_esr_2_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__19426\,
            in1 => \N__19364\,
            in2 => \N__19346\,
            in3 => \N__19342\,
            lcout => throttle_command_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36063\,
            ce => \N__19286\,
            sr => \N__19262\
        );

    \pid_alt.pid_prereg_esr_RNIIM0I_5_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19222\,
            in2 => \_gnd_net_\,
            in3 => \N__19198\,
            lcout => \pid_alt.N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25267\,
            in1 => \N__22482\,
            in2 => \N__22406\,
            in3 => \N__30024\,
            lcout => \ppm_encoder_1.init_pulses_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22543\,
            in1 => \N__22527\,
            in2 => \N__30025\,
            in3 => \N__22407\,
            lcout => \ppm_encoder_1.init_pulses_1_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_1_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNIHFK13_0_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__22002\,
            in1 => \N__22433\,
            in2 => \N__19133\,
            in3 => \N__29928\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIALN65_1_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001111"
        )
    port map (
            in0 => \N__25058\,
            in1 => \N__19130\,
            in2 => \N__19103\,
            in3 => \N__22222\,
            lcout => \ppm_encoder_1.throttle_RNIALN65Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIMGR62_4_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__19774\,
            in1 => \N__26677\,
            in2 => \N__22016\,
            in3 => \N__22095\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_esr_RNIV9IN5_4_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__20164\,
            in1 => \_gnd_net_\,
            in2 => \N__19529\,
            in3 => \N__19514\,
            lcout => \ppm_encoder_1.aileron_esr_RNIV9IN5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI6LFQ_0_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__22450\,
            in1 => \N__22576\,
            in2 => \N__22529\,
            in3 => \N__22542\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI5QE01_0_0_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__29927\,
            in1 => \_gnd_net_\,
            in2 => \N__19520\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.init_pulses_3_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_3_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_RNITVNJ2_4_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__21844\,
            in1 => \N__22202\,
            in2 => \N__19517\,
            in3 => \N__26641\,
            lcout => \ppm_encoder_1.un2_throttle_iv_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_RNI7RM01_0_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22481\,
            in1 => \N__25266\,
            in2 => \N__22405\,
            in3 => \N__29879\,
            lcout => \ppm_encoder_1.init_pulses_0_sqmuxa_0\,
            ltout => \ppm_encoder_1.init_pulses_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIR7352_2_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__20533\,
            in1 => \N__22771\,
            in2 => \N__19508\,
            in3 => \N__19917\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI5V123_2_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19505\,
            in3 => \N__19552\,
            lcout => \ppm_encoder_1.throttle_RNI5V123Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_3_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29880\,
            in1 => \N__25185\,
            in2 => \_gnd_net_\,
            in3 => \N__22948\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIT9352_3_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010100101"
        )
    port map (
            in0 => \N__25186\,
            in1 => \N__24769\,
            in2 => \N__19935\,
            in3 => \N__22249\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un1_init_pulses_0_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNI82223_3_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19493\,
            in3 => \N__19651\,
            lcout => \ppm_encoder_1.throttle_RNI82223Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_12_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22950\,
            in1 => \N__27838\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIGTUS_8_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29881\,
            in1 => \N__24258\,
            in2 => \_gnd_net_\,
            in3 => \N__22949\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_1_1_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23253\,
            in2 => \_gnd_net_\,
            in3 => \N__29885\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI8J2H_2_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22575\,
            in2 => \_gnd_net_\,
            in3 => \N__25215\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_d_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI7O1N_0_2_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19619\,
            in3 => \N__29883\,
            lcout => \ppm_encoder_1.un1_init_pulses_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_10_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29888\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__22947\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIHUUS_9_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22945\,
            in1 => \N__19598\,
            in2 => \_gnd_net_\,
            in3 => \N__29886\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIANUS_2_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29884\,
            in1 => \N__20529\,
            in2 => \_gnd_net_\,
            in3 => \N__22944\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIPCRP_0_10_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__22946\,
            in1 => \_gnd_net_\,
            in2 => \N__25490\,
            in3 => \N__29887\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_4_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29253\,
            in1 => \N__21824\,
            in2 => \_gnd_net_\,
            in3 => \N__19775\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_3_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20124\,
            in1 => \N__19757\,
            in2 => \N__23228\,
            in3 => \N__19751\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36033\,
            ce => 'H',
            sr => \N__36763\
        );

    \ppm_encoder_1.init_pulses_RNIBOUS_0_3_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__25184\,
            in1 => \N__22978\,
            in2 => \_gnd_net_\,
            in3 => \N__29912\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_7_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20125\,
            in1 => \N__19736\,
            in2 => \N__23229\,
            in3 => \N__19730\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36033\,
            ce => 'H',
            sr => \N__36763\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_0_7_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__19693\,
            in1 => \N__22982\,
            in2 => \_gnd_net_\,
            in3 => \N__29914\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIFSUS_7_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__29913\,
            in1 => \_gnd_net_\,
            in2 => \N__23044\,
            in3 => \N__19692\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_7_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__19694\,
            in1 => \N__27941\,
            in2 => \N__30579\,
            in3 => \N__21446\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_8_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__23201\,
            in1 => \N__19682\,
            in2 => \N__19673\,
            in3 => \N__20126\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36033\,
            ce => 'H',
            sr => \N__36763\
        );

    \ppm_encoder_1.init_pulses_RNO_1_0_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19938\,
            in1 => \N__23293\,
            in2 => \N__24386\,
            in3 => \N__30028\,
            lcout => \ppm_encoder_1.un1_init_pulses_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIC1OR2_2_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23294\,
            in1 => \N__20528\,
            in2 => \N__30087\,
            in3 => \N__19936\,
            lcout => \ppm_encoder_1.init_pulses_RNIC1OR2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_2_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23193\,
            in1 => \N__20122\,
            in2 => \N__19964\,
            in3 => \N__19952\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36023\,
            ce => 'H',
            sr => \N__36767\
        );

    \ppm_encoder_1.init_pulses_RNIG5OR2_6_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__23295\,
            in1 => \N__24622\,
            in2 => \N__30088\,
            in3 => \N__19937\,
            lcout => \ppm_encoder_1.init_pulses_RNIG5OR2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_6_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23194\,
            in1 => \N__20123\,
            in2 => \N__19883\,
            in3 => \N__19868\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36023\,
            ce => 'H',
            sr => \N__36767\
        );

    \ppm_encoder_1.init_pulses_RNIERUS_6_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__30027\,
            in1 => \N__24621\,
            in2 => \_gnd_net_\,
            in3 => \N__23030\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNI8LUS_0_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__23029\,
            in1 => \N__24381\,
            in2 => \_gnd_net_\,
            in3 => \N__30026\,
            lcout => \ppm_encoder_1.un1_init_pulses_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_16_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__20105\,
            in2 => \N__19811\,
            in3 => \N__19799\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36018\,
            ce => 'H',
            sr => \N__36770\
        );

    \ppm_encoder_1.init_pulses_4_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20106\,
            in1 => \N__19793\,
            in2 => \N__23191\,
            in3 => \N__19787\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36018\,
            ce => 'H',
            sr => \N__36770\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_4_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20136\,
            in1 => \N__23076\,
            in2 => \_gnd_net_\,
            in3 => \N__30035\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNICPUS_0_4_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__30036\,
            in1 => \_gnd_net_\,
            in2 => \N__23090\,
            in3 => \N__20137\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_4_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__20138\,
            in1 => \N__27924\,
            in2 => \N__30584\,
            in3 => \N__26648\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_5_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__20107\,
            in1 => \N__20027\,
            in2 => \N__23192\,
            in3 => \N__20021\,
            lcout => \ppm_encoder_1.init_pulsesZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36018\,
            ce => 'H',
            sr => \N__36770\
        );

    \ppm_encoder_1.PPM_STATE_RNISH5F_1_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36877\,
            lcout => \ppm_encoder_1.N_1014_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNITGRP_0_14_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__23087\,
            in1 => \N__24301\,
            in2 => \_gnd_net_\,
            in3 => \N__30041\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIE3D21_3_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25296\,
            in1 => \N__22504\,
            in2 => \N__27923\,
            in3 => \N__25238\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_159_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_11_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27894\,
            in1 => \N__23338\,
            in2 => \_gnd_net_\,
            in3 => \N__21476\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_11_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__30607\,
            in1 => \_gnd_net_\,
            in2 => \N__19982\,
            in3 => \N__30569\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIRERP_0_12_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__30040\,
            in1 => \_gnd_net_\,
            in2 => \N__27839\,
            in3 => \N__23086\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_2_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__30608\,
            in1 => \N__27895\,
            in2 => \N__20537\,
            in3 => \N__30570\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_e_0_6_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30989\,
            in2 => \_gnd_net_\,
            in3 => \N__21634\,
            lcout => alt_kp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36160\,
            ce => \N__25755\,
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_alt_kp_4_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__20485\,
            in1 => \N__33644\,
            in2 => \N__28187\,
            in3 => \N__31690\,
            lcout => alt_kp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36146\,
            ce => 'H',
            sr => \N__36690\
        );

    \pid_alt.error_i_reg_esr_6_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20471\,
            lcout => \pid_alt.error_i_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36142\,
            ce => \N__20300\,
            sr => \N__21570\
        );

    \pid_alt.error_p_reg_esr_RNI69J71_6_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__20459\,
            in1 => \N__20421\,
            in2 => \_gnd_net_\,
            in3 => \N__20399\,
            lcout => \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6\,
            ltout => \pid_alt.error_p_reg_esr_RNI69J71Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNIFL6F2_7_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20263\,
            in1 => \N__20238\,
            in2 => \N__20342\,
            in3 => \N__20224\,
            lcout => \pid_alt.error_p_reg_esr_RNIFL6F2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_i_reg_esr_7_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \pid_alt.error_i_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36142\,
            ce => \N__20300\,
            sr => \N__21570\
        );

    \pid_alt.error_p_reg_esr_RNI9CJ71_7_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__20264\,
            in1 => \N__20239\,
            in2 => \_gnd_net_\,
            in3 => \N__20225\,
            lcout => \pid_alt.error_p_reg_esr_RNI9CJ71Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_11_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26009\,
            lcout => \dron_frame_decoder_1.drone_altitude_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36137\,
            ce => \N__25636\,
            sr => \N__36696\
        );

    \dron_frame_decoder_1.source_Altitude_esr_9_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26089\,
            lcout => \dron_frame_decoder_1.drone_altitude_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36137\,
            ce => \N__25636\,
            sr => \N__36696\
        );

    \dron_frame_decoder_1.source_Altitude_esr_10_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26051\,
            lcout => \dron_frame_decoder_1.drone_altitude_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36137\,
            ce => \N__25636\,
            sr => \N__36696\
        );

    \dron_frame_decoder_1.source_Altitude_esr_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26126\,
            lcout => \dron_frame_decoder_1.drone_altitude_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36137\,
            ce => \N__25636\,
            sr => \N__36696\
        );

    \dron_frame_decoder_1.source_Altitude_esr_14_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26231\,
            lcout => drone_altitude_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36137\,
            ce => \N__25636\,
            sr => \N__36696\
        );

    \dron_frame_decoder_1.source_Altitude_esr_2_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26046\,
            lcout => drone_altitude_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36133\,
            ce => \N__25704\,
            sr => \N__36702\
        );

    \dron_frame_decoder_1.source_Altitude_esr_5_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26260\,
            lcout => \dron_frame_decoder_1.drone_altitude_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36133\,
            ce => \N__25704\,
            sr => \N__36702\
        );

    \dron_frame_decoder_1.source_Altitude_esr_3_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26005\,
            lcout => drone_altitude_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36133\,
            ce => \N__25704\,
            sr => \N__36702\
        );

    \pid_alt.error_p_reg_esr_RNIF43K_18_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20622\,
            in2 => \_gnd_net_\,
            in3 => \N__20572\,
            lcout => \pid_alt.error_p_reg_esr_RNIF43KZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.error_p_reg_esr_RNI1O4K_20_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20861\,
            in2 => \_gnd_net_\,
            in3 => \N__20803\,
            lcout => \pid_alt.error_p_reg_esr_RNI1O4KZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH2data_esr_0_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31475\,
            lcout => \frame_decoder_CH2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_2_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30867\,
            lcout => \frame_decoder_CH2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_3_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31199\,
            lcout => \frame_decoder_CH2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_4_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31691\,
            lcout => \frame_decoder_CH2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_5_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30737\,
            lcout => \frame_decoder_CH2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_esr_6_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \Commands_frame_decoder.source_CH2data_ess_7_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30988\,
            lcout => \frame_decoder_CH2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36123\,
            ce => \N__23555\,
            sr => \N__36708\
        );

    \scaler_2.un2_source_data_0_cry_1_c_RNO_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23804\,
            in1 => \N__21042\,
            in2 => \_gnd_net_\,
            in3 => \N__23762\,
            lcout => \scaler_2.un2_source_data_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.N_881_i_l_ofx_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21071\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23651\,
            lcout => \scaler_2.N_881_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un3_source_data_un3_source_data_0_axb_7_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__23650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21070\,
            lcout => \scaler_2.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_axb_7_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29087\,
            in2 => \_gnd_net_\,
            in3 => \N__29066\,
            lcout => \scaler_3.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.un2_source_data_0_cry_1_c_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21050\,
            in2 => \N__21043\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_6_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20992\,
            in2 => \N__21044\,
            in3 => \N__20999\,
            lcout => scaler_2_data_6,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_1\,
            carryout => \scaler_2.un2_source_data_0_cry_2\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_7_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20950\,
            in2 => \N__20996\,
            in3 => \N__20957\,
            lcout => scaler_2_data_7,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_2\,
            carryout => \scaler_2.un2_source_data_0_cry_3\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_8_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20929\,
            in2 => \N__20954\,
            in3 => \N__20936\,
            lcout => scaler_2_data_8,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_3\,
            carryout => \scaler_2.un2_source_data_0_cry_4\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_9_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21295\,
            in2 => \N__20933\,
            in3 => \N__20885\,
            lcout => scaler_2_data_9,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_4\,
            carryout => \scaler_2.un2_source_data_0_cry_5\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_10_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21274\,
            in2 => \N__21299\,
            in3 => \N__21281\,
            lcout => scaler_2_data_10,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_5\,
            carryout => \scaler_2.un2_source_data_0_cry_6\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_11_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21226\,
            in2 => \N__21278\,
            in3 => \N__21233\,
            lcout => scaler_2_data_11,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_6\,
            carryout => \scaler_2.un2_source_data_0_cry_7\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_12_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21208\,
            in2 => \N__21230\,
            in3 => \N__21212\,
            lcout => scaler_2_data_12,
            ltout => OPEN,
            carryin => \scaler_2.un2_source_data_0_cry_7\,
            carryout => \scaler_2.un2_source_data_0_cry_8\,
            clk => \N__36112\,
            ce => \N__29573\,
            sr => \N__36714\
        );

    \scaler_2.source_data_1_esr_13_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21209\,
            in2 => \N__21185\,
            in3 => \N__21170\,
            lcout => scaler_2_data_13,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \scaler_2.un2_source_data_0_cry_9\,
            clk => \N__36106\,
            ce => \N__29571\,
            sr => \N__36719\
        );

    \scaler_2.source_data_1_esr_14_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21167\,
            lcout => scaler_2_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36106\,
            ce => \N__29571\,
            sr => \N__36719\
        );

    \Commands_frame_decoder.source_alt_ki_7_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30987\,
            in2 => \_gnd_net_\,
            in3 => \N__21624\,
            lcout => alt_ki_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36098\,
            ce => \N__28041\,
            sr => \_gnd_net_\
        );

    \pid_alt.pid_prereg_1_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__34132\,
            in1 => \N__21137\,
            in2 => \N__21119\,
            in3 => \N__21097\,
            lcout => \pid_alt.pid_preregZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36091\,
            ce => 'H',
            sr => \N__36727\
        );

    \pid_alt.source_data_valid_esr_RNO_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34131\,
            in2 => \_gnd_net_\,
            in3 => \N__36895\,
            lcout => \pid_alt.state_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_1_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34133\,
            lcout => \pid_alt.N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36091\,
            ce => 'H',
            sr => \N__36727\
        );

    \pid_alt.state_RNICP2N1_0_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23825\,
            in2 => \_gnd_net_\,
            in3 => \N__21623\,
            lcout => \pid_alt.N_422_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.source_data_valid_esr_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23885\,
            lcout => pid_altitude_dv,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36083\,
            ce => \N__21482\,
            sr => \N__36730\
        );

    \ppm_encoder_1.elevator_13_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__24419\,
            in1 => \N__29657\,
            in2 => \N__24936\,
            in3 => \N__24328\,
            lcout => \ppm_encoder_1.elevatorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.rudder_11_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__26908\,
            in1 => \N__24858\,
            in2 => \N__25529\,
            in3 => \N__21468\,
            lcout => \ppm_encoder_1.rudderZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.rudder_7_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__25595\,
            in1 => \N__26566\,
            in2 => \N__24937\,
            in3 => \N__21432\,
            lcout => \ppm_encoder_1.rudderZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.throttle_10_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__21416\,
            in1 => \N__24859\,
            in2 => \N__21386\,
            in3 => \N__22599\,
            lcout => \ppm_encoder_1.throttleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.throttle_13_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__21371\,
            in1 => \N__21350\,
            in2 => \N__24938\,
            in3 => \N__23689\,
            lcout => \ppm_encoder_1.throttleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.throttle_2_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111101101001000"
        )
    port map (
            in0 => \N__21338\,
            in1 => \N__24860\,
            in2 => \N__21326\,
            in3 => \N__22764\,
            lcout => \ppm_encoder_1.throttleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.throttle_4_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21815\,
            in1 => \N__21800\,
            in2 => \N__24939\,
            in3 => \N__21843\,
            lcout => \ppm_encoder_1.throttleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36075\,
            ce => 'H',
            sr => \N__36736\
        );

    \ppm_encoder_1.throttle_RNII6JI2_12_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__21648\,
            in1 => \N__27789\,
            in2 => \N__22359\,
            in3 => \N__22251\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNIFQRT5_12_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21788\,
            in2 => \N__21770\,
            in3 => \N__21752\,
            lcout => \ppm_encoder_1.elevator_RNIFQRT5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNI25DH2_12_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__21696\,
            in1 => \N__21708\,
            in2 => \N__22124\,
            in3 => \N__22006\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_3_12_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29489\,
            in1 => \N__21649\,
            in2 => \_gnd_net_\,
            in3 => \N__21697\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_12_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29223\,
            in1 => \_gnd_net_\,
            in2 => \N__21746\,
            in3 => \N__21709\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_12_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__21710\,
            in1 => \N__24929\,
            in2 => \N__21743\,
            in3 => \N__21719\,
            lcout => \ppm_encoder_1.aileronZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36064\,
            ce => 'H',
            sr => \N__36740\
        );

    \ppm_encoder_1.elevator_12_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__21698\,
            in1 => \N__29705\,
            in2 => \N__24983\,
            in3 => \N__24428\,
            lcout => \ppm_encoder_1.elevatorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36064\,
            ce => 'H',
            sr => \N__36740\
        );

    \ppm_encoder_1.throttle_12_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21686\,
            in1 => \N__21662\,
            in2 => \N__24984\,
            in3 => \N__21650\,
            lcout => \ppm_encoder_1.throttleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36064\,
            ce => 'H',
            sr => \N__36740\
        );

    \ppm_encoder_1.throttle_RNIS5KK2_8_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__24225\,
            in1 => \N__21882\,
            in2 => \N__22343\,
            in3 => \N__22250\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.un2_throttle_iv_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_RNIONI96_8_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__22163\,
            in1 => \_gnd_net_\,
            in2 => \N__22148\,
            in3 => \N__21944\,
            lcout => \ppm_encoder_1.throttle_RNIONI96Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_RNICKVN2_8_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__21936\,
            in1 => \N__22791\,
            in2 => \N__22110\,
            in3 => \N__22000\,
            lcout => \ppm_encoder_1.un2_throttle_iv_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_8_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21883\,
            in1 => \N__29480\,
            in2 => \_gnd_net_\,
            in3 => \N__21937\,
            lcout => \ppm_encoder_1.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_8_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101011001010"
        )
    port map (
            in0 => \N__21938\,
            in1 => \N__24476\,
            in2 => \N__24982\,
            in3 => \N__28943\,
            lcout => \ppm_encoder_1.elevatorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36056\,
            ce => 'H',
            sr => \N__36745\
        );

    \ppm_encoder_1.throttle_8_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111011100010"
        )
    port map (
            in0 => \N__21884\,
            in1 => \N__24921\,
            in2 => \N__21926\,
            in3 => \N__21893\,
            lcout => \ppm_encoder_1.throttleZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36056\,
            ce => 'H',
            sr => \N__36745\
        );

    \ppm_encoder_1.aileron_8_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__21872\,
            in1 => \N__21854\,
            in2 => \N__24981\,
            in3 => \N__22792\,
            lcout => \ppm_encoder_1.aileronZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36056\,
            ce => 'H',
            sr => \N__36745\
        );

    \ppm_encoder_1.rudder_8_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011001100"
        )
    port map (
            in0 => \N__25577\,
            in1 => \N__24226\,
            in2 => \N__26525\,
            in3 => \N__24928\,
            lcout => \ppm_encoder_1.rudderZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36056\,
            ce => 'H',
            sr => \N__36745\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_4_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26678\,
            in1 => \N__21845\,
            in2 => \_gnd_net_\,
            in3 => \N__22483\,
            lcout => \ppm_encoder_1.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_0_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111111100"
        )
    port map (
            in0 => \N__23046\,
            in1 => \N__22544\,
            in2 => \N__36914\,
            in3 => \N__29967\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011011110"
        )
    port map (
            in0 => \N__29963\,
            in1 => \N__36901\,
            in2 => \N__29252\,
            in3 => \N__23047\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_1_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__36900\,
            in1 => \N__29218\,
            in2 => \N__22528\,
            in3 => \N__29966\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_3_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__29962\,
            in1 => \N__22640\,
            in2 => \N__22451\,
            in3 => \N__36909\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_1_rep1_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__22484\,
            in1 => \N__29217\,
            in2 => \N__36913\,
            in3 => \N__29965\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_0_rep1_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000110"
        )
    port map (
            in0 => \N__29964\,
            in1 => \N__25279\,
            in2 => \N__23083\,
            in3 => \N__36902\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNILS7D_3_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22574\,
            in2 => \_gnd_net_\,
            in3 => \N__22446\,
            lcout => \ppm_encoder_1.N_227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m9_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110000000"
        )
    port map (
            in0 => \N__27955\,
            in1 => \N__29482\,
            in2 => \N__29222\,
            in3 => \N__25225\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1_0_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22432\,
            in1 => \N__22942\,
            in2 => \_gnd_net_\,
            in3 => \N__22401\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_fast_RNI35QO1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI2APU1_2_1_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22658\,
            in3 => \N__29908\,
            lcout => \ppm_encoder_1.PPM_STATE_RNI2APU1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_3_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__29910\,
            in1 => \N__22639\,
            in2 => \N__25236\,
            in3 => \N__36911\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_11_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22943\,
            in1 => \N__23339\,
            in2 => \_gnd_net_\,
            in3 => \N__29909\,
            lcout => \ppm_encoder_1.un1_init_pulses_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_10_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29481\,
            in1 => \N__22607\,
            in2 => \_gnd_net_\,
            in3 => \N__24107\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_10_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29181\,
            in1 => \_gnd_net_\,
            in2 => \N__22580\,
            in3 => \N__24164\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_fast_2_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__29911\,
            in1 => \N__35063\,
            in2 => \N__23384\,
            in3 => \N__22577\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36042\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIUS1G_4_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27422\,
            in1 => \N__27451\,
            in2 => \N__27398\,
            in3 => \N__27481\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIDBJ8_13_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30437\,
            in2 => \_gnd_net_\,
            in3 => \N__27605\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_17_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIAEV01_8_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__22553\,
            in1 => \N__27635\,
            in2 => \N__22547\,
            in3 => \N__27371\,
            lcout => \ppm_encoder_1.N_145_17\,
            ltout => \ppm_encoder_1.N_145_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_1_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30176\,
            in1 => \N__24680\,
            in2 => \N__22727\,
            in3 => \N__25142\,
            lcout => \ppm_encoder_1.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_RNI09RH2_1_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30175\,
            in1 => \N__24746\,
            in2 => \N__22724\,
            in3 => \N__25141\,
            lcout => \ppm_encoder_1.N_238\,
            ltout => \ppm_encoder_1.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_0_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__25334\,
            in1 => \N__25396\,
            in2 => \N__22715\,
            in3 => \N__24740\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36034\,
            ce => 'H',
            sr => \N__36758\
        );

    \ppm_encoder_1.PPM_STATE_RNIV4V5_1_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24737\,
            in2 => \_gnd_net_\,
            in3 => \N__25333\,
            lcout => \ppm_encoder_1.PPM_STATE_59_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_RNO_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22694\,
            in1 => \N__27452\,
            in2 => \N__22667\,
            in3 => \N__27482\,
            lcout => \ppm_encoder_1.counter24_0_I_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_4_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22712\,
            in1 => \N__22700\,
            in2 => \_gnd_net_\,
            in3 => \N__27110\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.pulses2count_esr_5_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__22688\,
            in1 => \N__22679\,
            in2 => \N__27122\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.pulses2count_esr_0_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24491\,
            in1 => \N__27111\,
            in2 => \_gnd_net_\,
            in3 => \N__24344\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.pulses2count_esr_1_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27109\,
            in1 => \N__25100\,
            in2 => \_gnd_net_\,
            in3 => \N__23348\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.pulses2count_esr_10_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22862\,
            in1 => \N__27112\,
            in2 => \_gnd_net_\,
            in3 => \N__25424\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.counter24_0_I_33_c_RNO_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__22853\,
            in1 => \N__27694\,
            in2 => \N__22817\,
            in3 => \N__27661\,
            lcout => \ppm_encoder_1.counter24_0_I_33_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_11_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22847\,
            in1 => \N__27113\,
            in2 => \_gnd_net_\,
            in3 => \N__22829\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36024\,
            ce => \N__27014\,
            sr => \N__36760\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_8_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29260\,
            in1 => \N__22808\,
            in2 => \_gnd_net_\,
            in3 => \N__22796\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_8_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27107\,
            in2 => \N__22778\,
            in3 => \N__24212\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36019\,
            ce => \N__26997\,
            sr => \N__36764\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_2_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__29259\,
            in1 => \N__29461\,
            in2 => \_gnd_net_\,
            in3 => \N__22775\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_2_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27106\,
            in2 => \N__22748\,
            in3 => \N__22745\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36019\,
            ce => \N__26997\,
            sr => \N__36764\
        );

    \ppm_encoder_1.pulses2count_esr_3_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27105\,
            in1 => \N__23096\,
            in2 => \_gnd_net_\,
            in3 => \N__25163\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36019\,
            ce => \N__26997\,
            sr => \N__36764\
        );

    \ppm_encoder_1.counter24_0_I_27_c_RNO_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__22733\,
            in1 => \N__27730\,
            in2 => \N__23393\,
            in3 => \N__27367\,
            lcout => \ppm_encoder_1.counter24_0_I_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_9_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29261\,
            in1 => \N__23441\,
            in2 => \_gnd_net_\,
            in3 => \N__23429\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_9_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27108\,
            in2 => \N__23408\,
            in3 => \N__23405\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36019\,
            ce => \N__26997\,
            sr => \N__36764\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_ns_3_0__m6_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__23081\,
            in1 => \N__29273\,
            in2 => \N__29484\,
            in3 => \N__27897\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2\,
            ltout => \ppm_encoder_1.CHOOSE_CHANNEL_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_2_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__27898\,
            in1 => \N__35078\,
            in2 => \N__23369\,
            in3 => \N__30039\,
            lcout => \ppm_encoder_1.CHOOSE_CHANNELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_1_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__30531\,
            in1 => \N__27896\,
            in2 => \N__30618\,
            in3 => \N__23366\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIQDRP_0_11_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__23337\,
            in1 => \N__23080\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNIGD613_3_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30038\,
            in1 => \N__30112\,
            in2 => \_gnd_net_\,
            in3 => \N__23297\,
            lcout => \ppm_encoder_1.un1_init_pulses_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_3_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__29272\,
            in1 => \N__29460\,
            in2 => \_gnd_net_\,
            in3 => \N__24773\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.init_pulses_RNIVIRP_16_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__30390\,
            in1 => \N__23082\,
            in2 => \_gnd_net_\,
            in3 => \N__30043\,
            lcout => \ppm_encoder_1.un1_init_pulses_3_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_3_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__25297\,
            in1 => \N__29392\,
            in2 => \_gnd_net_\,
            in3 => \N__25237\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_10_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__34129\,
            in1 => \N__23996\,
            in2 => \_gnd_net_\,
            in3 => \N__23956\,
            lcout => \pid_alt.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36143\,
            ce => 'H',
            sr => \N__36689\
        );

    \dron_frame_decoder_1.source_Altitude_esr_6_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26229\,
            lcout => \dron_frame_decoder_1.drone_altitude_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36138\,
            ce => \N__25705\,
            sr => \N__36691\
        );

    \dron_frame_decoder_1.source_Altitude_esr_4_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25964\,
            lcout => \dron_frame_decoder_1.drone_altitude_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36138\,
            ce => \N__25705\,
            sr => \N__36691\
        );

    \Commands_frame_decoder.source_CH1data8lto7_1_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30969\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \Commands_frame_decoder.state_ns_i_a2_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIHIDC_4_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23501\,
            lcout => drone_altitude_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIIJDC_5_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23486\,
            lcout => drone_altitude_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_Altitude_esr_RNIJKDC_6_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23471\,
            lcout => drone_altitude_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH1data_esr_4_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31696\,
            lcout => alt_command_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36128\,
            ce => \N__25877\,
            sr => \N__36697\
        );

    \Commands_frame_decoder.source_CH1data_esr_5_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30738\,
            lcout => alt_command_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36128\,
            ce => \N__25877\,
            sr => \N__36697\
        );

    \Commands_frame_decoder.source_CH1data_esr_6_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31362\,
            lcout => alt_command_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36128\,
            ce => \N__25877\,
            sr => \N__36697\
        );

    \Commands_frame_decoder.source_CH1data_esr_7_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30983\,
            lcout => alt_command_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36128\,
            ce => \N__25877\,
            sr => \N__36697\
        );

    \Commands_frame_decoder.state_RNIC08S_3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__36889\,
            in1 => \N__28148\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIG48S_7_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36888\,
            in2 => \_gnd_net_\,
            in3 => \N__28268\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset2data_esr_0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31474\,
            lcout => \frame_decoder_OFF2data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_1_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31822\,
            lcout => \frame_decoder_OFF2data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_2_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30857\,
            lcout => \frame_decoder_OFF2data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF2data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_4_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31695\,
            lcout => \frame_decoder_OFF2data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_5_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30736\,
            lcout => \frame_decoder_OFF2data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_esr_6_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31343\,
            lcout => \frame_decoder_OFF2data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \Commands_frame_decoder.source_offset2data_ess_7_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30982\,
            lcout => \frame_decoder_OFF2data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36118\,
            ce => \N__23642\,
            sr => \N__36706\
        );

    \dron_frame_decoder_1.state_RNO_2_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__25911\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24063\,
            lcout => \dron_frame_decoder_1.state_ns_i_i_a2_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNO_1_0_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25912\,
            in1 => \N__24064\,
            in2 => \N__24029\,
            in3 => \N__32421\,
            lcout => \dron_frame_decoder_1.state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_data_valid_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__36942\,
            in1 => \N__33628\,
            in2 => \N__32813\,
            in3 => \N__31892\,
            lcout => \debug_CH3_20A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36107\,
            ce => 'H',
            sr => \N__36712\
        );

    \dron_frame_decoder_1.state_0_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__24065\,
            in1 => \N__32186\,
            in2 => \N__23627\,
            in3 => \N__23597\,
            lcout => \dron_frame_decoder_1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36107\,
            ce => 'H',
            sr => \N__36712\
        );

    \dron_frame_decoder_1.source_data_valid_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__25916\,
            in1 => \N__32422\,
            in2 => \_gnd_net_\,
            in3 => \N__23981\,
            lcout => \debug_CH1_0A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36107\,
            ce => 'H',
            sr => \N__36712\
        );

    \dron_frame_decoder_1.state_RNO_0_0_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__24040\,
            in2 => \N__23609\,
            in3 => \N__23704\,
            lcout => \dron_frame_decoder_1.state_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1_1_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25958\,
            in2 => \_gnd_net_\,
            in3 => \N__26081\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_0_0_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNIN9KQ1_0_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26225\,
            in1 => \N__24062\,
            in2 => \N__24044\,
            in3 => \N__26004\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_1_3_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26118\,
            in1 => \N__32416\,
            in2 => \N__26050\,
            in3 => \N__24002\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3\,
            ltout => \dron_frame_decoder_1.state_ns_0_i_a2_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_1_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__24024\,
            in1 => \N__24041\,
            in2 => \N__24032\,
            in3 => \N__32174\,
            lcout => \dron_frame_decoder_1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36099\,
            ce => 'H',
            sr => \N__36715\
        );

    \dron_frame_decoder_1.state_ns_0_i_a2_1_0_3_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26178\,
            in2 => \_gnd_net_\,
            in3 => \N__26259\,
            lcout => \dron_frame_decoder_1.state_ns_0_i_a2_1_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pid_alt.state_RNIFCSD1_0_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__23985\,
            in1 => \N__23867\,
            in2 => \N__34130\,
            in3 => \N__36875\,
            lcout => \pid_alt.state_RNIFCSD1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_4_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__36958\,
            in1 => \N__23819\,
            in2 => \N__23737\,
            in3 => \N__23779\,
            lcout => scaler_2_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36084\,
            ce => 'H',
            sr => \N__36724\
        );

    \dron_frame_decoder_1.state_3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32161\,
            in1 => \N__23720\,
            in2 => \N__32206\,
            in3 => \N__23708\,
            lcout => \dron_frame_decoder_1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36084\,
            ce => 'H',
            sr => \N__36724\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_13_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29485\,
            in1 => \N__23688\,
            in2 => \_gnd_net_\,
            in3 => \N__24327\,
            lcout => \ppm_encoder_1.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_14_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__27958\,
            in1 => \N__30568\,
            in2 => \N__24308\,
            in3 => \N__25777\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_8_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__30567\,
            in1 => \N__24266\,
            in2 => \N__24236\,
            in3 => \N__27959\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_12_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__26869\,
            in1 => \N__25508\,
            in2 => \N__27799\,
            in3 => \N__24879\,
            lcout => \ppm_encoder_1.rudderZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36065\,
            ce => 'H',
            sr => \N__36731\
        );

    \ppm_encoder_1.aileron_10_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__24200\,
            in1 => \N__24176\,
            in2 => \N__24940\,
            in3 => \N__24153\,
            lcout => \ppm_encoder_1.aileronZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36065\,
            ce => 'H',
            sr => \N__36731\
        );

    \ppm_encoder_1.aileron_13_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__24137\,
            in1 => \N__24116\,
            in2 => \N__24942\,
            in3 => \N__29523\,
            lcout => \ppm_encoder_1.aileronZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36065\,
            ce => 'H',
            sr => \N__36731\
        );

    \ppm_encoder_1.elevator_10_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110111101100000"
        )
    port map (
            in0 => \N__28868\,
            in1 => \N__24449\,
            in2 => \N__24941\,
            in3 => \N__24096\,
            lcout => \ppm_encoder_1.elevatorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36065\,
            ce => 'H',
            sr => \N__36731\
        );

    \ppm_encoder_1.un1_elevator_cry_6_c_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29023\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \ppm_encoder_1.un1_elevator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_6_THRU_LUT4_0_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28978\,
            in2 => \_gnd_net_\,
            in3 => \N__24068\,
            lcout => \ppm_encoder_1.un1_elevator_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_6\,
            carryout => \ppm_encoder_1.un1_elevator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_7_THRU_LUT4_0_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28939\,
            in2 => \_gnd_net_\,
            in3 => \N__24470\,
            lcout => \ppm_encoder_1.un1_elevator_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_7\,
            carryout => \ppm_encoder_1.un1_elevator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_8_THRU_LUT4_0_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28903\,
            in2 => \_gnd_net_\,
            in3 => \N__24452\,
            lcout => \ppm_encoder_1.un1_elevator_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_8\,
            carryout => \ppm_encoder_1.un1_elevator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_9_THRU_LUT4_0_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28864\,
            in2 => \_gnd_net_\,
            in3 => \N__24443\,
            lcout => \ppm_encoder_1.un1_elevator_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_9\,
            carryout => \ppm_encoder_1.un1_elevator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_10_THRU_LUT4_0_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29737\,
            in2 => \_gnd_net_\,
            in3 => \N__24431\,
            lcout => \ppm_encoder_1.un1_elevator_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_10\,
            carryout => \ppm_encoder_1.un1_elevator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_11_THRU_LUT4_0_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29704\,
            in2 => \_gnd_net_\,
            in3 => \N__24422\,
            lcout => \ppm_encoder_1.un1_elevator_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_11\,
            carryout => \ppm_encoder_1.un1_elevator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_elevator_cry_12_THRU_LUT4_0_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29656\,
            in2 => \N__28674\,
            in3 => \N__24413\,
            lcout => \ppm_encoder_1.un1_elevator_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_elevator_cry_12\,
            carryout => \ppm_encoder_1.un1_elevator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.elevator_esr_14_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29627\,
            in2 => \_gnd_net_\,
            in3 => \N__24410\,
            lcout => \ppm_encoder_1.elevatorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36050\,
            ce => \N__27267\,
            sr => \N__36741\
        );

    \ppm_encoder_1.rudder_10_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011110000"
        )
    port map (
            in0 => \N__26431\,
            in1 => \N__25541\,
            in2 => \N__25455\,
            in3 => \N__24947\,
            lcout => \ppm_encoder_1.rudderZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36043\,
            ce => 'H',
            sr => \N__36746\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_0_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__27948\,
            in2 => \_gnd_net_\,
            in3 => \N__24385\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_ctle_14_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24943\,
            in2 => \_gnd_net_\,
            in3 => \N__36890\,
            lcout => \ppm_encoder_1.pid_altitude_dv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.aileron_6_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__24944\,
            in1 => \N__24656\,
            in2 => \_gnd_net_\,
            in3 => \N__29112\,
            lcout => \ppm_encoder_1.aileronZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36043\,
            ce => 'H',
            sr => \N__36746\
        );

    \ppm_encoder_1.elevator_6_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__29301\,
            in1 => \N__29027\,
            in2 => \_gnd_net_\,
            in3 => \N__24946\,
            lcout => \ppm_encoder_1.elevatorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36043\,
            ce => 'H',
            sr => \N__36746\
        );

    \ppm_encoder_1.rudder_6_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__24945\,
            in1 => \N__24606\,
            in2 => \_gnd_net_\,
            in3 => \N__26608\,
            lcout => \ppm_encoder_1.rudderZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36043\,
            ce => 'H',
            sr => \N__36746\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_6_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__27949\,
            in1 => \N__24632\,
            in2 => \N__24608\,
            in3 => \N__30557\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_13_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__27947\,
            in1 => \N__24587\,
            in2 => \N__24559\,
            in3 => \N__30545\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_13_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__24985\,
            in1 => \N__24555\,
            in2 => \N__26816\,
            in3 => \N__25802\,
            lcout => \ppm_encoder_1.rudderZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36035\,
            ce => 'H',
            sr => \N__36752\
        );

    \ppm_encoder_1.throttle_0_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__24508\,
            in1 => \N__24987\,
            in2 => \_gnd_net_\,
            in3 => \N__24536\,
            lcout => \ppm_encoder_1.throttleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36035\,
            ce => 'H',
            sr => \N__36752\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_0_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__29195\,
            in1 => \N__29466\,
            in2 => \_gnd_net_\,
            in3 => \N__24507\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_1_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__29467\,
            in1 => \N__29196\,
            in2 => \_gnd_net_\,
            in3 => \N__25053\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.throttle_1_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__24986\,
            in1 => \N__25054\,
            in2 => \N__25091\,
            in3 => \N__25076\,
            lcout => \ppm_encoder_1.throttleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36035\,
            ce => 'H',
            sr => \N__36752\
        );

    \ppm_encoder_1.throttle_3_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__25034\,
            in1 => \N__25022\,
            in2 => \N__25000\,
            in3 => \N__24768\,
            lcout => \ppm_encoder_1.throttleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36035\,
            ce => 'H',
            sr => \N__36752\
        );

    \ppm_encoder_1.PPM_STATE_RNISL0F_1_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27505\,
            in1 => \N__24738\,
            in2 => \N__27563\,
            in3 => \N__27531\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.PPM_STATE_1_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25358\,
            in2 => \_gnd_net_\,
            in3 => \N__25411\,
            lcout => \ppm_encoder_1.PPM_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36025\,
            ce => 'H',
            sr => \N__36755\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_0_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__25357\,
            in1 => \N__25395\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_140_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.ppm_output_reg_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011110100"
        )
    port map (
            in0 => \N__24739\,
            in1 => \N__24691\,
            in2 => \N__24719\,
            in3 => \N__24716\,
            lcout => ppm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36025\,
            ce => 'H',
            sr => \N__36755\
        );

    \ppm_encoder_1.ppm_output_reg_RNO_2_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27506\,
            in1 => \N__27562\,
            in2 => \N__25363\,
            in3 => \N__27532\,
            lcout => \ppm_encoder_1.un1_PPM_STATE_1_sqmuxa_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_RNO_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__24674\,
            in1 => \N__24665\,
            in2 => \N__27533\,
            in3 => \N__27504\,
            lcout => \ppm_encoder_1.counter24_0_I_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_RNO_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__27558\,
            in1 => \N__25157\,
            in2 => \N__25151\,
            in3 => \N__26944\,
            lcout => \ppm_encoder_1.counter24_0_I_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNIK1KG_0_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26945\,
            in1 => \N__27698\,
            in2 => \N__27668\,
            in3 => \N__27731\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_1_c_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25133\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_9_c_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28686\,
            in2 => \N__25127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_0\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_15_c_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25118\,
            in2 => \N__28700\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_1\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_21_c_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28678\,
            in2 => \N__27239\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_2\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_27_c_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25112\,
            in2 => \N__28701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_3\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_33_c_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25106\,
            in2 => \N__28658\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_4\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_39_c_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27152\,
            in2 => \N__28702\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_5\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28685\,
            in2 => \N__30413\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_6\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25601\,
            in2 => \N__28672\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_28_0_\,
            carryout => \ppm_encoder_1.counter24_0_data_tmp_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30263\,
            in2 => \N__28703\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ppm_encoder_1.counter24_0_data_tmp_8\,
            carryout => \ppm_encoder_1.counter24_0_N_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_N_2_THRU_LUT4_0_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25493\,
            lcout => \ppm_encoder_1.counter24_0_N_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_10_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__27925\,
            in1 => \N__25489\,
            in2 => \N__25460\,
            in3 => \N__30533\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNIGCO83_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__25412\,
            in1 => \N__25382\,
            in2 => \N__25364\,
            in3 => \N__35059\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNIGCOZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.CHOOSE_CHANNEL_RNI33GU_0_3_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29427\,
            in1 => \N__25292\,
            in2 => \_gnd_net_\,
            in3 => \N__25229\,
            lcout => \ppm_encoder_1.pulses2count_9_sn_N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_3_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__30532\,
            in1 => \N__27926\,
            in2 => \N__30626\,
            in3 => \N__25190\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_51_c_RNO_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__30236\,
            in1 => \N__30214\,
            in2 => \N__30329\,
            in3 => \N__30371\,
            lcout => \ppm_encoder_1.counter24_0_I_51_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_c_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26609\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_29_0_\,
            carryout => \ppm_encoder_1.un1_rudder_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_6_THRU_LUT4_0_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26567\,
            in2 => \_gnd_net_\,
            in3 => \N__25580\,
            lcout => \ppm_encoder_1.un1_rudder_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_6\,
            carryout => \ppm_encoder_1.un1_rudder_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_7_THRU_LUT4_0_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26524\,
            in2 => \_gnd_net_\,
            in3 => \N__25562\,
            lcout => \ppm_encoder_1.un1_rudder_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_7\,
            carryout => \ppm_encoder_1.un1_rudder_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_8_THRU_LUT4_0_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26473\,
            in2 => \_gnd_net_\,
            in3 => \N__25544\,
            lcout => \ppm_encoder_1.un1_rudder_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_8\,
            carryout => \ppm_encoder_1.un1_rudder_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_9_THRU_LUT4_0_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26432\,
            in2 => \_gnd_net_\,
            in3 => \N__25532\,
            lcout => \ppm_encoder_1.un1_rudder_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_9\,
            carryout => \ppm_encoder_1.un1_rudder_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_10_THRU_LUT4_0_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26912\,
            in2 => \_gnd_net_\,
            in3 => \N__25511\,
            lcout => \ppm_encoder_1.un1_rudder_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_10\,
            carryout => \ppm_encoder_1.un1_rudder_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_11_THRU_LUT4_0_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26870\,
            in2 => \_gnd_net_\,
            in3 => \N__25496\,
            lcout => \ppm_encoder_1.un1_rudder_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_11\,
            carryout => \ppm_encoder_1.un1_rudder_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.un1_rudder_cry_12_THRU_LUT4_0_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26815\,
            in2 => \N__28673\,
            in3 => \N__25790\,
            lcout => \ppm_encoder_1.un1_rudder_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_rudder_cry_12\,
            carryout => \ppm_encoder_1.un1_rudder_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.rudder_esr_14_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26786\,
            in2 => \_gnd_net_\,
            in3 => \N__25787\,
            lcout => \ppm_encoder_1.rudderZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36010\,
            ce => \N__27293\,
            sr => \N__36768\
        );

    \Commands_frame_decoder.state_RNIF38S_6_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__28177\,
            in1 => \N__33643\,
            in2 => \_gnd_net_\,
            in3 => \N__36887\,
            lcout => \Commands_frame_decoder.state_RNIF38SZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_offset4data_esr_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31223\,
            lcout => \frame_decoder_OFF4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36129\,
            ce => \N__28111\,
            sr => \N__36692\
        );

    \dron_frame_decoder_1.state_RNI0TLI1_5_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__28079\,
            in1 => \N__28240\,
            in2 => \N__25910\,
            in3 => \N__36882\,
            lcout => \dron_frame_decoder_1.N_390_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__32413\,
            in1 => \N__28241\,
            in2 => \N__28099\,
            in3 => \N__32187\,
            lcout => \dron_frame_decoder_1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36124\,
            ce => 'H',
            sr => \N__36694\
        );

    \dron_frame_decoder_1.state_RNI3T3K1_7_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28239\,
            in1 => \N__25897\,
            in2 => \N__25618\,
            in3 => \N__28078\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.state_RNI3T3K1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI0AAT1_7_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25655\,
            in3 => \N__35075\,
            lcout => \dron_frame_decoder_1.N_382_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32415\,
            in1 => \N__25617\,
            in2 => \N__28100\,
            in3 => \N__32189\,
            lcout => \dron_frame_decoder_1.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36124\,
            ce => 'H',
            sr => \N__36694\
        );

    \dron_frame_decoder_1.state_6_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__32188\,
            in1 => \N__25901\,
            in2 => \N__25619\,
            in3 => \N__32414\,
            lcout => \dron_frame_decoder_1.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36124\,
            ce => 'H',
            sr => \N__36694\
        );

    \Commands_frame_decoder.state_RNIBV7S_2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25828\,
            in2 => \_gnd_net_\,
            in3 => \N__36891\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__25862\,
            in1 => \N__31106\,
            in2 => \N__25856\,
            in3 => \N__32881\,
            lcout => \Commands_frame_decoder.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36119\,
            ce => 'H',
            sr => \N__36698\
        );

    \Commands_frame_decoder.state_RNO_1_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31449\,
            in2 => \_gnd_net_\,
            in3 => \N__30945\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_2_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30852\,
            in1 => \N__31088\,
            in2 => \N__25865\,
            in3 => \N__30711\,
            lcout => \Commands_frame_decoder.state_ns_0_a3_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIEI1J_2_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25852\,
            in2 => \_gnd_net_\,
            in3 => \N__33631\,
            lcout => \Commands_frame_decoder.un1_sink_data_valid_2_0\,
            ltout => \Commands_frame_decoder.un1_sink_data_valid_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_3_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25814\,
            in2 => \N__25817\,
            in3 => \N__32882\,
            lcout => \Commands_frame_decoder.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36119\,
            ce => 'H',
            sr => \N__36698\
        );

    \Commands_frame_decoder.state_RNIFJ1J_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33563\,
            lcout => \Commands_frame_decoder.source_CH2data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNID18S_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28216\,
            in2 => \_gnd_net_\,
            in3 => \N__36884\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIHL1J_5_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28204\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIE28S_5_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__36874\,
            in1 => \_gnd_net_\,
            in2 => \N__26144\,
            in3 => \_gnd_net_\,
            lcout => \Commands_frame_decoder.source_CH4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_reset_system_g_THRU_LUT4_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36873\,
            lcout => \GB_BUFFER_reset_system_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNIGK1J_4_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28132\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => \Commands_frame_decoder.source_CH3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_CH3data_esr_4_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31652\,
            lcout => \frame_decoder_CH3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36100\,
            ce => \N__28464\,
            sr => \N__36709\
        );

    \uart_drone.data_esr_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28321\,
            lcout => uart_drone_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28307\,
            lcout => uart_drone_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28291\,
            lcout => uart_drone_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28415\,
            lcout => uart_drone_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_4_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34226\,
            lcout => uart_drone_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28403\,
            lcout => uart_drone_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_6_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28390\,
            lcout => uart_drone_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \uart_drone.data_esr_7_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34409\,
            lcout => uart_drone_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36092\,
            ce => \N__31520\,
            sr => \N__31562\
        );

    \Commands_frame_decoder.source_offset4data_esr_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31491\,
            lcout => \frame_decoder_OFF4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_esr_1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31827\,
            lcout => \frame_decoder_OFF4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_esr_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30844\,
            lcout => \frame_decoder_OFF4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_esr_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31697\,
            lcout => \frame_decoder_OFF4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_esr_5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30716\,
            lcout => \frame_decoder_OFF4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_esr_6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31358\,
            lcout => \frame_decoder_OFF4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_offset4data_ess_7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30959\,
            lcout => \frame_decoder_OFF4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36085\,
            ce => \N__28121\,
            sr => \N__36716\
        );

    \Commands_frame_decoder.source_CH4data_esr_0_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31494\,
            lcout => \frame_decoder_CH4data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_1_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31828\,
            lcout => \frame_decoder_CH4data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_2_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30856\,
            lcout => \frame_decoder_CH4data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_3_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH4data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_4_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31670\,
            lcout => \frame_decoder_CH4data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_5_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30717\,
            lcout => \frame_decoder_CH4data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_esr_6_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31359\,
            lcout => \frame_decoder_CH4data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \Commands_frame_decoder.source_CH4data_ess_7_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30981\,
            lcout => \frame_decoder_CH4data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36076\,
            ce => \N__26291\,
            sr => \N__36720\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26696\,
            in2 => \N__26738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_0_c_RNI40BL_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26279\,
            in2 => \N__26273\,
            in3 => \N__26408\,
            lcout => \scaler_4.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_0\,
            carryout => \scaler_4.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_1_c_RNI74CL_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26405\,
            in2 => \N__26396\,
            in3 => \N__26387\,
            lcout => \scaler_4.un3_source_data_0_cry_1_c_RNI74CL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_1\,
            carryout => \scaler_4.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_2_c_RNIA8DL_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26384\,
            in2 => \N__26378\,
            in3 => \N__26366\,
            lcout => \scaler_4.un3_source_data_0_cry_2_c_RNIA8DL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_2\,
            carryout => \scaler_4.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_3_c_RNIDCEL_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26363\,
            in2 => \N__26354\,
            in3 => \N__26345\,
            lcout => \scaler_4.un3_source_data_0_cry_3_c_RNIDCEL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_3\,
            carryout => \scaler_4.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_4_c_RNIGGFL_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26342\,
            in2 => \N__26336\,
            in3 => \N__26324\,
            lcout => \scaler_4.un3_source_data_0_cry_4_c_RNIGGFL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_4\,
            carryout => \scaler_4.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_5_c_RNIJKGL_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26321\,
            in2 => \N__26315\,
            in3 => \N__26303\,
            lcout => \scaler_4.un3_source_data_0_cry_5_c_RNIJKGL\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_5\,
            carryout => \scaler_4.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_6_c_RNIOUNN_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28334\,
            in2 => \_gnd_net_\,
            in3 => \N__26300\,
            lcout => \scaler_4.un3_source_data_0_cry_6_c_RNIOUNN\,
            ltout => OPEN,
            carryin => \scaler_4.un3_source_data_0_cry_6\,
            carryout => \scaler_4.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_7_c_RNIP0PN_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26624\,
            in2 => \N__28671\,
            in3 => \N__26297\,
            lcout => \scaler_4.un3_source_data_0_cry_7_c_RNIP0PN\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \scaler_4.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_cry_8_c_RNIS918_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26294\,
            lcout => \scaler_4.un3_source_data_0_cry_8_c_RNIS918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_RNO_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__26762\,
            in1 => \N__26739\,
            in2 => \_gnd_net_\,
            in3 => \N__26706\,
            lcout => \scaler_4.un2_source_data_0_cry_1_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.N_905_i_l_ofx_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28373\,
            in2 => \_gnd_net_\,
            in3 => \N__28354\,
            lcout => \scaler_4.N_905_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un2_source_data_0_cry_1_c_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26763\,
            in2 => \N__26618\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.source_data_1_esr_6_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26578\,
            in2 => \N__26770\,
            in3 => \N__26585\,
            lcout => scaler_4_data_6,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_1\,
            carryout => \scaler_4.un2_source_data_0_cry_2\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_7_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26536\,
            in2 => \N__26582\,
            in3 => \N__26543\,
            lcout => scaler_4_data_7,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_2\,
            carryout => \scaler_4.un2_source_data_0_cry_3\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_8_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26488\,
            in2 => \N__26540\,
            in3 => \N__26495\,
            lcout => scaler_4_data_8,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_3\,
            carryout => \scaler_4.un2_source_data_0_cry_4\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_9_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26443\,
            in2 => \N__26492\,
            in3 => \N__26450\,
            lcout => scaler_4_data_9,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_4\,
            carryout => \scaler_4.un2_source_data_0_cry_5\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_10_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26923\,
            in2 => \N__26447\,
            in3 => \N__26411\,
            lcout => scaler_4_data_10,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_5\,
            carryout => \scaler_4.un2_source_data_0_cry_6\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_11_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26881\,
            in2 => \N__26927\,
            in3 => \N__26888\,
            lcout => scaler_4_data_11,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_6\,
            carryout => \scaler_4.un2_source_data_0_cry_7\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_12_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26839\,
            in2 => \N__26885\,
            in3 => \N__26846\,
            lcout => scaler_4_data_12,
            ltout => OPEN,
            carryin => \scaler_4.un2_source_data_0_cry_7\,
            carryout => \scaler_4.un2_source_data_0_cry_8\,
            clk => \N__36051\,
            ce => \N__29570\,
            sr => \N__36732\
        );

    \scaler_4.source_data_1_esr_13_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26843\,
            in2 => \N__26828\,
            in3 => \N__26792\,
            lcout => scaler_4_data_13,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \scaler_4.un2_source_data_0_cry_9\,
            clk => \N__36044\,
            ce => \N__29569\,
            sr => \N__36737\
        );

    \scaler_4.source_data_1_esr_14_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26789\,
            lcout => scaler_4_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36044\,
            ce => \N__29569\,
            sr => \N__36737\
        );

    \scaler_4.source_data_1_esr_5_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26771\,
            in1 => \N__26740\,
            in2 => \_gnd_net_\,
            in3 => \N__26708\,
            lcout => scaler_4_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36044\,
            ce => \N__29569\,
            sr => \N__36737\
        );

    \scaler_4.source_data_1_4_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__36977\,
            in1 => \N__26741\,
            in2 => \N__26663\,
            in3 => \N__26707\,
            lcout => scaler_4_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36036\,
            ce => 'H',
            sr => \N__36742\
        );

    \ppm_encoder_1.elevator_esr_4_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32027\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.elevatorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36026\,
            ce => \N__27283\,
            sr => \N__36747\
        );

    \ppm_encoder_1.rudder_esr_4_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26662\,
            lcout => \ppm_encoder_1.rudderZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36026\,
            ce => \N__27283\,
            sr => \N__36747\
        );

    \ppm_encoder_1.rudder_esr_5_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27335\,
            lcout => \ppm_encoder_1.rudderZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36026\,
            ce => \N__27283\,
            sr => \N__36747\
        );

    \ppm_encoder_1.counter24_0_I_21_c_RNO_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__27212\,
            in2 => \N__27179\,
            in3 => \N__27417\,
            lcout => \ppm_encoder_1.counter24_0_I_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_6_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27224\,
            in1 => \N__27121\,
            in2 => \_gnd_net_\,
            in3 => \N__29093\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36020\,
            ce => \N__27013\,
            sr => \N__36753\
        );

    \ppm_encoder_1.pulses2count_esr_7_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27206\,
            in1 => \N__27118\,
            in2 => \_gnd_net_\,
            in3 => \N__27191\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36020\,
            ce => \N__27013\,
            sr => \N__36753\
        );

    \ppm_encoder_1.pulses2count_esr_12_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27170\,
            in1 => \N__27120\,
            in2 => \_gnd_net_\,
            in3 => \N__30452\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36020\,
            ce => \N__27013\,
            sr => \N__36753\
        );

    \ppm_encoder_1.counter24_0_I_39_c_RNO_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__27601\,
            in1 => \N__27158\,
            in2 => \N__27131\,
            in3 => \N__27631\,
            lcout => \ppm_encoder_1.counter24_0_I_39_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_13_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27117\,
            in1 => \N__29504\,
            in2 => \_gnd_net_\,
            in3 => \N__27140\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36020\,
            ce => \N__27013\,
            sr => \N__36753\
        );

    \ppm_encoder_1.pulses2count_esr_14_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27119\,
            in1 => \N__27044\,
            in2 => \_gnd_net_\,
            in3 => \N__27026\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36020\,
            ce => \N__27013\,
            sr => \N__36753\
        );

    \ppm_encoder_1.counter_0_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26943\,
            in2 => \N__26969\,
            in3 => \N__26968\,
            lcout => \ppm_encoder_1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_0\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_1_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27557\,
            in2 => \_gnd_net_\,
            in3 => \N__27536\,
            lcout => \ppm_encoder_1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_0\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_1\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_2_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27527\,
            in2 => \_gnd_net_\,
            in3 => \N__27509\,
            lcout => \ppm_encoder_1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_1\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_2\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_3_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27503\,
            in2 => \_gnd_net_\,
            in3 => \N__27485\,
            lcout => \ppm_encoder_1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_2\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_3\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_4_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27477\,
            in2 => \_gnd_net_\,
            in3 => \N__27455\,
            lcout => \ppm_encoder_1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_3\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_4\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_5_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27447\,
            in2 => \_gnd_net_\,
            in3 => \N__27425\,
            lcout => \ppm_encoder_1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_4\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_5\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_6_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27421\,
            in2 => \_gnd_net_\,
            in3 => \N__27401\,
            lcout => \ppm_encoder_1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_5\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_6\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_7_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27394\,
            in2 => \_gnd_net_\,
            in3 => \N__27374\,
            lcout => \ppm_encoder_1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_6\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_7\,
            clk => \N__36015\,
            ce => 'H',
            sr => \N__27974\
        );

    \ppm_encoder_1.counter_8_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27360\,
            in2 => \_gnd_net_\,
            in3 => \N__27338\,
            lcout => \ppm_encoder_1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_8\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_9_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27723\,
            in2 => \_gnd_net_\,
            in3 => \N__27701\,
            lcout => \ppm_encoder_1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_8\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_9\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_10_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27693\,
            in2 => \_gnd_net_\,
            in3 => \N__27671\,
            lcout => \ppm_encoder_1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_9\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_10\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_11_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27660\,
            in2 => \_gnd_net_\,
            in3 => \N__27638\,
            lcout => \ppm_encoder_1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_10\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_11\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_12_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27630\,
            in2 => \_gnd_net_\,
            in3 => \N__27608\,
            lcout => \ppm_encoder_1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_11\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_12\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_13_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27600\,
            in2 => \_gnd_net_\,
            in3 => \N__27578\,
            lcout => \ppm_encoder_1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_12\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_13\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_14_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30433\,
            in2 => \_gnd_net_\,
            in3 => \N__27575\,
            lcout => \ppm_encoder_1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_13\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_14\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_15_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30251\,
            in2 => \_gnd_net_\,
            in3 => \N__27572\,
            lcout => \ppm_encoder_1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_14\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_15\,
            clk => \N__36013\,
            ce => 'H',
            sr => \N__27973\
        );

    \ppm_encoder_1.counter_16_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30213\,
            in2 => \_gnd_net_\,
            in3 => \N__27569\,
            lcout => \ppm_encoder_1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_16\,
            clk => \N__36011\,
            ce => 'H',
            sr => \N__27972\
        );

    \ppm_encoder_1.counter_17_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30235\,
            in2 => \_gnd_net_\,
            in3 => \N__27566\,
            lcout => \ppm_encoder_1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \ppm_encoder_1.un1_counter_13_cry_16\,
            carryout => \ppm_encoder_1.un1_counter_13_cry_17\,
            clk => \N__36011\,
            ce => 'H',
            sr => \N__27972\
        );

    \ppm_encoder_1.counter_18_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30191\,
            in2 => \_gnd_net_\,
            in3 => \N__27977\,
            lcout => \ppm_encoder_1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36011\,
            ce => 'H',
            sr => \N__27972\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_12_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27922\,
            in1 => \N__27837\,
            in2 => \_gnd_net_\,
            in3 => \N__27803\,
            lcout => \ppm_encoder_1.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_3__0__0_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27773\,
            lcout => \uart_pc_sync.aux_3__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_2__0__0_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31022\,
            lcout => \uart_pc_sync.aux_2__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.Q_0__0_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27767\,
            lcout => \debug_CH2_18A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_0__0__0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone_sync.aux_0__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36150\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_1__0__0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27752\,
            lcout => \uart_drone_sync.aux_1__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_2__0__0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27743\,
            lcout => \uart_drone_sync.aux_2__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.aux_3__0__0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27737\,
            lcout => \uart_drone_sync.aux_3__0__0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNILP1J_9_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31988\,
            in2 => \_gnd_net_\,
            in3 => \N__33632\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.un1_state51_i_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__33633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36880\,
            lcout => \Commands_frame_decoder.un1_state51_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNII68S_9_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__36881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \Commands_frame_decoder.source_offset4data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_RNI6P6K_4_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32356\,
            in2 => \_gnd_net_\,
            in3 => \N__28092\,
            lcout => \dron_frame_decoder_1.un1_sink_data_valid_5_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_2_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__30821\,
            in1 => \N__31079\,
            in2 => \N__31477\,
            in3 => \N__28066\,
            lcout => \Commands_frame_decoder.N_338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_11_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__33624\,
            in1 => \N__27988\,
            in2 => \N__32300\,
            in3 => \N__32909\,
            lcout => \Commands_frame_decoder.stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36113\,
            ce => 'H',
            sr => \N__36703\
        );

    \Commands_frame_decoder.state_RNIQRI31_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__33623\,
            in1 => \N__27987\,
            in2 => \_gnd_net_\,
            in3 => \N__36879\,
            lcout => \Commands_frame_decoder.state_RNIQRI31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_10_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__28004\,
            in2 => \_gnd_net_\,
            in3 => \N__32873\,
            lcout => \Commands_frame_decoder.stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36113\,
            ce => 'H',
            sr => \N__36703\
        );

    \Commands_frame_decoder.state_7_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__32874\,
            in1 => \N__28176\,
            in2 => \N__33642\,
            in3 => \N__28277\,
            lcout => \Commands_frame_decoder.stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36113\,
            ce => 'H',
            sr => \N__36703\
        );

    \Commands_frame_decoder.state_RNIJN1J_7_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33622\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28276\,
            lcout => \Commands_frame_decoder.source_offset2data_1_sqmuxa\,
            ltout => \Commands_frame_decoder.source_offset2data_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_8_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28253\,
            in2 => \N__28256\,
            in3 => \N__32875\,
            lcout => \Commands_frame_decoder.stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36113\,
            ce => 'H',
            sr => \N__36703\
        );

    \Commands_frame_decoder.state_RNIKO1J_8_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28252\,
            in2 => \_gnd_net_\,
            in3 => \N__33562\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIMQ8T1_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33955\,
            in2 => \_gnd_net_\,
            in3 => \N__35076\,
            lcout => \uart_pc.timer_Count_RNIMQ8T1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_5_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__32406\,
            in1 => \N__28238\,
            in2 => \N__32120\,
            in3 => \N__32178\,
            lcout => \dron_frame_decoder_1.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36101\,
            ce => 'H',
            sr => \N__36710\
        );

    \Commands_frame_decoder.state_5_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__32868\,
            in1 => \N__28205\,
            in2 => \_gnd_net_\,
            in3 => \N__28217\,
            lcout => \Commands_frame_decoder.stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36101\,
            ce => 'H',
            sr => \N__36710\
        );

    \uart_pc.data_rdy_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36324\,
            in2 => \_gnd_net_\,
            in3 => \N__33956\,
            lcout => uart_pc_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36101\,
            ce => 'H',
            sr => \N__36710\
        );

    \Commands_frame_decoder.state_6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__32869\,
            in1 => \N__28169\,
            in2 => \_gnd_net_\,
            in3 => \N__28193\,
            lcout => \Commands_frame_decoder.stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36101\,
            ce => 'H',
            sr => \N__36710\
        );

    \Commands_frame_decoder.state_4_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__28133\,
            in1 => \N__28147\,
            in2 => \_gnd_net_\,
            in3 => \N__32867\,
            lcout => \Commands_frame_decoder.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36101\,
            ce => 'H',
            sr => \N__36710\
        );

    \uart_pc.data_6_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__31877\,
            in1 => \N__31725\,
            in2 => \N__31946\,
            in3 => \N__30921\,
            lcout => uart_pc_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNILR1B2_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__36314\,
            in1 => \N__35077\,
            in2 => \_gnd_net_\,
            in3 => \N__33953\,
            lcout => \uart_pc.timer_Count_RNILR1B2Z0Z_2\,
            ltout => \uart_pc.timer_Count_RNILR1B2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_4_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__31875\,
            in1 => \N__32696\,
            in2 => \N__28376\,
            in3 => \N__30682\,
            lcout => uart_pc_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIOU0N_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__37255\,
            in1 => \N__32471\,
            in2 => \_gnd_net_\,
            in3 => \N__36885\,
            lcout => \uart_drone.state_RNIOU0NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_4.un3_source_data_un3_source_data_0_axb_7_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28372\,
            in2 => \_gnd_net_\,
            in3 => \N__28355\,
            lcout => \scaler_4.un3_source_data_0_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__31876\,
            in1 => \N__30853\,
            in2 => \N__32732\,
            in3 => \N__31724\,
            lcout => uart_pc_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__31919\,
            in1 => \N__34362\,
            in2 => \N__28322\,
            in3 => \N__34264\,
            lcout => \uart_drone.data_AuxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \uart_drone.data_Aux_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__34265\,
            in1 => \N__28306\,
            in2 => \N__34379\,
            in3 => \N__32768\,
            lcout => \uart_drone.data_AuxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \uart_drone.data_Aux_2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__31586\,
            in1 => \N__34363\,
            in2 => \N__28295\,
            in3 => \N__34266\,
            lcout => \uart_drone.data_AuxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \uart_drone.data_Aux_3_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__34267\,
            in1 => \N__28414\,
            in2 => \N__34380\,
            in3 => \N__31568\,
            lcout => \uart_drone.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \uart_drone.data_Aux_5_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__34268\,
            in1 => \N__28402\,
            in2 => \N__34381\,
            in3 => \N__31574\,
            lcout => \uart_drone.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \uart_drone.data_Aux_6_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__31580\,
            in1 => \N__34364\,
            in2 => \N__28391\,
            in3 => \N__34269\,
            lcout => \uart_drone.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36086\,
            ce => 'H',
            sr => \N__34182\
        );

    \Commands_frame_decoder.source_CH3data_esr_0_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31492\,
            lcout => \frame_decoder_CH3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36077\,
            ce => \N__28472\,
            sr => \N__36721\
        );

    \Commands_frame_decoder.source_offset3data_esr_0_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31490\,
            lcout => \frame_decoder_OFF3data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_1_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_2_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_OFF3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_3_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31200\,
            lcout => \frame_decoder_OFF3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_4_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31651\,
            lcout => \frame_decoder_OFF3data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_5_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30715\,
            lcout => \frame_decoder_OFF3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_esr_6_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31356\,
            lcout => \frame_decoder_OFF3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_offset3data_ess_7_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30957\,
            lcout => \frame_decoder_OFF3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36066\,
            ce => \N__31928\,
            sr => \N__36725\
        );

    \Commands_frame_decoder.source_CH3data_esr_3_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31201\,
            lcout => \frame_decoder_CH3data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \Commands_frame_decoder.source_CH3data_esr_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \frame_decoder_CH3data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \Commands_frame_decoder.source_CH3data_esr_2_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30828\,
            lcout => \frame_decoder_CH3data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \Commands_frame_decoder.source_CH3data_esr_5_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30724\,
            lcout => \frame_decoder_CH3data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \Commands_frame_decoder.source_CH3data_esr_6_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31357\,
            lcout => \frame_decoder_CH3data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \Commands_frame_decoder.source_CH3data_ess_7_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30958\,
            lcout => \frame_decoder_CH3data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36057\,
            ce => \N__28468\,
            sr => \N__36728\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32045\,
            in2 => \N__32090\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_0_c_RNI10UK_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28436\,
            in2 => \N__28430\,
            in3 => \N__28418\,
            lcout => \scaler_3.un2_source_data_0\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_0\,
            carryout => \scaler_3.un3_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_1_c_RNI44VK_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28847\,
            in2 => \N__28841\,
            in3 => \N__28829\,
            lcout => \scaler_3.un3_source_data_0_cry_1_c_RNI44VK\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_1\,
            carryout => \scaler_3.un3_source_data_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_2_c_RNI780L_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28826\,
            in2 => \N__28817\,
            in3 => \N__28808\,
            lcout => \scaler_3.un3_source_data_0_cry_2_c_RNI780L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_2\,
            carryout => \scaler_3.un3_source_data_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_3_c_RNIAC1L_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28805\,
            in2 => \N__28793\,
            in3 => \N__28781\,
            lcout => \scaler_3.un3_source_data_0_cry_3_c_RNIAC1L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_3\,
            carryout => \scaler_3.un3_source_data_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_4_c_RNIDG2L_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28778\,
            in2 => \N__28772\,
            in3 => \N__28760\,
            lcout => \scaler_3.un3_source_data_0_cry_4_c_RNIDG2L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_4\,
            carryout => \scaler_3.un3_source_data_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_5_c_RNIGK3L_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28757\,
            in2 => \N__28751\,
            in3 => \N__28739\,
            lcout => \scaler_3.un3_source_data_0_cry_5_c_RNIGK3L\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_5\,
            carryout => \scaler_3.un3_source_data_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_6_c_RNILUAN_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28736\,
            in2 => \_gnd_net_\,
            in3 => \N__28721\,
            lcout => \scaler_3.un3_source_data_0_cry_6_c_RNILUAN\,
            ltout => OPEN,
            carryin => \scaler_3.un3_source_data_0_cry_6\,
            carryout => \scaler_3.un3_source_data_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_7_c_RNIM0CN_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29042\,
            in2 => \N__28657\,
            in3 => \N__28478\,
            lcout => \scaler_3.un3_source_data_0_cry_7_c_RNIM0CN\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \scaler_3.un3_source_data_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un3_source_data_un3_source_data_0_cry_8_c_RNIRV25_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28475\,
            lcout => \scaler_3.un3_source_data_0_cry_8_c_RNIRV25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.N_893_i_l_ofx_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29086\,
            in2 => \_gnd_net_\,
            in3 => \N__29062\,
            lcout => \scaler_3.N_893_i_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_RNO_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__29609\,
            in1 => \N__32091\,
            in2 => \_gnd_net_\,
            in3 => \N__32055\,
            lcout => \scaler_3.un2_source_data_0_cry_1_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.un2_source_data_0_cry_1_c_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29610\,
            in2 => \N__29036\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_3.source_data_1_esr_6_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28999\,
            in2 => \N__29617\,
            in3 => \N__29006\,
            lcout => scaler_3_data_6,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_1\,
            carryout => \scaler_3.un2_source_data_0_cry_2\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_7_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28954\,
            in2 => \N__29003\,
            in3 => \N__28961\,
            lcout => scaler_3_data_7,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_2\,
            carryout => \scaler_3.un2_source_data_0_cry_3\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_8_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28918\,
            in2 => \N__28958\,
            in3 => \N__28925\,
            lcout => scaler_3_data_8,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_3\,
            carryout => \scaler_3.un2_source_data_0_cry_4\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_9_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28879\,
            in2 => \N__28922\,
            in3 => \N__28886\,
            lcout => scaler_3_data_9,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_4\,
            carryout => \scaler_3.un2_source_data_0_cry_5\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_10_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29749\,
            in2 => \N__28883\,
            in3 => \N__28850\,
            lcout => scaler_3_data_10,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_5\,
            carryout => \scaler_3.un2_source_data_0_cry_6\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_11_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29716\,
            in2 => \N__29753\,
            in3 => \N__29723\,
            lcout => scaler_3_data_11,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_6\,
            carryout => \scaler_3.un2_source_data_0_cry_7\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_12_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29680\,
            in2 => \N__29720\,
            in3 => \N__29687\,
            lcout => scaler_3_data_12,
            ltout => OPEN,
            carryin => \scaler_3.un2_source_data_0_cry_7\,
            carryout => \scaler_3.un2_source_data_0_cry_8\,
            clk => \N__36037\,
            ce => \N__29568\,
            sr => \N__36743\
        );

    \scaler_3.source_data_1_esr_13_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29684\,
            in2 => \N__29669\,
            in3 => \N__29633\,
            lcout => scaler_3_data_13,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \scaler_3.un2_source_data_0_cry_9\,
            clk => \N__36027\,
            ce => \N__29567\,
            sr => \N__36748\
        );

    \scaler_3.source_data_1_esr_14_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29630\,
            lcout => scaler_3_data_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36027\,
            ce => \N__29567\,
            sr => \N__36748\
        );

    \scaler_3.source_data_1_esr_5_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__29618\,
            in1 => \N__32092\,
            in2 => \_gnd_net_\,
            in3 => \N__32059\,
            lcout => scaler_3_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36027\,
            ce => \N__29567\,
            sr => \N__36748\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_13_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29244\,
            in1 => \N__29546\,
            in2 => \_gnd_net_\,
            in3 => \N__29533\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_2_6_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29498\,
            in1 => \N__29333\,
            in2 => \_gnd_net_\,
            in3 => \N__29303\,
            lcout => OPEN,
            ltout => \ppm_encoder_1.N_298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_1_6_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29245\,
            in1 => \_gnd_net_\,
            in2 => \N__29126\,
            in3 => \N__29122\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_esr_RNO_0_12_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__30625\,
            in1 => \N__30571\,
            in2 => \_gnd_net_\,
            in3 => \N__30464\,
            lcout => \ppm_encoder_1.pulses2count_esr_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter24_0_I_45_c_RNO_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__30446\,
            in1 => \N__30249\,
            in2 => \N__29768\,
            in3 => \N__30429\,
            lcout => \ppm_encoder_1.counter24_0_I_45_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_16_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__30401\,
            in1 => \N__30367\,
            in2 => \N__30139\,
            in3 => \N__30085\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36012\,
            ce => 'H',
            sr => \N__36761\
        );

    \ppm_encoder_1.pulses2count_17_LC_8_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__30353\,
            in1 => \N__30322\,
            in2 => \N__30140\,
            in3 => \N__30086\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36012\,
            ce => 'H',
            sr => \N__36761\
        );

    \ppm_encoder_1.pulses2count_18_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__30084\,
            in1 => \N__30308\,
            in2 => \N__30275\,
            in3 => \N__30137\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36012\,
            ce => 'H',
            sr => \N__36761\
        );

    \ppm_encoder_1.counter24_0_I_57_c_RNO_LC_8_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__30189\,
            in1 => \N__30271\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ppm_encoder_1.counter24_0_I_57_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.counter_RNI637H_18_LC_8_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__30234\,
            in2 => \N__30215\,
            in3 => \N__30190\,
            lcout => \ppm_encoder_1.PPM_STATE_ns_0_a3_0_2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ppm_encoder_1.pulses2count_15_LC_8_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__30161\,
            in1 => \N__29767\,
            in2 => \N__30138\,
            in3 => \N__30083\,
            lcout => \ppm_encoder_1.pulses2countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36009\,
            ce => 'H',
            sr => \N__36765\
        );

    \uart_pc_sync.aux_1__0__0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31007\,
            lcout => \uart_pc_sync.aux_1__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc_sync.aux_0__0__0_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31016\,
            lcout => \uart_pc_sync.aux_0__0_Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_rdy_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34335\,
            in2 => \_gnd_net_\,
            in3 => \N__31544\,
            lcout => uart_drone_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36120\,
            ce => 'H',
            sr => \N__36699\
        );

    \Commands_frame_decoder.state_RNO_3_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30854\,
            in1 => \N__30973\,
            in2 => \N__31476\,
            in3 => \N__30729\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_i_a2_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__31055\,
            in1 => \N__31101\,
            in2 => \N__31001\,
            in3 => \N__30998\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__32872\,
            in1 => \N__31083\,
            in2 => \N__30992\,
            in3 => \N__31031\,
            lcout => \Commands_frame_decoder.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36114\,
            ce => 'H',
            sr => \N__36704\
        );

    \Commands_frame_decoder.state_RNO_1_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__30974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31445\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_0_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30855\,
            in1 => \N__31046\,
            in2 => \N__30752\,
            in3 => \N__30730\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_0_a3_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__31084\,
            in1 => \N__31102\,
            in2 => \N__30629\,
            in3 => \N__32871\,
            lcout => \Commands_frame_decoder.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36114\,
            ce => 'H',
            sr => \N__36704\
        );

    \uart_pc.state_RNO_0_2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110100"
        )
    port map (
            in0 => \N__36339\,
            in1 => \N__33250\,
            in2 => \N__33420\,
            in3 => \N__36894\,
            lcout => \uart_pc.state_srsts_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNI9E9J_2_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32590\,
            lcout => \uart_drone.N_126_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_1_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31636\,
            in2 => \_gnd_net_\,
            in3 => \N__31818\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.state_ns_i_a2_2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_ns_i_a2_2_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33621\,
            in1 => \N__31311\,
            in2 => \N__31109\,
            in3 => \N__31158\,
            lcout => \Commands_frame_decoder.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNI3NPK_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33467\,
            in2 => \_gnd_net_\,
            in3 => \N__31078\,
            lcout => \Commands_frame_decoder.N_308_2\,
            ltout => \Commands_frame_decoder.N_308_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.state_RNO_1_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100011"
        )
    port map (
            in0 => \N__31045\,
            in1 => \N__32290\,
            in2 => \N__31034\,
            in3 => \N__32908\,
            lcout => \Commands_frame_decoder.state_ns_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__31510\,
            in1 => \N__34324\,
            in2 => \_gnd_net_\,
            in3 => \N__36896\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100001111"
        )
    port map (
            in0 => \N__32278\,
            in1 => \N__32628\,
            in2 => \N__31025\,
            in3 => \N__32466\,
            lcout => \uart_drone.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIDGR31_2_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__32587\,
            in1 => \N__32325\,
            in2 => \N__32467\,
            in3 => \N__32627\,
            lcout => \uart_drone.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__31254\,
            in1 => \N__31511\,
            in2 => \N__34352\,
            in3 => \N__36899\,
            lcout => \uart_drone.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI40411_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__37236\,
            in1 => \N__32649\,
            in2 => \N__32543\,
            in3 => \N__32597\,
            lcout => \uart_drone.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__31415\,
            in1 => \N__31866\,
            in2 => \N__36194\,
            in3 => \N__31726\,
            lcout => uart_pc_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_5_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__31727\,
            in1 => \N__31964\,
            in2 => \N__31878\,
            in3 => \N__31307\,
            lcout => uart_pc_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__32534\,
            in1 => \N__34323\,
            in2 => \N__31256\,
            in3 => \N__36898\,
            lcout => OPEN,
            ltout => \uart_drone.state_srsts_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_2_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__31255\,
            in1 => \N__32650\,
            in2 => \N__31238\,
            in3 => \N__32598\,
            lcout => \uart_drone.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone_sync.Q_0__0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31235\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \debug_CH0_16A_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_3_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__31723\,
            in1 => \N__31143\,
            in2 => \N__35372\,
            in3 => \N__31880\,
            lcout => uart_pc_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36087\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIES9Q1_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__34331\,
            in1 => \N__31539\,
            in2 => \_gnd_net_\,
            in3 => \N__35020\,
            lcout => \uart_drone.timer_Count_RNIES9Q1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.source_data_valid_RNO_0_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33166\,
            in2 => \_gnd_net_\,
            in3 => \N__33492\,
            lcout => \Commands_frame_decoder.count_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNO_0_3_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__32600\,
            in1 => \N__37227\,
            in2 => \N__32542\,
            in3 => \N__32651\,
            lcout => \uart_drone.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__31879\,
            in1 => \N__31722\,
            in2 => \N__32753\,
            in3 => \N__31786\,
            lcout => uart_pc_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36087\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_4_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__31721\,
            in1 => \N__33954\,
            in2 => \N__31653\,
            in3 => \N__32710\,
            lcout => uart_pc_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36087\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_2_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__37189\,
            in1 => \N__37118\,
            in2 => \_gnd_net_\,
            in3 => \N__37061\,
            lcout => \uart_drone.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_6_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__37064\,
            in1 => \_gnd_net_\,
            in2 => \N__37132\,
            in3 => \N__37192\,
            lcout => \uart_drone.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_5_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__37063\,
            in1 => \_gnd_net_\,
            in2 => \N__37131\,
            in3 => \N__37191\,
            lcout => \uart_drone.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_3_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__37190\,
            in1 => \N__37119\,
            in2 => \_gnd_net_\,
            in3 => \N__37062\,
            lcout => \uart_drone.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIRC5U2_2_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31555\,
            in2 => \_gnd_net_\,
            in3 => \N__31540\,
            lcout => \uart_drone.data_rdyc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_6_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__32792\,
            in1 => \N__36352\,
            in2 => \N__31963\,
            in3 => \N__36234\,
            lcout => \uart_pc.data_AuxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36067\,
            ce => 'H',
            sr => \N__35675\
        );

    \uart_pc.data_Aux_7_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__36235\,
            in1 => \N__31939\,
            in2 => \N__36356\,
            in3 => \N__33859\,
            lcout => \uart_pc.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36067\,
            ce => 'H',
            sr => \N__35675\
        );

    \Commands_frame_decoder.state_RNIH58S_8_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32008\,
            in2 => \_gnd_net_\,
            in3 => \N__36893\,
            lcout => \Commands_frame_decoder.source_offset3data_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_0_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__37193\,
            in1 => \N__37133\,
            in2 => \_gnd_net_\,
            in3 => \N__37051\,
            lcout => \uart_drone.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI3M4C3_15_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__33312\,
            in1 => \N__33291\,
            in2 => \_gnd_net_\,
            in3 => \N__31901\,
            lcout => \dron_frame_decoder_1.WDT10_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI0JQQ_6_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33030\,
            in1 => \N__33051\,
            in2 => \_gnd_net_\,
            in3 => \N__33130\,
            lcout => \dron_frame_decoder_1.WDT10lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIM3K1_4_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32935\,
            in1 => \N__33100\,
            in2 => \N__33086\,
            in3 => \N__32920\,
            lcout => OPEN,
            ltout => \dron_frame_decoder_1.WDT_RNIM3K1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIATMH2_7_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__33115\,
            in1 => \N__32219\,
            in2 => \N__31910\,
            in3 => \N__31907\,
            lcout => \dron_frame_decoder_1.WDT10lt14_0\,
            ltout => \dron_frame_decoder_1.WDT10lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNIC5NL3_15_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__33292\,
            in1 => \N__33313\,
            in2 => \N__31895\,
            in3 => \N__32417\,
            lcout => \dron_frame_decoder_1.WDT_RNIC5NL3Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_RNI65RK1_10_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__33067\,
            in1 => \N__33031\,
            in2 => \N__33011\,
            in3 => \N__33052\,
            lcout => \dron_frame_decoder_1.WDT_RNI65RK1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.state_2_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__32107\,
            in1 => \N__32423\,
            in2 => \N__32213\,
            in3 => \N__32160\,
            lcout => \dron_frame_decoder_1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36028\,
            ce => 'H',
            sr => \N__36749\
        );

    \scaler_3.source_data_1_4_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011011000"
        )
    port map (
            in0 => \N__36969\,
            in1 => \N__32096\,
            in2 => \N__32026\,
            in3 => \N__32060\,
            lcout => scaler_3_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36016\,
            ce => 'H',
            sr => \N__36756\
        );

    \Commands_frame_decoder.state_9_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__32009\,
            in2 => \_gnd_net_\,
            in3 => \N__32870\,
            lcout => \Commands_frame_decoder.stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36108\,
            ce => 'H',
            sr => \N__36700\
        );

    \uart_drone.timer_Count_RNI5A9J_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__33224\,
            in1 => \N__33202\,
            in2 => \N__33227\,
            in3 => \_gnd_net_\,
            lcout => \uart_drone.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_10_11_0_\,
            carryout => \uart_drone.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32327\,
            in2 => \_gnd_net_\,
            in3 => \N__31973\,
            lcout => \uart_drone.timer_Count_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_1\,
            carryout => \uart_drone.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32599\,
            in2 => \_gnd_net_\,
            in3 => \N__31970\,
            lcout => \uart_drone.timer_Count_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_drone.un4_timer_Count_1_cry_2\,
            carryout => \uart_drone.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_4_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32643\,
            in2 => \_gnd_net_\,
            in3 => \N__31967\,
            lcout => \uart_drone.timer_Count_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__33191\,
            in1 => \N__32492\,
            in2 => \N__32261\,
            in3 => \N__35057\,
            lcout => \uart_drone.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__33226\,
            in1 => \N__32491\,
            in2 => \N__32260\,
            in3 => \N__35056\,
            lcout => \uart_drone.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_4_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__35055\,
            in1 => \N__32259\,
            in2 => \N__32501\,
            in3 => \N__32429\,
            lcout => \uart_drone.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.source_data_valid_2_sqmuxa_i_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32389\,
            in2 => \_gnd_net_\,
            in3 => \N__36883\,
            lcout => \dron_frame_decoder_1.source_data_valid_2_sqmuxa_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__35054\,
            in1 => \N__32258\,
            in2 => \N__32500\,
            in3 => \N__32333\,
            lcout => \uart_drone.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI9ADK1_4_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__32464\,
            in1 => \N__32309\,
            in2 => \N__32279\,
            in3 => \N__37247\,
            lcout => \uart_drone.un1_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNIG8P51_2_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__33629\,
            in1 => \N__33149\,
            in2 => \_gnd_net_\,
            in3 => \N__33490\,
            lcout => \Commands_frame_decoder.state_ns_i_a3_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNIDLVE1_2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__33630\,
            in2 => \N__33159\,
            in3 => \N__36892\,
            lcout => \Commands_frame_decoder.count_RNIDLVE1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNIAT1D1_4_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__32642\,
            in1 => \N__32465\,
            in2 => \N__35065\,
            in3 => \N__32274\,
            lcout => \uart_drone.N_143\,
            ltout => \uart_drone.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_3_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__35032\,
            in1 => \N__32242\,
            in2 => \N__32231\,
            in3 => \N__32228\,
            lcout => \uart_drone.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__35270\,
            in1 => \N__35348\,
            in2 => \N__33251\,
            in3 => \N__32660\,
            lcout => \uart_pc.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_RNI62411_4_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__32588\,
            in1 => \N__32644\,
            in2 => \N__37240\,
            in3 => \N__32460\,
            lcout => \uart_drone.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__33830\,
            in1 => \N__34472\,
            in2 => \_gnd_net_\,
            in3 => \N__34571\,
            lcout => \uart_pc.data_Auxce_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__35344\,
            in1 => \N__35269\,
            in2 => \N__33425\,
            in3 => \N__33903\,
            lcout => OPEN,
            ltout => \uart_pc.N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_3_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__35035\,
            in1 => \N__33971\,
            in2 => \N__32654\,
            in3 => \N__33424\,
            lcout => \uart_pc.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNIU8TV1_3_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32645\,
            in1 => \N__37327\,
            in2 => \_gnd_net_\,
            in3 => \N__32589\,
            lcout => \uart_drone.N_144_1\,
            ltout => \uart_drone.N_144_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_3_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__32552\,
            in1 => \N__32535\,
            in2 => \N__32510\,
            in3 => \N__35034\,
            lcout => \uart_drone.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.state_4_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__35033\,
            in1 => \N__32507\,
            in2 => \N__32499\,
            in3 => \N__37226\,
            lcout => \uart_drone.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIBLRB2_4_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__35297\,
            in1 => \N__34757\,
            in2 => \N__34697\,
            in3 => \N__33901\,
            lcout => \uart_pc.un1_state_2_0\,
            ltout => \uart_pc.un1_state_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_1_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__32749\,
            in1 => \N__32786\,
            in2 => \N__32756\,
            in3 => \N__36325\,
            lcout => \uart_pc.data_AuxZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36069\,
            ce => 'H',
            sr => \N__35679\
        );

    \uart_pc.data_Aux_2_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__36326\,
            in1 => \N__32738\,
            in2 => \N__32728\,
            in3 => \N__36216\,
            lcout => \uart_pc.data_AuxZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36069\,
            ce => 'H',
            sr => \N__35679\
        );

    \uart_pc.data_Aux_4_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__36327\,
            in1 => \N__32777\,
            in2 => \N__32711\,
            in3 => \N__36217\,
            lcout => \uart_pc.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36069\,
            ce => 'H',
            sr => \N__35679\
        );

    \uart_pc.data_Aux_5_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__36218\,
            in1 => \N__32993\,
            in2 => \N__32695\,
            in3 => \N__36328\,
            lcout => \uart_pc.data_AuxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36069\,
            ce => 'H',
            sr => \N__35679\
        );

    \Commands_frame_decoder.WDT_RNII19A1_4_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33745\,
            in1 => \N__33328\,
            in2 => \N__33731\,
            in3 => \N__33343\,
            lcout => \Commands_frame_decoder.WDT_RNII19A1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNID7P31_6_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33697\,
            in1 => \N__33775\,
            in2 => \_gnd_net_\,
            in3 => \N__33679\,
            lcout => OPEN,
            ltout => \Commands_frame_decoder.WDT8lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIUG2B4_7_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__33760\,
            in1 => \N__32666\,
            in2 => \N__32678\,
            in3 => \N__32675\,
            lcout => \Commands_frame_decoder.WDT8lt14_0\,
            ltout => \Commands_frame_decoder.WDT8lt14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_RNIF92K5_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__32805\,
            in1 => \N__34040\,
            in2 => \N__32669\,
            in3 => \N__34010\,
            lcout => \Commands_frame_decoder.state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNI2VDI1_10_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__33678\,
            in1 => \N__33696\,
            in2 => \N__33662\,
            in3 => \N__33712\,
            lcout => \Commands_frame_decoder.WDT_RNI2VDI1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_15_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__34041\,
            in1 => \N__34011\,
            in2 => \N__33640\,
            in3 => \N__32890\,
            lcout => \Commands_frame_decoder.N_303_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_RNIPRJG5_0_15_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010011"
        )
    port map (
            in0 => \N__32891\,
            in1 => \N__33617\,
            in2 => \N__34016\,
            in3 => \N__34042\,
            lcout => \Commands_frame_decoder.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.preinit_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__32806\,
            in1 => \_gnd_net_\,
            in2 => \N__33641\,
            in3 => \_gnd_net_\,
            lcout => \Commands_frame_decoder.preinitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36059\,
            ce => 'H',
            sr => \N__36722\
        );

    \uart_pc.state_RNIEAGS_4_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__33905\,
            in1 => \_gnd_net_\,
            in2 => \N__34756\,
            in3 => \N__36886\,
            lcout => \uart_pc.state_RNIEAGSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_6_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__34560\,
            in1 => \N__33814\,
            in2 => \_gnd_net_\,
            in3 => \N__34452\,
            lcout => \uart_pc.data_Auxce_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__33812\,
            in1 => \N__34450\,
            in2 => \_gnd_net_\,
            in3 => \N__34558\,
            lcout => \uart_pc.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_4_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__34559\,
            in1 => \N__33813\,
            in2 => \_gnd_net_\,
            in3 => \N__34451\,
            lcout => \uart_pc.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNI5UFA2_3_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__35326\,
            in1 => \_gnd_net_\,
            in2 => \N__35264\,
            in3 => \N__33858\,
            lcout => \uart_pc.N_144_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.data_Aux_RNO_0_1_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__37185\,
            in1 => \N__37127\,
            in2 => \_gnd_net_\,
            in3 => \N__37043\,
            lcout => \uart_drone.data_Auxce_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIITIF1_4_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110011"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__34747\,
            in2 => \N__35263\,
            in3 => \N__33904\,
            lcout => \uart_pc.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_5_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__33811\,
            in1 => \N__34449\,
            in2 => \_gnd_net_\,
            in3 => \N__34547\,
            lcout => \uart_pc.data_Auxce_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNO_0_2_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34500\,
            in2 => \_gnd_net_\,
            in3 => \N__34548\,
            lcout => \uart_pc.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_RNI4U6E1_2_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33810\,
            in1 => \N__34448\,
            in2 => \_gnd_net_\,
            in3 => \N__34546\,
            lcout => \uart_pc.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dron_frame_decoder_1.WDT_0_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32969\,
            in2 => \N__32984\,
            in3 => \N__32983\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_0\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32963\,
            in2 => \_gnd_net_\,
            in3 => \N__32957\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_0\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_1\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_2_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32954\,
            in2 => \_gnd_net_\,
            in3 => \N__32948\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_1\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_2\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_3_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32945\,
            in2 => \_gnd_net_\,
            in3 => \N__32939\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_2\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_3\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_4_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32936\,
            in2 => \_gnd_net_\,
            in3 => \N__32924\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_3\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_4\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_5_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32921\,
            in2 => \_gnd_net_\,
            in3 => \N__33134\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_4\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_5\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_6_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33131\,
            in2 => \_gnd_net_\,
            in3 => \N__33119\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_5\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_6\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_7_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33116\,
            in2 => \_gnd_net_\,
            in3 => \N__33104\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_6\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_7\,
            clk => \N__36039\,
            ce => 'H',
            sr => \N__33277\
        );

    \dron_frame_decoder_1.WDT_8_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33101\,
            in2 => \_gnd_net_\,
            in3 => \N__33089\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_8\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_9_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33085\,
            in2 => \_gnd_net_\,
            in3 => \N__33071\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_8\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_9\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_10_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33068\,
            in2 => \_gnd_net_\,
            in3 => \N__33056\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_9\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_10\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_11_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33053\,
            in2 => \_gnd_net_\,
            in3 => \N__33035\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_10\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_11\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_12_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33032\,
            in2 => \_gnd_net_\,
            in3 => \N__33014\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_11\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_12\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_13_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \_gnd_net_\,
            in3 => \N__32996\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_12\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_13\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_14_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33314\,
            in2 => \_gnd_net_\,
            in3 => \N__33299\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \dron_frame_decoder_1.un1_WDT_cry_13\,
            carryout => \dron_frame_decoder_1.un1_WDT_cry_14\,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \dron_frame_decoder_1.WDT_15_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33293\,
            in2 => \_gnd_net_\,
            in3 => \N__33296\,
            lcout => \dron_frame_decoder_1.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36030\,
            ce => 'H',
            sr => \N__33278\
        );

    \uart_pc.state_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__33249\,
            in1 => \N__36343\,
            in2 => \N__34718\,
            in3 => \N__36910\,
            lcout => \uart_pc.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.timer_Count_RNO_0_1_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33225\,
            in2 => \_gnd_net_\,
            in3 => \N__33203\,
            lcout => \uart_drone.timer_Count_RNO_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33826\,
            in1 => \N__34467\,
            in2 => \_gnd_net_\,
            in3 => \N__34566\,
            lcout => \uart_pc.data_Auxce_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_RNIE6P51_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33433\,
            in1 => \N__33612\,
            in2 => \_gnd_net_\,
            in3 => \N__33493\,
            lcout => \Commands_frame_decoder.CO0\,
            ltout => \Commands_frame_decoder.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__33448\,
            in1 => \_gnd_net_\,
            in2 => \N__33185\,
            in3 => \N__33175\,
            lcout => \Commands_frame_decoder.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_RNO_0_3_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__33825\,
            in1 => \N__34466\,
            in2 => \_gnd_net_\,
            in3 => \N__34565\,
            lcout => \uart_pc.data_Auxce_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_2_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__33449\,
            in1 => \N__33182\,
            in2 => \N__33167\,
            in3 => \N__33176\,
            lcout => \Commands_frame_decoder.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.count_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__33613\,
            in1 => \N__33494\,
            in2 => \N__33437\,
            in3 => \N__33447\,
            lcout => \Commands_frame_decoder.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIGRIF1_2_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__35268\,
            in1 => \N__35337\,
            in2 => \N__33419\,
            in3 => \N__33902\,
            lcout => \uart_pc.timer_Count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Commands_frame_decoder.WDT_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33377\,
            in2 => \N__33392\,
            in3 => \N__33391\,
            lcout => \Commands_frame_decoder.WDTZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_0\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33371\,
            in2 => \_gnd_net_\,
            in3 => \N__33365\,
            lcout => \Commands_frame_decoder.WDTZ0Z_1\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_0\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_1\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33362\,
            in2 => \_gnd_net_\,
            in3 => \N__33356\,
            lcout => \Commands_frame_decoder.WDTZ0Z_2\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_1\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_2\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33353\,
            in2 => \_gnd_net_\,
            in3 => \N__33347\,
            lcout => \Commands_frame_decoder.WDTZ0Z_3\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_2\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_3\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33344\,
            in2 => \_gnd_net_\,
            in3 => \N__33332\,
            lcout => \Commands_frame_decoder.WDTZ0Z_4\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_3\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_4\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_5_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33329\,
            in2 => \_gnd_net_\,
            in3 => \N__33317\,
            lcout => \Commands_frame_decoder.WDTZ0Z_5\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_4\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_5\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_6_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33776\,
            in2 => \_gnd_net_\,
            in3 => \N__33764\,
            lcout => \Commands_frame_decoder.WDTZ0Z_6\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_5\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_6\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_7_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33761\,
            in2 => \_gnd_net_\,
            in3 => \N__33749\,
            lcout => \Commands_frame_decoder.WDTZ0Z_7\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_6\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_7\,
            clk => \N__36060\,
            ce => 'H',
            sr => \N__33991\
        );

    \Commands_frame_decoder.WDT_8_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33746\,
            in2 => \_gnd_net_\,
            in3 => \N__33734\,
            lcout => \Commands_frame_decoder.WDTZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_8\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_9_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33730\,
            in2 => \_gnd_net_\,
            in3 => \N__33716\,
            lcout => \Commands_frame_decoder.WDTZ0Z_9\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_8\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_9\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_10_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33713\,
            in2 => \_gnd_net_\,
            in3 => \N__33701\,
            lcout => \Commands_frame_decoder.WDTZ0Z_10\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_9\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_10\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_11_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33698\,
            in2 => \_gnd_net_\,
            in3 => \N__33683\,
            lcout => \Commands_frame_decoder.WDTZ0Z_11\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_10\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_11\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_12_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33680\,
            in2 => \_gnd_net_\,
            in3 => \N__33665\,
            lcout => \Commands_frame_decoder.WDTZ0Z_12\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_11\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_12\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_13_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33661\,
            in2 => \_gnd_net_\,
            in3 => \N__33647\,
            lcout => \Commands_frame_decoder.WDTZ0Z_13\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_12\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_13\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_14_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34043\,
            in2 => \_gnd_net_\,
            in3 => \N__34022\,
            lcout => \Commands_frame_decoder.WDTZ0Z_14\,
            ltout => OPEN,
            carryin => \Commands_frame_decoder.un1_WDT_cry_13\,
            carryout => \Commands_frame_decoder.un1_WDT_cry_14\,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \Commands_frame_decoder.WDT_15_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34015\,
            in2 => \_gnd_net_\,
            in3 => \N__34019\,
            lcout => \Commands_frame_decoder.WDTZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36053\,
            ce => 'H',
            sr => \N__33995\
        );

    \uart_pc.state_4_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__33907\,
            in1 => \N__33970\,
            in2 => \N__35064\,
            in3 => \N__35152\,
            lcout => \uart_pc.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIPD2K1_2_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__35184\,
            in1 => \N__35324\,
            in2 => \N__35246\,
            in3 => \N__34746\,
            lcout => \uart_pc.data_rdyc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNIJOJC1_2_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37175\,
            in1 => \N__37126\,
            in2 => \_gnd_net_\,
            in3 => \N__37042\,
            lcout => \uart_drone.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIUPE73_3_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__34499\,
            in1 => \N__33906\,
            in2 => \_gnd_net_\,
            in3 => \N__33857\,
            lcout => \uart_pc.un1_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_3_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__35058\,
            in1 => \N__35114\,
            in2 => \N__35156\,
            in3 => \N__34679\,
            lcout => \uart_pc.timer_CountZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.bit_Count_0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000111000"
        )
    port map (
            in0 => \N__33911\,
            in1 => \N__34504\,
            in2 => \N__34570\,
            in3 => \N__33860\,
            lcout => \uart_pc.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36040\,
            ce => 'H',
            sr => \N__36733\
        );

    \uart_pc.bit_Count_2_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__34481\,
            in1 => \N__33824\,
            in2 => \N__34471\,
            in3 => \N__33836\,
            lcout => \uart_pc.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36040\,
            ce => 'H',
            sr => \N__36733\
        );

    \uart_pc.bit_Count_1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__34561\,
            in1 => \N__34462\,
            in2 => \N__34505\,
            in3 => \N__34480\,
            lcout => \uart_pc.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36040\,
            ce => 'H',
            sr => \N__36733\
        );

    \uart_drone.data_Aux_7_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__34378\,
            in1 => \N__34270\,
            in2 => \N__34405\,
            in3 => \N__37325\,
            lcout => \uart_drone.data_AuxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36031\,
            ce => 'H',
            sr => \N__34201\
        );

    \uart_drone.data_Aux_4_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__36989\,
            in1 => \N__34377\,
            in2 => \N__34219\,
            in3 => \N__34274\,
            lcout => \uart_drone.data_AuxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36021\,
            ce => 'H',
            sr => \N__34202\
        );

    \pid_alt.state_RNIH1EN_0_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34166\,
            in2 => \_gnd_net_\,
            in3 => \N__36878\,
            lcout => \pid_alt.state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__35548\,
            in1 => \N__34052\,
            in2 => \N__35468\,
            in3 => \N__35565\,
            lcout => \reset_module_System.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36078\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI9O1P_2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__34601\,
            in1 => \N__34622\,
            in2 => \N__34643\,
            in3 => \N__34064\,
            lcout => \reset_module_System.reset6_15\,
            ltout => \reset_module_System.reset6_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.reset_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35464\,
            in2 => \N__34067\,
            in3 => \N__35547\,
            lcout => reset_system,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36078\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_cry_1_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35534\,
            in2 => \N__35588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \reset_module_System.count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34063\,
            in2 => \_gnd_net_\,
            in3 => \N__34046\,
            lcout => \reset_module_System.count_1_2\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_1\,
            carryout => \reset_module_System.count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_3_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34621\,
            in2 => \_gnd_net_\,
            in3 => \N__34610\,
            lcout => \reset_module_System.countZ0Z_3\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_2\,
            carryout => \reset_module_System.count_1_cry_3\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_4_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34772\,
            in2 => \_gnd_net_\,
            in3 => \N__34607\,
            lcout => \reset_module_System.countZ0Z_4\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_3\,
            carryout => \reset_module_System.count_1_cry_4\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_5_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34798\,
            in2 => \_gnd_net_\,
            in3 => \N__34604\,
            lcout => \reset_module_System.countZ0Z_5\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_4\,
            carryout => \reset_module_System.count_1_cry_5\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_6_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34600\,
            in2 => \_gnd_net_\,
            in3 => \N__34589\,
            lcout => \reset_module_System.countZ0Z_6\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_5\,
            carryout => \reset_module_System.count_1_cry_6\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_7_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34814\,
            in2 => \_gnd_net_\,
            in3 => \N__34586\,
            lcout => \reset_module_System.countZ0Z_7\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_6\,
            carryout => \reset_module_System.count_1_cry_7\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_8_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34826\,
            in2 => \_gnd_net_\,
            in3 => \N__34583\,
            lcout => \reset_module_System.countZ0Z_8\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_7\,
            carryout => \reset_module_System.count_1_cry_8\,
            clk => \N__36068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34784\,
            in2 => \_gnd_net_\,
            in3 => \N__34580\,
            lcout => \reset_module_System.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \reset_module_System.count_1_cry_9\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_10_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35479\,
            in2 => \_gnd_net_\,
            in3 => \N__34577\,
            lcout => \reset_module_System.countZ0Z_10\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_9\,
            carryout => \reset_module_System.count_1_cry_10\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_11_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35506\,
            in2 => \_gnd_net_\,
            in3 => \N__34574\,
            lcout => \reset_module_System.countZ0Z_11\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_10\,
            carryout => \reset_module_System.count_1_cry_11\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_12_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35605\,
            in2 => \_gnd_net_\,
            in3 => \N__34667\,
            lcout => \reset_module_System.countZ0Z_12\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_11\,
            carryout => \reset_module_System.count_1_cry_12\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_13_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35402\,
            in2 => \_gnd_net_\,
            in3 => \N__34664\,
            lcout => \reset_module_System.countZ0Z_13\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_12\,
            carryout => \reset_module_System.count_1_cry_13\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_14_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35518\,
            in2 => \_gnd_net_\,
            in3 => \N__34661\,
            lcout => \reset_module_System.countZ0Z_14\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_13\,
            carryout => \reset_module_System.count_1_cry_14\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_15_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35429\,
            in2 => \_gnd_net_\,
            in3 => \N__34658\,
            lcout => \reset_module_System.countZ0Z_15\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_14\,
            carryout => \reset_module_System.count_1_cry_15\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_16_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35630\,
            in2 => \_gnd_net_\,
            in3 => \N__34655\,
            lcout => \reset_module_System.countZ0Z_16\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_15\,
            carryout => \reset_module_System.count_1_cry_16\,
            clk => \N__36058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_17_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35491\,
            in2 => \_gnd_net_\,
            in3 => \N__34652\,
            lcout => \reset_module_System.countZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \reset_module_System.count_1_cry_17\,
            clk => \N__36052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_18_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35644\,
            in2 => \_gnd_net_\,
            in3 => \N__34649\,
            lcout => \reset_module_System.countZ0Z_18\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_17\,
            carryout => \reset_module_System.count_1_cry_18\,
            clk => \N__36052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_19_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35441\,
            in2 => \_gnd_net_\,
            in3 => \N__34646\,
            lcout => \reset_module_System.countZ0Z_19\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_18\,
            carryout => \reset_module_System.count_1_cry_19\,
            clk => \N__36052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_20_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34639\,
            in2 => \_gnd_net_\,
            in3 => \N__34625\,
            lcout => \reset_module_System.countZ0Z_20\,
            ltout => OPEN,
            carryin => \reset_module_System.count_1_cry_19\,
            carryout => \reset_module_System.count_1_cry_20\,
            clk => \N__36052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_21_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35416\,
            in2 => \_gnd_net_\,
            in3 => \N__34760\,
            lcout => \reset_module_System.countZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_RNO_0_2_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37028\,
            in2 => \_gnd_net_\,
            in3 => \N__37286\,
            lcout => \uart_drone.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNIMQ8T1_4_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35292\,
            in1 => \N__34751\,
            in2 => \N__35256\,
            in3 => \N__35021\,
            lcout => \uart_pc.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_RNO_0_0_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__34708\,
            in1 => \N__36351\,
            in2 => \_gnd_net_\,
            in3 => \N__36897\,
            lcout => OPEN,
            ltout => \uart_pc.state_srsts_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.state_0_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__34752\,
            in1 => \N__35240\,
            in2 => \N__34721\,
            in3 => \N__35293\,
            lcout => \uart_pc.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIRP8S_1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__34847\,
            in1 => \N__35167\,
            in2 => \N__34850\,
            in3 => \_gnd_net_\,
            lcout => \uart_pc.un1_state_2_0_a3_0\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \uart_pc.un4_timer_Count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_2_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35189\,
            in3 => \N__34682\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_1\,
            carryout => \uart_pc.un4_timer_Count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35328\,
            in2 => \_gnd_net_\,
            in3 => \N__34673\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_pc.un4_timer_Count_1_cry_2\,
            carryout => \uart_pc.un4_timer_Count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_4_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35236\,
            in2 => \_gnd_net_\,
            in3 => \N__34670\,
            lcout => \uart_pc.timer_Count_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNIVT8S_2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35327\,
            in2 => \_gnd_net_\,
            in3 => \N__35185\,
            lcout => \uart_pc.N_126_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_4_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__35022\,
            in1 => \N__35108\,
            in2 => \N__35155\,
            in3 => \N__35276\,
            lcout => \uart_pc.timer_CountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_2_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__35195\,
            in1 => \N__35145\,
            in2 => \N__35115\,
            in3 => \N__35023\,
            lcout => \uart_pc.timer_CountZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_RNO_0_1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34848\,
            in2 => \_gnd_net_\,
            in3 => \N__35168\,
            lcout => OPEN,
            ltout => \uart_pc.timer_Count_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_1_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__35154\,
            in1 => \N__35024\,
            in2 => \N__35171\,
            in3 => \N__35119\,
            lcout => \uart_pc.timer_CountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.timer_Count_0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__34849\,
            in1 => \N__35153\,
            in2 => \N__35120\,
            in3 => \N__35025\,
            lcout => \uart_pc.timer_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36029\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI97FD_5_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34825\,
            in1 => \N__34813\,
            in2 => \N__34802\,
            in3 => \N__34783\,
            lcout => \reset_module_System.reset6_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIR9N6_1_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34771\,
            in2 => \_gnd_net_\,
            in3 => \N__35532\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIA72I1_16_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35645\,
            in1 => \N__35629\,
            in2 => \N__35618\,
            in3 => \N__35615\,
            lcout => OPEN,
            ltout => \reset_module_System.reset6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNIMJ304_12_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__35390\,
            in1 => \N__35609\,
            in2 => \N__35594\,
            in3 => \N__35585\,
            lcout => \reset_module_System.reset6_19\,
            ltout => \reset_module_System.reset6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__35587\,
            in1 => \N__35566\,
            in2 => \N__35591\,
            in3 => \N__35463\,
            lcout => \reset_module_System.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNO_0_1_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35586\,
            in2 => \_gnd_net_\,
            in3 => \N__35533\,
            lcout => OPEN,
            ltout => \reset_module_System.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__35462\,
            in1 => \N__35567\,
            in2 => \N__35552\,
            in3 => \N__35549\,
            lcout => \reset_module_System.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNISRMR1_10_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35519\,
            in1 => \N__35507\,
            in2 => \N__35495\,
            in3 => \N__35480\,
            lcout => \reset_module_System.reset6_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_module_System.count_RNI34OR1_21_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35440\,
            in1 => \N__35428\,
            in2 => \N__35417\,
            in3 => \N__35401\,
            lcout => \reset_module_System.reset6_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_3_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__35384\,
            in1 => \N__36344\,
            in2 => \N__35365\,
            in3 => \N__36230\,
            lcout => \uart_pc.data_AuxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36061\,
            ce => 'H',
            sr => \N__35683\
        );

    \uart_drone.state_RNI63LK2_3_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__37287\,
            in1 => \N__37328\,
            in2 => \_gnd_net_\,
            in3 => \N__37251\,
            lcout => \uart_drone.un1_state_7_0\,
            ltout => \uart_drone.un1_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_drone.bit_Count_1_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__37106\,
            in1 => \N__37041\,
            in2 => \N__37346\,
            in3 => \N__37288\,
            lcout => \uart_drone.bit_CountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36054\,
            ce => 'H',
            sr => \N__36734\
        );

    \uart_drone.bit_Count_2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__37107\,
            in1 => \N__37161\,
            in2 => \N__37343\,
            in3 => \N__37334\,
            lcout => \uart_drone.bit_CountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36054\,
            ce => 'H',
            sr => \N__36734\
        );

    \uart_drone.bit_Count_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010000110000"
        )
    port map (
            in0 => \N__37326\,
            in1 => \N__37289\,
            in2 => \N__37050\,
            in3 => \N__37256\,
            lcout => \uart_drone.bit_CountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36047\,
            ce => 'H',
            sr => \N__36738\
        );

    \uart_drone.data_Aux_RNO_0_4_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37174\,
            in1 => \N__37117\,
            in2 => \_gnd_net_\,
            in3 => \N__37029\,
            lcout => \uart_drone.data_Auxce_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \scaler_2.source_data_1_esr_ctle_14_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36965\,
            in2 => \_gnd_net_\,
            in3 => \N__36876\,
            lcout => \debug_CH3_20A_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_pc.data_Aux_0_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__36368\,
            in1 => \N__36345\,
            in2 => \N__36184\,
            in3 => \N__36236\,
            lcout => \uart_pc.data_AuxZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36071\,
            ce => 'H',
            sr => \N__35684\
        );
end \INTERFACE\;
